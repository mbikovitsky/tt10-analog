magic
tech sky130A
magscale 1 2
timestamp 1757770450
<< viali >>
rect 2145 17289 2179 17323
rect 2789 17289 2823 17323
rect 4077 17289 4111 17323
rect 7297 17289 7331 17323
rect 7941 17289 7975 17323
rect 9321 17289 9355 17323
rect 10149 17289 10183 17323
rect 12449 17289 12483 17323
rect 12909 17289 12943 17323
rect 18429 17289 18463 17323
rect 17233 17221 17267 17255
rect 24685 17221 24719 17255
rect 3433 17153 3467 17187
rect 4721 17153 4755 17187
rect 5365 17153 5399 17187
rect 15761 17153 15795 17187
rect 8769 17085 8803 17119
rect 8861 17085 8895 17119
rect 9229 17085 9263 17119
rect 10333 17085 10367 17119
rect 12081 17085 12115 17119
rect 12265 17085 12299 17119
rect 12725 17085 12759 17119
rect 16589 17085 16623 17119
rect 16773 17085 16807 17119
rect 17049 17085 17083 17119
rect 17417 17085 17451 17119
rect 17877 17085 17911 17119
rect 18245 17085 18279 17119
rect 19717 17085 19751 17119
rect 21649 17085 21683 17119
rect 22293 17085 22327 17119
rect 23029 17085 23063 17119
rect 23121 17085 23155 17119
rect 23489 17085 23523 17119
rect 24041 17085 24075 17119
rect 24317 17085 24351 17119
rect 24869 17085 24903 17119
rect 25513 17085 25547 17119
rect 26157 17085 26191 17119
rect 26801 17085 26835 17119
rect 15485 17017 15519 17051
rect 26617 17017 26651 17051
rect 8953 16949 8987 16983
rect 11897 16949 11931 16983
rect 15117 16949 15151 16983
rect 15577 16949 15611 16983
rect 16681 16949 16715 16983
rect 17601 16949 17635 16983
rect 17693 16949 17727 16983
rect 19533 16949 19567 16983
rect 21465 16949 21499 16983
rect 22109 16949 22143 16983
rect 22845 16949 22879 16983
rect 23305 16949 23339 16983
rect 23857 16949 23891 16983
rect 24133 16949 24167 16983
rect 25329 16949 25363 16983
rect 25973 16949 26007 16983
rect 1685 16745 1719 16779
rect 2145 16745 2179 16779
rect 5641 16745 5675 16779
rect 6285 16745 6319 16779
rect 9413 16745 9447 16779
rect 9873 16745 9907 16779
rect 11161 16745 11195 16779
rect 11529 16745 11563 16779
rect 13461 16745 13495 16779
rect 13829 16745 13863 16779
rect 15209 16745 15243 16779
rect 16313 16745 16347 16779
rect 16957 16745 16991 16779
rect 17509 16745 17543 16779
rect 19717 16745 19751 16779
rect 24685 16745 24719 16779
rect 10149 16677 10183 16711
rect 12050 16677 12084 16711
rect 16773 16677 16807 16711
rect 17233 16677 17267 16711
rect 17417 16677 17451 16711
rect 23029 16677 23063 16711
rect 1869 16609 1903 16643
rect 2329 16609 2363 16643
rect 4261 16609 4295 16643
rect 4528 16609 4562 16643
rect 6009 16609 6043 16643
rect 6469 16609 6503 16643
rect 6561 16609 6595 16643
rect 6745 16609 6779 16643
rect 7021 16609 7055 16643
rect 8300 16609 8334 16643
rect 9505 16609 9539 16643
rect 10517 16609 10551 16643
rect 11345 16609 11379 16643
rect 11713 16609 11747 16643
rect 11805 16609 11839 16643
rect 13645 16609 13679 16643
rect 14013 16609 14047 16643
rect 14473 16609 14507 16643
rect 15117 16609 15151 16643
rect 15577 16609 15611 16643
rect 15761 16609 15795 16643
rect 15945 16609 15979 16643
rect 16129 16609 16163 16643
rect 19266 16609 19300 16643
rect 20830 16609 20864 16643
rect 21465 16609 21499 16643
rect 21649 16609 21683 16643
rect 21925 16609 21959 16643
rect 22109 16609 22143 16643
rect 22477 16609 22511 16643
rect 22661 16609 22695 16643
rect 23213 16609 23247 16643
rect 23673 16609 23707 16643
rect 24041 16609 24075 16643
rect 24409 16609 24443 16643
rect 24961 16609 24995 16643
rect 6929 16541 6963 16575
rect 8033 16541 8067 16575
rect 15301 16541 15335 16575
rect 16865 16541 16899 16575
rect 17601 16541 17635 16575
rect 19533 16541 19567 16575
rect 21097 16541 21131 16575
rect 21281 16541 21315 16575
rect 22293 16541 22327 16575
rect 22845 16541 22879 16575
rect 23397 16541 23431 16575
rect 23489 16541 23523 16575
rect 5825 16473 5859 16507
rect 14289 16473 14323 16507
rect 14749 16473 14783 16507
rect 18153 16473 18187 16507
rect 7665 16405 7699 16439
rect 9873 16405 9907 16439
rect 10057 16405 10091 16439
rect 13185 16405 13219 16439
rect 16589 16405 16623 16439
rect 17969 16405 18003 16439
rect 23857 16405 23891 16439
rect 6469 16201 6503 16235
rect 8677 16201 8711 16235
rect 9045 16201 9079 16235
rect 12357 16201 12391 16235
rect 13921 16201 13955 16235
rect 18521 16201 18555 16235
rect 20361 16201 20395 16235
rect 4629 16133 4663 16167
rect 16589 16133 16623 16167
rect 17785 16133 17819 16167
rect 19993 16133 20027 16167
rect 3249 16065 3283 16099
rect 7849 16065 7883 16099
rect 10241 16065 10275 16099
rect 13001 16065 13035 16099
rect 14473 16065 14507 16099
rect 16773 16065 16807 16099
rect 2881 15997 2915 16031
rect 5273 15997 5307 16031
rect 5365 15997 5399 16031
rect 5457 15997 5491 16031
rect 5641 15997 5675 16031
rect 6285 15997 6319 16031
rect 8861 15997 8895 16031
rect 9137 15997 9171 16031
rect 11713 15997 11747 16031
rect 12081 15997 12115 16031
rect 15393 15997 15427 16031
rect 16313 15997 16347 16031
rect 16497 15997 16531 16031
rect 17233 15997 17267 16031
rect 17509 15997 17543 16031
rect 17601 15997 17635 16031
rect 17877 15997 17911 16031
rect 18061 15997 18095 16031
rect 18245 15997 18279 16031
rect 18337 15997 18371 16031
rect 19625 15997 19659 16031
rect 19901 15997 19935 16031
rect 20269 15997 20303 16031
rect 20361 15997 20395 16031
rect 20545 15997 20579 16031
rect 22937 15997 22971 16031
rect 23029 15997 23063 16031
rect 24041 15997 24075 16031
rect 3494 15929 3528 15963
rect 5733 15929 5767 15963
rect 7582 15929 7616 15963
rect 10486 15929 10520 15963
rect 11897 15929 11931 15963
rect 11989 15929 12023 15963
rect 12725 15929 12759 15963
rect 15025 15929 15059 15963
rect 17417 15929 17451 15963
rect 19533 15929 19567 15963
rect 19993 15929 20027 15963
rect 3065 15861 3099 15895
rect 4997 15861 5031 15895
rect 11621 15861 11655 15895
rect 12265 15861 12299 15895
rect 12817 15861 12851 15895
rect 14289 15861 14323 15895
rect 14381 15861 14415 15895
rect 16221 15861 16255 15895
rect 16957 15861 16991 15895
rect 20177 15861 20211 15895
rect 22753 15861 22787 15895
rect 23949 15861 23983 15895
rect 3341 15657 3375 15691
rect 7205 15657 7239 15691
rect 7297 15657 7331 15691
rect 10057 15657 10091 15691
rect 11345 15657 11379 15691
rect 13185 15657 13219 15691
rect 13553 15657 13587 15691
rect 14473 15657 14507 15691
rect 14933 15657 14967 15691
rect 19625 15657 19659 15691
rect 23213 15657 23247 15691
rect 4537 15589 4571 15623
rect 4629 15589 4663 15623
rect 5181 15589 5215 15623
rect 14841 15589 14875 15623
rect 15301 15589 15335 15623
rect 16405 15589 16439 15623
rect 17969 15589 18003 15623
rect 19962 15589 19996 15623
rect 3525 15521 3559 15555
rect 4445 15521 4479 15555
rect 4813 15521 4847 15555
rect 5089 15521 5123 15555
rect 5273 15521 5307 15555
rect 5457 15521 5491 15555
rect 5825 15521 5859 15555
rect 6081 15521 6115 15555
rect 7573 15521 7607 15555
rect 7665 15521 7699 15555
rect 7757 15521 7791 15555
rect 7941 15521 7975 15555
rect 11805 15521 11839 15555
rect 12633 15521 12667 15555
rect 15669 15521 15703 15555
rect 16129 15521 16163 15555
rect 16773 15521 16807 15555
rect 17785 15521 17819 15555
rect 18613 15521 18647 15555
rect 18797 15521 18831 15555
rect 19441 15521 19475 15555
rect 21833 15521 21867 15555
rect 22100 15521 22134 15555
rect 23857 15521 23891 15555
rect 24041 15521 24075 15555
rect 24308 15521 24342 15555
rect 3709 15453 3743 15487
rect 9413 15453 9447 15487
rect 9597 15453 9631 15487
rect 9689 15453 9723 15487
rect 11713 15453 11747 15487
rect 13645 15453 13679 15487
rect 13829 15453 13863 15487
rect 15025 15453 15059 15487
rect 18429 15453 18463 15487
rect 19717 15453 19751 15487
rect 4261 15385 4295 15419
rect 12081 15385 12115 15419
rect 23305 15385 23339 15419
rect 4905 15317 4939 15351
rect 11989 15317 12023 15351
rect 16957 15317 16991 15351
rect 21097 15317 21131 15351
rect 25421 15317 25455 15351
rect 4997 15113 5031 15147
rect 9413 15113 9447 15147
rect 10701 15113 10735 15147
rect 12633 15113 12667 15147
rect 14933 15113 14967 15147
rect 17693 15113 17727 15147
rect 24777 15113 24811 15147
rect 18153 15045 18187 15079
rect 20085 15045 20119 15079
rect 24317 15045 24351 15079
rect 5825 14977 5859 15011
rect 9689 14977 9723 15011
rect 13185 14977 13219 15011
rect 14105 14977 14139 15011
rect 25053 14977 25087 15011
rect 4629 14909 4663 14943
rect 4813 14909 4847 14943
rect 5365 14909 5399 14943
rect 5457 14909 5491 14943
rect 5549 14909 5583 14943
rect 5733 14909 5767 14943
rect 6377 14909 6411 14943
rect 9229 14909 9263 14943
rect 9597 14909 9631 14943
rect 10057 14909 10091 14943
rect 10149 14909 10183 14943
rect 10977 14909 11011 14943
rect 11069 14909 11103 14943
rect 11161 14909 11195 14943
rect 11345 14909 11379 14943
rect 12081 14909 12115 14943
rect 12265 14909 12299 14943
rect 12449 14909 12483 14943
rect 13001 14909 13035 14943
rect 15117 14909 15151 14943
rect 16037 14909 16071 14943
rect 16313 14909 16347 14943
rect 16405 14909 16439 14943
rect 17141 14909 17175 14943
rect 17509 14909 17543 14943
rect 18337 14909 18371 14943
rect 18705 14909 18739 14943
rect 24041 14909 24075 14943
rect 24317 14909 24351 14943
rect 24961 14909 24995 14943
rect 25605 14909 25639 14943
rect 5089 14841 5123 14875
rect 13921 14841 13955 14875
rect 16221 14841 16255 14875
rect 17325 14841 17359 14875
rect 17417 14841 17451 14875
rect 17877 14841 17911 14875
rect 18961 14841 18995 14875
rect 24133 14841 24167 14875
rect 24593 14841 24627 14875
rect 8677 14773 8711 14807
rect 10333 14773 10367 14807
rect 13093 14773 13127 14807
rect 13553 14773 13587 14807
rect 14013 14773 14047 14807
rect 16589 14773 16623 14807
rect 18521 14773 18555 14807
rect 24501 14773 24535 14807
rect 3709 14569 3743 14603
rect 7205 14569 7239 14603
rect 8953 14569 8987 14603
rect 9781 14569 9815 14603
rect 10701 14569 10735 14603
rect 12357 14569 12391 14603
rect 12817 14569 12851 14603
rect 13185 14569 13219 14603
rect 14565 14569 14599 14603
rect 17325 14569 17359 14603
rect 19349 14569 19383 14603
rect 21833 14569 21867 14603
rect 23121 14569 23155 14603
rect 24593 14569 24627 14603
rect 4629 14501 4663 14535
rect 4721 14501 4755 14535
rect 10057 14501 10091 14535
rect 13553 14501 13587 14535
rect 19789 14501 19823 14535
rect 22569 14501 22603 14535
rect 22937 14501 22971 14535
rect 23949 14501 23983 14535
rect 2596 14433 2630 14467
rect 3985 14433 4019 14467
rect 4537 14433 4571 14467
rect 4905 14433 4939 14467
rect 5825 14433 5859 14467
rect 6081 14433 6115 14467
rect 7573 14433 7607 14467
rect 7840 14433 7874 14467
rect 9413 14433 9447 14467
rect 12725 14433 12759 14467
rect 14933 14433 14967 14467
rect 17141 14433 17175 14467
rect 18245 14433 18279 14467
rect 18337 14433 18371 14467
rect 18521 14433 18555 14467
rect 19165 14433 19199 14467
rect 22109 14433 22143 14467
rect 22201 14433 22235 14467
rect 22293 14433 22327 14467
rect 22477 14433 22511 14467
rect 22753 14433 22787 14467
rect 23029 14433 23063 14467
rect 23121 14433 23155 14467
rect 23305 14433 23339 14467
rect 24409 14433 24443 14467
rect 25982 14433 26016 14467
rect 26249 14433 26283 14467
rect 2329 14365 2363 14399
rect 4169 14365 4203 14399
rect 9321 14365 9355 14399
rect 10241 14365 10275 14399
rect 10333 14365 10367 14399
rect 12909 14365 12943 14399
rect 13645 14365 13679 14399
rect 13737 14365 13771 14399
rect 15025 14365 15059 14399
rect 15117 14365 15151 14399
rect 16957 14365 16991 14399
rect 19533 14365 19567 14399
rect 24317 14365 24351 14399
rect 3801 14297 3835 14331
rect 4353 14297 4387 14331
rect 24869 14297 24903 14331
rect 9137 14229 9171 14263
rect 20913 14229 20947 14263
rect 24041 14229 24075 14263
rect 2789 14025 2823 14059
rect 11989 14025 12023 14059
rect 14749 14025 14783 14059
rect 18153 14025 18187 14059
rect 21189 14025 21223 14059
rect 23857 14025 23891 14059
rect 25421 14025 25455 14059
rect 25513 14025 25547 14059
rect 25697 14025 25731 14059
rect 3893 13957 3927 13991
rect 8401 13957 8435 13991
rect 9137 13957 9171 13991
rect 14657 13957 14691 13991
rect 17509 13957 17543 13991
rect 19533 13957 19567 13991
rect 5273 13889 5307 13923
rect 9781 13889 9815 13923
rect 10057 13889 10091 13923
rect 10425 13889 10459 13923
rect 12633 13889 12667 13923
rect 14013 13889 14047 13923
rect 15301 13889 15335 13923
rect 21925 13889 21959 13923
rect 22385 13889 22419 13923
rect 25237 13889 25271 13923
rect 25605 13889 25639 13923
rect 2973 13821 3007 13855
rect 5641 13821 5675 13855
rect 5733 13821 5767 13855
rect 5825 13821 5859 13855
rect 6009 13821 6043 13855
rect 7849 13821 7883 13855
rect 8033 13821 8067 13855
rect 8677 13821 8711 13855
rect 8769 13821 8803 13855
rect 8861 13821 8895 13855
rect 9045 13821 9079 13855
rect 9321 13821 9355 13855
rect 9413 13821 9447 13855
rect 9505 13821 9539 13855
rect 9689 13821 9723 13855
rect 9965 13821 9999 13855
rect 11621 13821 11655 13855
rect 11713 13821 11747 13855
rect 16957 13821 16991 13855
rect 17233 13821 17267 13855
rect 17325 13821 17359 13855
rect 17601 13821 17635 13855
rect 17969 13821 18003 13855
rect 18705 13821 18739 13855
rect 18889 13821 18923 13855
rect 19073 13821 19107 13855
rect 19349 13821 19383 13855
rect 19809 13821 19843 13855
rect 20065 13821 20099 13855
rect 21281 13821 21315 13855
rect 21465 13821 21499 13855
rect 21833 13821 21867 13855
rect 25329 13821 25363 13855
rect 25697 13821 25731 13855
rect 25881 13821 25915 13855
rect 5028 13753 5062 13787
rect 5365 13753 5399 13787
rect 8217 13753 8251 13787
rect 11253 13753 11287 13787
rect 15117 13753 15151 13787
rect 17141 13753 17175 13787
rect 17785 13753 17819 13787
rect 17877 13753 17911 13787
rect 24970 13753 25004 13787
rect 11897 13685 11931 13719
rect 12357 13685 12391 13719
rect 12449 13685 12483 13719
rect 14197 13685 14231 13719
rect 14289 13685 14323 13719
rect 15209 13685 15243 13719
rect 5457 13481 5491 13515
rect 8953 13481 8987 13515
rect 13093 13481 13127 13515
rect 13461 13481 13495 13515
rect 14565 13481 14599 13515
rect 24317 13481 24351 13515
rect 25237 13481 25271 13515
rect 4445 13413 4479 13447
rect 12725 13413 12759 13447
rect 16313 13413 16347 13447
rect 25605 13413 25639 13447
rect 4353 13345 4387 13379
rect 4537 13345 4571 13379
rect 4721 13345 4755 13379
rect 4813 13345 4847 13379
rect 7573 13345 7607 13379
rect 7840 13345 7874 13379
rect 9229 13345 9263 13379
rect 11233 13345 11267 13379
rect 12449 13345 12483 13379
rect 12633 13345 12667 13379
rect 12817 13345 12851 13379
rect 14933 13345 14967 13379
rect 16129 13345 16163 13379
rect 16405 13345 16439 13379
rect 16497 13345 16531 13379
rect 16957 13345 16991 13379
rect 17509 13345 17543 13379
rect 21465 13345 21499 13379
rect 21833 13345 21867 13379
rect 24041 13345 24075 13379
rect 24777 13345 24811 13379
rect 25053 13345 25087 13379
rect 25145 13345 25179 13379
rect 25421 13345 25455 13379
rect 25697 13345 25731 13379
rect 25881 13345 25915 13379
rect 6377 13277 6411 13311
rect 9321 13277 9355 13311
rect 9689 13277 9723 13311
rect 10977 13277 11011 13311
rect 13553 13277 13587 13311
rect 13737 13277 13771 13311
rect 15025 13277 15059 13311
rect 15117 13277 15151 13311
rect 17141 13277 17175 13311
rect 17785 13277 17819 13311
rect 21557 13277 21591 13311
rect 21741 13277 21775 13311
rect 22477 13277 22511 13311
rect 23857 13277 23891 13311
rect 23949 13277 23983 13311
rect 24133 13277 24167 13311
rect 9045 13209 9079 13243
rect 12357 13209 12391 13243
rect 16681 13209 16715 13243
rect 4169 13141 4203 13175
rect 5825 13141 5859 13175
rect 13001 13141 13035 13175
rect 16773 13141 16807 13175
rect 24593 13141 24627 13175
rect 24961 13141 24995 13175
rect 25789 13141 25823 13175
rect 4997 12937 5031 12971
rect 6929 12937 6963 12971
rect 8401 12937 8435 12971
rect 10977 12937 11011 12971
rect 17601 12937 17635 12971
rect 20545 12937 20579 12971
rect 23949 12937 23983 12971
rect 24133 12937 24167 12971
rect 25145 12937 25179 12971
rect 18245 12869 18279 12903
rect 3709 12801 3743 12835
rect 6377 12801 6411 12835
rect 12357 12801 12391 12835
rect 12541 12801 12575 12835
rect 16221 12801 16255 12835
rect 19165 12801 19199 12835
rect 21281 12801 21315 12835
rect 21465 12801 21499 12835
rect 23581 12801 23615 12835
rect 25513 12801 25547 12835
rect 3065 12733 3099 12767
rect 3433 12733 3467 12767
rect 3617 12733 3651 12767
rect 3893 12733 3927 12767
rect 3985 12733 4019 12767
rect 4445 12733 4479 12767
rect 4537 12733 4571 12767
rect 4813 12733 4847 12767
rect 8585 12733 8619 12767
rect 9505 12733 9539 12767
rect 9689 12733 9723 12767
rect 9781 12733 9815 12767
rect 9873 12733 9907 12767
rect 10333 12733 10367 12767
rect 10517 12733 10551 12767
rect 11253 12733 11287 12767
rect 11345 12733 11379 12767
rect 11437 12733 11471 12767
rect 11621 12733 11655 12767
rect 12725 12733 12759 12767
rect 12909 12733 12943 12767
rect 13001 12733 13035 12767
rect 14841 12733 14875 12767
rect 15945 12733 15979 12767
rect 17693 12733 17727 12767
rect 17877 12733 17911 12767
rect 18061 12733 18095 12767
rect 18705 12733 18739 12767
rect 18889 12733 18923 12767
rect 21189 12733 21223 12767
rect 21557 12733 21591 12767
rect 23489 12733 23523 12767
rect 23673 12733 23707 12767
rect 24501 12733 24535 12767
rect 25329 12733 25363 12767
rect 25421 12733 25455 12767
rect 25780 12733 25814 12767
rect 4629 12665 4663 12699
rect 6110 12665 6144 12699
rect 8217 12665 8251 12699
rect 11805 12665 11839 12699
rect 16477 12665 16511 12699
rect 17969 12665 18003 12699
rect 19432 12665 19466 12699
rect 22201 12665 22235 12699
rect 24317 12665 24351 12699
rect 25145 12665 25179 12699
rect 2881 12597 2915 12631
rect 3249 12597 3283 12631
rect 4261 12597 4295 12631
rect 10057 12597 10091 12631
rect 10149 12597 10183 12631
rect 13185 12597 13219 12631
rect 14749 12597 14783 12631
rect 16129 12597 16163 12631
rect 19073 12597 19107 12631
rect 24107 12597 24141 12631
rect 25053 12597 25087 12631
rect 26893 12597 26927 12631
rect 5365 12393 5399 12427
rect 5825 12393 5859 12427
rect 8861 12393 8895 12427
rect 12265 12393 12299 12427
rect 18429 12393 18463 12427
rect 19165 12393 19199 12427
rect 23423 12393 23457 12427
rect 25605 12393 25639 12427
rect 23213 12325 23247 12359
rect 2780 12257 2814 12291
rect 3985 12257 4019 12291
rect 4252 12257 4286 12291
rect 6101 12257 6135 12291
rect 6193 12257 6227 12291
rect 6285 12257 6319 12291
rect 6469 12257 6503 12291
rect 7849 12257 7883 12291
rect 8033 12257 8067 12291
rect 8401 12257 8435 12291
rect 8677 12257 8711 12291
rect 9209 12257 9243 12291
rect 10977 12257 11011 12291
rect 13461 12257 13495 12291
rect 13829 12257 13863 12291
rect 14013 12257 14047 12291
rect 14841 12257 14875 12291
rect 14933 12257 14967 12291
rect 15301 12257 15335 12291
rect 15393 12257 15427 12291
rect 16773 12257 16807 12291
rect 17141 12257 17175 12291
rect 17233 12257 17267 12291
rect 17509 12257 17543 12291
rect 17693 12257 17727 12291
rect 18061 12257 18095 12291
rect 18245 12257 18279 12291
rect 18981 12257 19015 12291
rect 19441 12257 19475 12291
rect 19625 12257 19659 12291
rect 19993 12257 20027 12291
rect 20177 12257 20211 12291
rect 21465 12257 21499 12291
rect 21833 12257 21867 12291
rect 22477 12257 22511 12291
rect 24878 12257 24912 12291
rect 25145 12257 25179 12291
rect 25237 12257 25271 12291
rect 25513 12257 25547 12291
rect 2513 12189 2547 12223
rect 8309 12189 8343 12223
rect 8953 12189 8987 12223
rect 13277 12189 13311 12223
rect 16865 12189 16899 12223
rect 21557 12189 21591 12223
rect 21741 12189 21775 12223
rect 10333 12121 10367 12155
rect 14473 12121 14507 12155
rect 3893 12053 3927 12087
rect 7665 12053 7699 12087
rect 13093 12053 13127 12087
rect 16405 12053 16439 12087
rect 20361 12053 20395 12087
rect 23397 12053 23431 12087
rect 23581 12053 23615 12087
rect 23765 12053 23799 12087
rect 25329 12053 25363 12087
rect 2973 11849 3007 11883
rect 11989 11849 12023 11883
rect 21281 11849 21315 11883
rect 22937 11849 22971 11883
rect 5089 11713 5123 11747
rect 17693 11713 17727 11747
rect 2789 11645 2823 11679
rect 4997 11645 5031 11679
rect 5365 11645 5399 11679
rect 5549 11645 5583 11679
rect 6101 11645 6135 11679
rect 6285 11645 6319 11679
rect 6653 11645 6687 11679
rect 6745 11645 6779 11679
rect 7389 11645 7423 11679
rect 7481 11645 7515 11679
rect 7573 11645 7607 11679
rect 7665 11645 7699 11679
rect 7849 11645 7883 11679
rect 8401 11645 8435 11679
rect 9597 11645 9631 11679
rect 9781 11645 9815 11679
rect 10149 11645 10183 11679
rect 10333 11645 10367 11679
rect 11161 11645 11195 11679
rect 11345 11645 11379 11679
rect 11713 11645 11747 11679
rect 11805 11645 11839 11679
rect 13369 11645 13403 11679
rect 14473 11645 14507 11679
rect 14565 11645 14599 11679
rect 14933 11645 14967 11679
rect 15025 11645 15059 11679
rect 17049 11645 17083 11679
rect 17233 11645 17267 11679
rect 17509 11645 17543 11679
rect 18061 11645 18095 11679
rect 22661 11645 22695 11679
rect 23213 11645 23247 11679
rect 23397 11645 23431 11679
rect 24869 11645 24903 11679
rect 24961 11645 24995 11679
rect 13124 11577 13158 11611
rect 16405 11577 16439 11611
rect 16865 11577 16899 11611
rect 18705 11577 18739 11611
rect 22394 11577 22428 11611
rect 23121 11577 23155 11611
rect 25228 11577 25262 11611
rect 4629 11509 4663 11543
rect 5733 11509 5767 11543
rect 7205 11509 7239 11543
rect 9045 11509 9079 11543
rect 9413 11509 9447 11543
rect 10977 11509 11011 11543
rect 15485 11509 15519 11543
rect 16681 11509 16715 11543
rect 17325 11509 17359 11543
rect 18245 11509 18279 11543
rect 19993 11509 20027 11543
rect 22753 11509 22787 11543
rect 22921 11509 22955 11543
rect 23213 11509 23247 11543
rect 24225 11509 24259 11543
rect 26341 11509 26375 11543
rect 6193 11305 6227 11339
rect 8125 11305 8159 11339
rect 8217 11305 8251 11339
rect 9321 11305 9355 11339
rect 13737 11305 13771 11339
rect 23689 11305 23723 11339
rect 24501 11305 24535 11339
rect 25329 11305 25363 11339
rect 7012 11237 7046 11271
rect 8401 11237 8435 11271
rect 8861 11237 8895 11271
rect 11529 11237 11563 11271
rect 19257 11237 19291 11271
rect 21557 11237 21591 11271
rect 23489 11237 23523 11271
rect 24777 11237 24811 11271
rect 3157 11169 3191 11203
rect 3341 11169 3375 11203
rect 4905 11169 4939 11203
rect 5089 11169 5123 11203
rect 5457 11169 5491 11203
rect 6009 11169 6043 11203
rect 6745 11169 6779 11203
rect 8585 11169 8619 11203
rect 9045 11169 9079 11203
rect 11161 11169 11195 11203
rect 11254 11169 11288 11203
rect 11437 11169 11471 11203
rect 11667 11169 11701 11203
rect 12624 11169 12658 11203
rect 16221 11169 16255 11203
rect 16488 11169 16522 11203
rect 18337 11169 18371 11203
rect 18521 11169 18555 11203
rect 18889 11169 18923 11203
rect 19533 11169 19567 11203
rect 19625 11169 19659 11203
rect 19717 11169 19751 11203
rect 19901 11169 19935 11203
rect 23305 11169 23339 11203
rect 25513 11169 25547 11203
rect 26157 11169 26191 11203
rect 4445 11101 4479 11135
rect 5365 11101 5399 11135
rect 5825 11101 5859 11135
rect 9873 11101 9907 11135
rect 12357 11101 12391 11135
rect 18613 11101 18647 11135
rect 18705 11101 18739 11135
rect 24041 11101 24075 11135
rect 24133 11101 24167 11135
rect 24225 11101 24259 11135
rect 24317 11101 24351 11135
rect 25789 11101 25823 11135
rect 25881 11101 25915 11135
rect 17601 11033 17635 11067
rect 19073 11033 19107 11067
rect 23857 11033 23891 11067
rect 25145 11033 25179 11067
rect 3341 10965 3375 10999
rect 8677 10965 8711 10999
rect 11805 10965 11839 10999
rect 23673 10965 23707 10999
rect 25237 10965 25271 10999
rect 25697 10965 25731 10999
rect 25973 10965 26007 10999
rect 26065 10965 26099 10999
rect 9781 10761 9815 10795
rect 12633 10761 12667 10795
rect 15577 10761 15611 10795
rect 16313 10761 16347 10795
rect 18705 10761 18739 10795
rect 20177 10761 20211 10795
rect 21281 10761 21315 10795
rect 22109 10761 22143 10795
rect 22201 10761 22235 10795
rect 23949 10761 23983 10795
rect 4629 10693 4663 10727
rect 7941 10693 7975 10727
rect 16589 10693 16623 10727
rect 22937 10693 22971 10727
rect 24133 10693 24167 10727
rect 25789 10693 25823 10727
rect 5273 10625 5307 10659
rect 5457 10625 5491 10659
rect 17969 10625 18003 10659
rect 21465 10625 21499 10659
rect 22477 10625 22511 10659
rect 22569 10625 22603 10659
rect 1685 10557 1719 10591
rect 3249 10557 3283 10591
rect 3505 10557 3539 10591
rect 5641 10557 5675 10591
rect 7573 10557 7607 10591
rect 7757 10557 7791 10591
rect 7849 10557 7883 10591
rect 8033 10557 8067 10591
rect 8401 10557 8435 10591
rect 11253 10557 11287 10591
rect 11401 10557 11435 10591
rect 11718 10557 11752 10591
rect 11989 10557 12023 10591
rect 12173 10557 12207 10591
rect 12265 10557 12299 10591
rect 12357 10557 12391 10591
rect 12725 10557 12759 10591
rect 12909 10557 12943 10591
rect 13001 10557 13035 10591
rect 13093 10557 13127 10591
rect 14197 10557 14231 10591
rect 16497 10557 16531 10591
rect 16681 10557 16715 10591
rect 16773 10557 16807 10591
rect 16957 10557 16991 10591
rect 19829 10557 19863 10591
rect 20085 10557 20119 10591
rect 20361 10557 20395 10591
rect 20545 10557 20579 10591
rect 21097 10557 21131 10591
rect 21281 10557 21315 10591
rect 21741 10557 21775 10591
rect 22385 10557 22419 10591
rect 22661 10557 22695 10591
rect 23489 10557 23523 10591
rect 23683 10557 23717 10591
rect 23857 10557 23891 10591
rect 24041 10557 24075 10591
rect 24685 10557 24719 10591
rect 24777 10557 24811 10591
rect 25605 10557 25639 10591
rect 25881 10557 25915 10591
rect 1952 10489 1986 10523
rect 8217 10489 8251 10523
rect 8646 10489 8680 10523
rect 11529 10489 11563 10523
rect 11621 10489 11655 10523
rect 13369 10489 13403 10523
rect 14442 10489 14476 10523
rect 23305 10489 23339 10523
rect 24317 10489 24351 10523
rect 24501 10489 24535 10523
rect 3065 10421 3099 10455
rect 4721 10421 4755 10455
rect 5825 10421 5859 10455
rect 11897 10421 11931 10455
rect 17417 10421 17451 10455
rect 20913 10421 20947 10455
rect 21649 10421 21683 10455
rect 22845 10421 22879 10455
rect 23489 10421 23523 10455
rect 25421 10421 25455 10455
rect 2513 10217 2547 10251
rect 4261 10217 4295 10251
rect 6193 10217 6227 10251
rect 17049 10217 17083 10251
rect 18521 10217 18555 10251
rect 25237 10217 25271 10251
rect 9597 10149 9631 10183
rect 9873 10149 9907 10183
rect 11437 10149 11471 10183
rect 17233 10149 17267 10183
rect 17417 10149 17451 10183
rect 18245 10149 18279 10183
rect 19248 10149 19282 10183
rect 23489 10149 23523 10183
rect 23673 10149 23707 10183
rect 24409 10149 24443 10183
rect 2053 10081 2087 10115
rect 2237 10081 2271 10115
rect 2697 10081 2731 10115
rect 3709 10081 3743 10115
rect 3985 10081 4019 10115
rect 4169 10081 4203 10115
rect 4537 10081 4571 10115
rect 4905 10081 4939 10115
rect 5089 10081 5123 10115
rect 5457 10081 5491 10115
rect 5917 10081 5951 10115
rect 6009 10081 6043 10115
rect 7389 10081 7423 10115
rect 7656 10081 7690 10115
rect 10057 10081 10091 10115
rect 11069 10081 11103 10115
rect 11217 10081 11251 10115
rect 11345 10081 11379 10115
rect 11534 10081 11568 10115
rect 11805 10081 11839 10115
rect 11989 10081 12023 10115
rect 12081 10081 12115 10115
rect 12173 10081 12207 10115
rect 12541 10081 12575 10115
rect 12797 10081 12831 10115
rect 17969 10081 18003 10115
rect 18153 10081 18187 10115
rect 18383 10081 18417 10115
rect 21281 10081 21315 10115
rect 21548 10081 21582 10115
rect 23029 10081 23063 10115
rect 23305 10081 23339 10115
rect 24593 10081 24627 10115
rect 24869 10081 24903 10115
rect 25053 10081 25087 10115
rect 25145 10081 25179 10115
rect 25329 10081 25363 10115
rect 2973 10013 3007 10047
rect 3065 10013 3099 10047
rect 4261 10013 4295 10047
rect 4445 10013 4479 10047
rect 8953 10013 8987 10047
rect 12449 10013 12483 10047
rect 18981 10013 19015 10047
rect 23213 10013 23247 10047
rect 2881 9945 2915 9979
rect 3801 9945 3835 9979
rect 5273 9945 5307 9979
rect 8769 9945 8803 9979
rect 11713 9945 11747 9979
rect 13921 9945 13955 9979
rect 20361 9945 20395 9979
rect 2237 9877 2271 9911
rect 4721 9877 4755 9911
rect 9689 9877 9723 9911
rect 22661 9877 22695 9911
rect 22845 9877 22879 9911
rect 24777 9877 24811 9911
rect 24869 9877 24903 9911
rect 1869 9673 1903 9707
rect 3065 9673 3099 9707
rect 8217 9673 8251 9707
rect 21741 9673 21775 9707
rect 22937 9673 22971 9707
rect 25605 9673 25639 9707
rect 3249 9605 3283 9639
rect 3985 9605 4019 9639
rect 7205 9605 7239 9639
rect 8677 9605 8711 9639
rect 15853 9605 15887 9639
rect 19349 9605 19383 9639
rect 21373 9605 21407 9639
rect 21465 9605 21499 9639
rect 1961 9537 1995 9571
rect 2513 9537 2547 9571
rect 4169 9537 4203 9571
rect 5273 9537 5307 9571
rect 6561 9537 6595 9571
rect 7113 9537 7147 9571
rect 14013 9537 14047 9571
rect 24593 9537 24627 9571
rect 1593 9469 1627 9503
rect 2789 9469 2823 9503
rect 2881 9469 2915 9503
rect 3801 9469 3835 9503
rect 4261 9469 4295 9503
rect 4353 9469 4387 9503
rect 4445 9469 4479 9503
rect 5089 9469 5123 9503
rect 5181 9469 5215 9503
rect 5365 9469 5399 9503
rect 6101 9469 6135 9503
rect 6193 9469 6227 9503
rect 6377 9469 6411 9503
rect 6837 9469 6871 9503
rect 7021 9469 7055 9503
rect 7297 9469 7331 9503
rect 7481 9469 7515 9503
rect 7573 9469 7607 9503
rect 8585 9469 8619 9503
rect 8769 9469 8803 9503
rect 8861 9469 8895 9503
rect 9045 9469 9079 9503
rect 9321 9469 9355 9503
rect 9781 9469 9815 9503
rect 11529 9469 11563 9503
rect 11677 9469 11711 9503
rect 12035 9469 12069 9503
rect 12357 9469 12391 9503
rect 17233 9469 17267 9503
rect 17969 9469 18003 9503
rect 18981 9469 19015 9503
rect 19528 9469 19562 9503
rect 19900 9469 19934 9503
rect 19993 9469 20027 9503
rect 21281 9469 21315 9503
rect 21557 9469 21591 9503
rect 22017 9469 22051 9503
rect 22201 9469 22235 9503
rect 22385 9469 22419 9503
rect 22477 9469 22511 9503
rect 22937 9469 22971 9503
rect 23121 9469 23155 9503
rect 23857 9469 23891 9503
rect 24015 9469 24049 9503
rect 24133 9469 24167 9503
rect 24317 9469 24351 9503
rect 24501 9469 24535 9503
rect 24777 9469 24811 9503
rect 25053 9469 25087 9503
rect 25329 9469 25363 9503
rect 25697 9469 25731 9503
rect 25789 9469 25823 9503
rect 1869 9401 1903 9435
rect 3065 9401 3099 9435
rect 5733 9401 5767 9435
rect 5917 9401 5951 9435
rect 9505 9401 9539 9435
rect 11805 9401 11839 9435
rect 11897 9401 11931 9435
rect 15761 9401 15795 9435
rect 16966 9401 17000 9435
rect 19625 9401 19659 9435
rect 19717 9401 19751 9435
rect 24225 9401 24259 9435
rect 25881 9401 25915 9435
rect 1685 9333 1719 9367
rect 4905 9333 4939 9367
rect 5549 9333 5583 9367
rect 5825 9333 5859 9367
rect 8401 9333 8435 9367
rect 9137 9333 9171 9367
rect 10425 9333 10459 9367
rect 12173 9333 12207 9367
rect 12909 9333 12943 9367
rect 17785 9333 17819 9367
rect 18797 9333 18831 9367
rect 24961 9333 24995 9367
rect 25145 9333 25179 9367
rect 2881 9129 2915 9163
rect 5641 9129 5675 9163
rect 6561 9129 6595 9163
rect 9597 9129 9631 9163
rect 9689 9129 9723 9163
rect 12357 9129 12391 9163
rect 12633 9129 12667 9163
rect 13461 9129 13495 9163
rect 16865 9129 16899 9163
rect 1768 9061 1802 9095
rect 9873 9061 9907 9095
rect 10057 9061 10091 9095
rect 14197 9061 14231 9095
rect 14534 9061 14568 9095
rect 16497 9061 16531 9095
rect 26433 9061 26467 9095
rect 4528 8993 4562 9027
rect 6377 8993 6411 9027
rect 7481 8993 7515 9027
rect 7665 8993 7699 9027
rect 7849 8993 7883 9027
rect 7941 8993 7975 9027
rect 8217 8993 8251 9027
rect 8484 8993 8518 9027
rect 11244 8993 11278 9027
rect 12449 8993 12483 9027
rect 13553 8993 13587 9027
rect 13737 8993 13771 9027
rect 13829 8993 13863 9027
rect 13921 8993 13955 9027
rect 14289 8993 14323 9027
rect 16129 8993 16163 9027
rect 16222 8993 16256 9027
rect 16405 8993 16439 9027
rect 16635 8993 16669 9027
rect 17141 8993 17175 9027
rect 17233 8993 17267 9027
rect 17325 8993 17359 9027
rect 17509 8993 17543 9027
rect 17601 8993 17635 9027
rect 17969 8993 18003 9027
rect 18337 8993 18371 9027
rect 18521 8993 18555 9027
rect 19625 8993 19659 9027
rect 19809 8993 19843 9027
rect 20361 8993 20395 9027
rect 20453 8993 20487 9027
rect 23673 8993 23707 9027
rect 24685 8993 24719 9027
rect 24777 8993 24811 9027
rect 25053 8993 25087 9027
rect 25145 8993 25179 9027
rect 25329 8993 25363 9027
rect 25421 8993 25455 9027
rect 25513 8993 25547 9027
rect 25881 8993 25915 9027
rect 26065 8993 26099 9027
rect 26157 8993 26191 9027
rect 1501 8925 1535 8959
rect 4261 8925 4295 8959
rect 6193 8925 6227 8959
rect 10977 8925 11011 8959
rect 12817 8925 12851 8959
rect 19993 8925 20027 8959
rect 24133 8925 24167 8959
rect 24593 8925 24627 8959
rect 26985 8925 27019 8959
rect 7757 8857 7791 8891
rect 15669 8857 15703 8891
rect 16773 8857 16807 8891
rect 17785 8857 17819 8891
rect 18429 8857 18463 8891
rect 20177 8857 20211 8891
rect 24869 8857 24903 8891
rect 8125 8789 8159 8823
rect 18153 8789 18187 8823
rect 20637 8789 20671 8823
rect 23949 8789 23983 8823
rect 24317 8789 24351 8823
rect 24685 8789 24719 8823
rect 24777 8789 24811 8823
rect 25789 8789 25823 8823
rect 25881 8789 25915 8823
rect 4997 8585 5031 8619
rect 7021 8585 7055 8619
rect 7849 8585 7883 8619
rect 11253 8585 11287 8619
rect 13553 8585 13587 8619
rect 14197 8585 14231 8619
rect 17325 8585 17359 8619
rect 20085 8585 20119 8619
rect 21649 8585 21683 8619
rect 3341 8517 3375 8551
rect 4629 8517 4663 8551
rect 5181 8517 5215 8551
rect 11621 8517 11655 8551
rect 3525 8449 3559 8483
rect 4261 8449 4295 8483
rect 13369 8449 13403 8483
rect 15577 8449 15611 8483
rect 18705 8449 18739 8483
rect 23857 8449 23891 8483
rect 3249 8381 3283 8415
rect 4353 8381 4387 8415
rect 4537 8381 4571 8415
rect 5457 8381 5491 8415
rect 5917 8381 5951 8415
rect 6469 8381 6503 8415
rect 6653 8381 6687 8415
rect 6837 8381 6871 8415
rect 7481 8381 7515 8415
rect 7665 8381 7699 8415
rect 8401 8381 8435 8415
rect 11437 8381 11471 8415
rect 11529 8381 11563 8415
rect 11713 8381 11747 8415
rect 11897 8381 11931 8415
rect 11989 8381 12023 8415
rect 12082 8381 12116 8415
rect 12454 8381 12488 8415
rect 12749 8381 12783 8415
rect 12909 8381 12943 8415
rect 13001 8381 13035 8415
rect 13139 8381 13173 8415
rect 15310 8381 15344 8415
rect 17141 8381 17175 8415
rect 17785 8381 17819 8415
rect 17969 8381 18003 8415
rect 18061 8381 18095 8415
rect 18153 8381 18187 8415
rect 20269 8381 20303 8415
rect 22293 8381 22327 8415
rect 23029 8381 23063 8415
rect 25513 8381 25547 8415
rect 25780 8381 25814 8415
rect 3617 8313 3651 8347
rect 4997 8313 5031 8347
rect 8646 8313 8680 8347
rect 12265 8313 12299 8347
rect 12357 8313 12391 8347
rect 13737 8313 13771 8347
rect 13921 8313 13955 8347
rect 18429 8313 18463 8347
rect 18950 8313 18984 8347
rect 20536 8313 20570 8347
rect 21741 8313 21775 8347
rect 24102 8313 24136 8347
rect 3525 8245 3559 8279
rect 4445 8245 4479 8279
rect 5273 8245 5307 8279
rect 9781 8245 9815 8279
rect 12633 8245 12667 8279
rect 22477 8245 22511 8279
rect 25237 8245 25271 8279
rect 26893 8245 26927 8279
rect 4261 8041 4295 8075
rect 6193 8041 6227 8075
rect 6469 8041 6503 8075
rect 19165 8041 19199 8075
rect 21097 8041 21131 8075
rect 23673 8041 23707 8075
rect 2228 7973 2262 8007
rect 3525 7973 3559 8007
rect 4413 7973 4447 8007
rect 4629 7973 4663 8007
rect 6101 7973 6135 8007
rect 8953 7973 8987 8007
rect 9321 7973 9355 8007
rect 11713 7973 11747 8007
rect 24225 7973 24259 8007
rect 26617 7973 26651 8007
rect 1961 7905 1995 7939
rect 3433 7905 3467 7939
rect 3617 7905 3651 7939
rect 3893 7905 3927 7939
rect 4077 7905 4111 7939
rect 4813 7905 4847 7939
rect 6009 7905 6043 7939
rect 8861 7905 8895 7939
rect 9137 7905 9171 7939
rect 9413 7905 9447 7939
rect 9597 7905 9631 7939
rect 9689 7905 9723 7939
rect 9781 7905 9815 7939
rect 10149 7905 10183 7939
rect 10793 7905 10827 7939
rect 11345 7905 11379 7939
rect 11493 7905 11527 7939
rect 11621 7905 11655 7939
rect 11851 7905 11885 7939
rect 12348 7905 12382 7939
rect 13553 7905 13587 7939
rect 13701 7905 13735 7939
rect 13829 7905 13863 7939
rect 13921 7905 13955 7939
rect 14018 7905 14052 7939
rect 14295 7905 14329 7939
rect 14473 7905 14507 7939
rect 14565 7905 14599 7939
rect 14657 7905 14691 7939
rect 16129 7905 16163 7939
rect 17417 7905 17451 7939
rect 19809 7905 19843 7939
rect 19901 7905 19935 7939
rect 20453 7905 20487 7939
rect 20637 7905 20671 7939
rect 20729 7905 20763 7939
rect 20821 7905 20855 7939
rect 22394 7905 22428 7939
rect 22661 7905 22695 7939
rect 23029 7905 23063 7939
rect 23213 7905 23247 7939
rect 23305 7905 23339 7939
rect 23397 7905 23431 7939
rect 24317 7905 24351 7939
rect 24961 7905 24995 7939
rect 25329 7905 25363 7939
rect 25605 7905 25639 7939
rect 25881 7905 25915 7939
rect 26801 7905 26835 7939
rect 6377 7837 6411 7871
rect 7021 7837 7055 7871
rect 12081 7837 12115 7871
rect 14933 7837 14967 7871
rect 15577 7837 15611 7871
rect 16681 7837 16715 7871
rect 24409 7837 24443 7871
rect 25421 7837 25455 7871
rect 26157 7837 26191 7871
rect 3709 7769 3743 7803
rect 14197 7769 14231 7803
rect 17601 7769 17635 7803
rect 21281 7769 21315 7803
rect 26433 7769 26467 7803
rect 3341 7701 3375 7735
rect 4445 7701 4479 7735
rect 5365 7701 5399 7735
rect 5825 7701 5859 7735
rect 10057 7701 10091 7735
rect 11989 7701 12023 7735
rect 13461 7701 13495 7735
rect 15025 7701 15059 7735
rect 20085 7701 20119 7735
rect 25145 7701 25179 7735
rect 25605 7701 25639 7735
rect 25697 7701 25731 7735
rect 26065 7701 26099 7735
rect 5089 7497 5123 7531
rect 5181 7497 5215 7531
rect 5549 7497 5583 7531
rect 7205 7497 7239 7531
rect 12357 7497 12391 7531
rect 15945 7497 15979 7531
rect 20913 7497 20947 7531
rect 23857 7497 23891 7531
rect 24409 7497 24443 7531
rect 26065 7497 26099 7531
rect 4905 7429 4939 7463
rect 11345 7429 11379 7463
rect 16681 7429 16715 7463
rect 20085 7429 20119 7463
rect 22477 7429 22511 7463
rect 4997 7361 5031 7395
rect 5365 7361 5399 7395
rect 9137 7361 9171 7395
rect 9229 7361 9263 7395
rect 11989 7361 12023 7395
rect 13553 7361 13587 7395
rect 20729 7361 20763 7395
rect 3525 7293 3559 7327
rect 5273 7293 5307 7327
rect 5641 7293 5675 7327
rect 5825 7293 5859 7327
rect 8493 7293 8527 7327
rect 8677 7293 8711 7327
rect 8769 7293 8803 7327
rect 8861 7293 8895 7327
rect 9965 7293 9999 7327
rect 12909 7293 12943 7327
rect 13093 7293 13127 7327
rect 14565 7293 14599 7327
rect 14832 7293 14866 7327
rect 16037 7293 16071 7327
rect 16130 7293 16164 7327
rect 16543 7293 16577 7327
rect 16773 7293 16807 7327
rect 17693 7293 17727 7327
rect 17877 7293 17911 7327
rect 17969 7293 18003 7327
rect 18061 7293 18095 7327
rect 18705 7293 18739 7327
rect 20177 7293 20211 7327
rect 21092 7293 21126 7327
rect 21189 7293 21223 7327
rect 21281 7293 21315 7327
rect 21464 7293 21498 7327
rect 21557 7293 21591 7327
rect 21649 7293 21683 7327
rect 22661 7293 22695 7327
rect 24038 7293 24072 7327
rect 24501 7293 24535 7327
rect 24869 7293 24903 7327
rect 24961 7293 24995 7327
rect 25053 7293 25087 7327
rect 25237 7293 25271 7327
rect 25881 7293 25915 7327
rect 26617 7293 26651 7327
rect 3792 7225 3826 7259
rect 6070 7225 6104 7259
rect 9873 7225 9907 7259
rect 10210 7225 10244 7259
rect 14197 7225 14231 7259
rect 16313 7225 16347 7259
rect 16405 7225 16439 7259
rect 18972 7225 19006 7259
rect 22293 7225 22327 7259
rect 25329 7225 25363 7259
rect 5365 7157 5399 7191
rect 11437 7157 11471 7191
rect 13277 7157 13311 7191
rect 16957 7157 16991 7191
rect 18337 7157 18371 7191
rect 24041 7157 24075 7191
rect 24593 7157 24627 7191
rect 5917 6953 5951 6987
rect 8677 6953 8711 6987
rect 10793 6953 10827 6987
rect 15945 6953 15979 6987
rect 21281 6953 21315 6987
rect 25697 6953 25731 6987
rect 26249 6953 26283 6987
rect 24584 6885 24618 6919
rect 5457 6817 5491 6851
rect 5641 6817 5675 6851
rect 5825 6817 5859 6851
rect 6009 6817 6043 6851
rect 8125 6817 8159 6851
rect 8861 6817 8895 6851
rect 9045 6817 9079 6851
rect 9137 6817 9171 6851
rect 9413 6817 9447 6851
rect 9680 6817 9714 6851
rect 11897 6817 11931 6851
rect 11989 6817 12023 6851
rect 12173 6817 12207 6851
rect 12541 6817 12575 6851
rect 12633 6817 12667 6851
rect 12725 6817 12759 6851
rect 12909 6817 12943 6851
rect 13737 6817 13771 6851
rect 13829 6817 13863 6851
rect 14013 6817 14047 6851
rect 14197 6817 14231 6851
rect 14832 6817 14866 6851
rect 16681 6817 16715 6851
rect 17785 6817 17819 6851
rect 17877 6817 17911 6851
rect 18133 6817 18167 6851
rect 19349 6817 19383 6851
rect 19901 6817 19935 6851
rect 21097 6817 21131 6851
rect 22405 6817 22439 6851
rect 22753 6817 22787 6851
rect 25881 6817 25915 6851
rect 26065 6817 26099 6851
rect 26433 6817 26467 6851
rect 11713 6749 11747 6783
rect 12265 6749 12299 6783
rect 13553 6749 13587 6783
rect 14565 6749 14599 6783
rect 17233 6749 17267 6783
rect 20729 6749 20763 6783
rect 22661 6749 22695 6783
rect 23305 6749 23339 6783
rect 24317 6749 24351 6783
rect 25789 6749 25823 6783
rect 26985 6749 27019 6783
rect 12173 6681 12207 6715
rect 19257 6681 19291 6715
rect 20913 6681 20947 6715
rect 5457 6613 5491 6647
rect 6837 6613 6871 6647
rect 11161 6613 11195 6647
rect 13001 6613 13035 6647
rect 16129 6613 16163 6647
rect 20085 6613 20119 6647
rect 5549 6409 5583 6443
rect 6469 6409 6503 6443
rect 6653 6409 6687 6443
rect 7113 6409 7147 6443
rect 14933 6409 14967 6443
rect 18705 6409 18739 6443
rect 22477 6409 22511 6443
rect 25973 6409 26007 6443
rect 5457 6341 5491 6375
rect 7021 6341 7055 6375
rect 12357 6341 12391 6375
rect 5641 6273 5675 6307
rect 6101 6273 6135 6307
rect 8861 6273 8895 6307
rect 12909 6273 12943 6307
rect 21005 6273 21039 6307
rect 24593 6273 24627 6307
rect 4721 6205 4755 6239
rect 5273 6205 5307 6239
rect 5365 6205 5399 6239
rect 5917 6205 5951 6239
rect 6009 6205 6043 6239
rect 6193 6205 6227 6239
rect 7297 6205 7331 6239
rect 7481 6205 7515 6239
rect 7573 6205 7607 6239
rect 7757 6205 7791 6239
rect 8677 6205 8711 6239
rect 9413 6205 9447 6239
rect 9505 6205 9539 6239
rect 9873 6205 9907 6239
rect 11897 6205 11931 6239
rect 11989 6205 12023 6239
rect 12081 6205 12115 6239
rect 12173 6205 12207 6239
rect 14381 6205 14415 6239
rect 14657 6205 14691 6239
rect 15485 6205 15519 6239
rect 15761 6205 15795 6239
rect 17877 6205 17911 6239
rect 18245 6205 18279 6239
rect 18981 6205 19015 6239
rect 19073 6205 19107 6239
rect 19165 6205 19199 6239
rect 19349 6205 19383 6239
rect 21649 6205 21683 6239
rect 21833 6205 21867 6239
rect 21996 6205 22030 6239
rect 22112 6205 22146 6239
rect 22247 6205 22281 6239
rect 22845 6205 22879 6239
rect 23581 6205 23615 6239
rect 24409 6205 24443 6239
rect 24860 6205 24894 6239
rect 6653 6137 6687 6171
rect 7849 6137 7883 6171
rect 8033 6137 8067 6171
rect 14473 6137 14507 6171
rect 16028 6137 16062 6171
rect 20760 6137 20794 6171
rect 21097 6137 21131 6171
rect 6377 6069 6411 6103
rect 7757 6069 7791 6103
rect 8217 6069 8251 6103
rect 8493 6069 8527 6103
rect 9597 6069 9631 6103
rect 11161 6069 11195 6103
rect 11713 6069 11747 6103
rect 14841 6069 14875 6103
rect 17141 6069 17175 6103
rect 17233 6069 17267 6103
rect 18429 6069 18463 6103
rect 19625 6069 19659 6103
rect 22661 6069 22695 6103
rect 23397 6069 23431 6103
rect 23857 6069 23891 6103
rect 4261 5865 4295 5899
rect 6377 5865 6411 5899
rect 6469 5865 6503 5899
rect 8217 5865 8251 5899
rect 10149 5865 10183 5899
rect 13093 5865 13127 5899
rect 14933 5865 14967 5899
rect 16129 5865 16163 5899
rect 21925 5865 21959 5899
rect 23397 5865 23431 5899
rect 14105 5797 14139 5831
rect 19625 5797 19659 5831
rect 5374 5729 5408 5763
rect 6009 5729 6043 5763
rect 6285 5729 6319 5763
rect 7104 5729 7138 5763
rect 8309 5729 8343 5763
rect 8576 5729 8610 5763
rect 9873 5729 9907 5763
rect 10977 5729 11011 5763
rect 11161 5729 11195 5763
rect 11253 5729 11287 5763
rect 11437 5729 11471 5763
rect 11529 5729 11563 5763
rect 11621 5729 11655 5763
rect 11877 5729 11911 5763
rect 13829 5729 13863 5763
rect 14381 5729 14415 5763
rect 14473 5729 14507 5763
rect 14657 5729 14691 5763
rect 15209 5729 15243 5763
rect 15301 5729 15335 5763
rect 15393 5729 15427 5763
rect 15577 5729 15611 5763
rect 17141 5729 17175 5763
rect 17233 5729 17267 5763
rect 17325 5729 17359 5763
rect 17509 5729 17543 5763
rect 17877 5729 17911 5763
rect 18061 5729 18095 5763
rect 18153 5729 18187 5763
rect 18245 5729 18279 5763
rect 18889 5729 18923 5763
rect 18982 5729 19016 5763
rect 19165 5729 19199 5763
rect 19257 5729 19291 5763
rect 19395 5729 19429 5763
rect 20361 5729 20395 5763
rect 21281 5729 21315 5763
rect 21429 5729 21463 5763
rect 21557 5729 21591 5763
rect 21649 5729 21683 5763
rect 21787 5729 21821 5763
rect 22005 5729 22039 5763
rect 22385 5729 22419 5763
rect 22533 5729 22567 5763
rect 22661 5729 22695 5763
rect 22753 5729 22787 5763
rect 22891 5729 22925 5763
rect 24521 5729 24555 5763
rect 24777 5729 24811 5763
rect 5641 5661 5675 5695
rect 6837 5661 6871 5695
rect 11069 5661 11103 5695
rect 13645 5661 13679 5695
rect 14105 5661 14139 5695
rect 16773 5661 16807 5695
rect 16865 5661 16899 5695
rect 20177 5661 20211 5695
rect 24869 5661 24903 5695
rect 25421 5661 25455 5695
rect 6653 5593 6687 5627
rect 11253 5593 11287 5627
rect 13921 5593 13955 5627
rect 14841 5593 14875 5627
rect 19533 5593 19567 5627
rect 5825 5525 5859 5559
rect 6101 5525 6135 5559
rect 9689 5525 9723 5559
rect 13001 5525 13035 5559
rect 18521 5525 18555 5559
rect 21005 5525 21039 5559
rect 22201 5525 22235 5559
rect 23029 5525 23063 5559
rect 6009 5321 6043 5355
rect 7389 5321 7423 5355
rect 8585 5321 8619 5355
rect 8769 5321 8803 5355
rect 11345 5321 11379 5355
rect 14749 5321 14783 5355
rect 20085 5321 20119 5355
rect 20821 5321 20855 5355
rect 23581 5321 23615 5355
rect 22385 5253 22419 5287
rect 23857 5253 23891 5287
rect 9229 5185 9263 5219
rect 13553 5185 13587 5219
rect 4629 5117 4663 5151
rect 4896 5117 4930 5151
rect 7941 5117 7975 5151
rect 9045 5117 9079 5151
rect 12725 5117 12759 5151
rect 14289 5117 14323 5151
rect 14565 5117 14599 5151
rect 14841 5117 14875 5151
rect 15945 5117 15979 5151
rect 16497 5117 16531 5151
rect 17141 5117 17175 5151
rect 18705 5117 18739 5151
rect 20177 5117 20211 5151
rect 20361 5117 20395 5151
rect 20453 5117 20487 5151
rect 20545 5117 20579 5151
rect 21097 5117 21131 5151
rect 22937 5117 22971 5151
rect 23121 5117 23155 5151
rect 23213 5117 23247 5151
rect 23305 5117 23339 5151
rect 25237 5117 25271 5151
rect 25881 5117 25915 5151
rect 8401 5049 8435 5083
rect 8861 5049 8895 5083
rect 12458 5049 12492 5083
rect 17049 5049 17083 5083
rect 17386 5049 17420 5083
rect 18972 5049 19006 5083
rect 24992 5049 25026 5083
rect 25329 5049 25363 5083
rect 8601 4981 8635 5015
rect 14197 4981 14231 5015
rect 14381 4981 14415 5015
rect 15025 4981 15059 5015
rect 16129 4981 16163 5015
rect 18521 4981 18555 5015
rect 7573 4777 7607 4811
rect 13001 4777 13035 4811
rect 24133 4777 24167 4811
rect 8125 4709 8159 4743
rect 11345 4709 11379 4743
rect 13553 4709 13587 4743
rect 19441 4709 19475 4743
rect 20545 4709 20579 4743
rect 5273 4641 5307 4675
rect 5457 4641 5491 4675
rect 6101 4641 6135 4675
rect 6285 4641 6319 4675
rect 7389 4641 7423 4675
rect 7481 4641 7515 4675
rect 7665 4641 7699 4675
rect 7757 4641 7791 4675
rect 7849 4641 7883 4675
rect 8309 4641 8343 4675
rect 8585 4641 8619 4675
rect 8769 4641 8803 4675
rect 9045 4641 9079 4675
rect 12541 4641 12575 4675
rect 12633 4641 12667 4675
rect 12817 4641 12851 4675
rect 13093 4641 13127 4675
rect 13185 4641 13219 4675
rect 13369 4641 13403 4675
rect 14013 4641 14047 4675
rect 14105 4641 14139 4675
rect 14289 4641 14323 4675
rect 14832 4641 14866 4675
rect 16129 4641 16163 4675
rect 17141 4641 17175 4675
rect 17233 4641 17267 4675
rect 17325 4641 17359 4675
rect 17509 4641 17543 4675
rect 20085 4641 20119 4675
rect 20269 4641 20303 4675
rect 20362 4641 20396 4675
rect 20637 4641 20671 4675
rect 20775 4641 20809 4675
rect 22293 4641 22327 4675
rect 22385 4641 22419 4675
rect 22477 4641 22511 4675
rect 22661 4641 22695 4675
rect 23489 4641 23523 4675
rect 23673 4641 23707 4675
rect 23765 4641 23799 4675
rect 23857 4641 23891 4675
rect 24225 4641 24259 4675
rect 24777 4641 24811 4675
rect 6469 4573 6503 4607
rect 10149 4573 10183 4607
rect 10793 4573 10827 4607
rect 14565 4573 14599 4607
rect 16773 4573 16807 4607
rect 16865 4573 16899 4607
rect 19533 4573 19567 4607
rect 21925 4573 21959 4607
rect 22017 4573 22051 4607
rect 22753 4573 22787 4607
rect 11713 4505 11747 4539
rect 15945 4505 15979 4539
rect 20913 4505 20947 4539
rect 5273 4437 5307 4471
rect 8493 4437 8527 4471
rect 8677 4437 8711 4471
rect 9229 4437 9263 4471
rect 11161 4437 11195 4471
rect 11345 4437 11379 4471
rect 14473 4437 14507 4471
rect 18153 4437 18187 4471
rect 21281 4437 21315 4471
rect 23397 4437 23431 4471
rect 8585 4233 8619 4267
rect 8769 4233 8803 4267
rect 10425 4233 10459 4267
rect 12449 4233 12483 4267
rect 14841 4233 14875 4267
rect 22201 4233 22235 4267
rect 23305 4233 23339 4267
rect 6009 4165 6043 4199
rect 8125 4165 8159 4199
rect 7941 4097 7975 4131
rect 20821 4097 20855 4131
rect 4629 4029 4663 4063
rect 6469 4029 6503 4063
rect 7297 4029 7331 4063
rect 7665 4029 7699 4063
rect 8217 4029 8251 4063
rect 9045 4029 9079 4063
rect 9312 4029 9346 4063
rect 10793 4029 10827 4063
rect 11069 4029 11103 4063
rect 12725 4029 12759 4063
rect 13553 4029 13587 4063
rect 14105 4029 14139 4063
rect 14289 4029 14323 4063
rect 14565 4029 14599 4063
rect 15117 4029 15151 4063
rect 15209 4029 15243 4063
rect 15301 4029 15335 4063
rect 15485 4029 15519 4063
rect 15945 4029 15979 4063
rect 16129 4029 16163 4063
rect 16221 4029 16255 4063
rect 16313 4029 16347 4063
rect 16681 4029 16715 4063
rect 18981 4029 19015 4063
rect 21088 4029 21122 4063
rect 22385 4029 22419 4063
rect 22533 4029 22567 4063
rect 22850 4029 22884 4063
rect 23121 4029 23155 4063
rect 23995 4029 24029 4063
rect 24133 4029 24167 4063
rect 24225 4029 24259 4063
rect 24353 4029 24387 4063
rect 24501 4029 24535 4063
rect 25145 4029 25179 4063
rect 4896 3961 4930 3995
rect 7849 3961 7883 3995
rect 8401 3961 8435 3995
rect 11314 3961 11348 3995
rect 14381 3961 14415 3995
rect 14749 3961 14783 3995
rect 16948 3961 16982 3995
rect 19226 3961 19260 3995
rect 22661 3961 22695 3995
rect 22753 3961 22787 3995
rect 7113 3893 7147 3927
rect 7481 3893 7515 3927
rect 7573 3893 7607 3927
rect 7941 3893 7975 3927
rect 8601 3893 8635 3927
rect 10977 3893 11011 3927
rect 12633 3893 12667 3927
rect 16589 3893 16623 3927
rect 18061 3893 18095 3927
rect 20361 3893 20395 3927
rect 23029 3893 23063 3927
rect 23857 3893 23891 3927
rect 24593 3893 24627 3927
rect 5365 3689 5399 3723
rect 8309 3689 8343 3723
rect 17601 3689 17635 3723
rect 19073 3689 19107 3723
rect 22661 3689 22695 3723
rect 25605 3689 25639 3723
rect 7104 3621 7138 3655
rect 13185 3621 13219 3655
rect 13277 3621 13311 3655
rect 15209 3621 15243 3655
rect 23888 3621 23922 3655
rect 5549 3553 5583 3587
rect 5641 3553 5675 3587
rect 5825 3553 5859 3587
rect 6469 3553 6503 3587
rect 8953 3553 8987 3587
rect 9965 3553 9999 3587
rect 11529 3553 11563 3587
rect 11796 3553 11830 3587
rect 13093 3553 13127 3587
rect 13461 3553 13495 3587
rect 13553 3553 13587 3587
rect 14749 3553 14783 3587
rect 14841 3553 14875 3587
rect 15025 3553 15059 3587
rect 15301 3553 15335 3587
rect 15485 3553 15519 3587
rect 15577 3553 15611 3587
rect 15669 3553 15703 3587
rect 16129 3553 16163 3587
rect 16385 3553 16419 3587
rect 18153 3553 18187 3587
rect 18429 3553 18463 3587
rect 18613 3553 18647 3587
rect 18705 3553 18739 3587
rect 18797 3553 18831 3587
rect 19625 3553 19659 3587
rect 20269 3553 20303 3587
rect 21557 3553 21591 3587
rect 21649 3553 21683 3587
rect 21741 3553 21775 3587
rect 21925 3553 21959 3587
rect 22017 3553 22051 3587
rect 22201 3553 22235 3587
rect 22293 3553 22327 3587
rect 22385 3553 22419 3587
rect 24492 3553 24526 3587
rect 5365 3485 5399 3519
rect 6837 3485 6871 3519
rect 9045 3485 9079 3519
rect 10149 3485 10183 3519
rect 13001 3485 13035 3519
rect 15945 3485 15979 3519
rect 21005 3485 21039 3519
rect 21281 3485 21315 3519
rect 24133 3485 24167 3519
rect 24225 3485 24259 3519
rect 8217 3417 8251 3451
rect 9689 3417 9723 3451
rect 22753 3417 22787 3451
rect 9781 3349 9815 3383
rect 12909 3349 12943 3383
rect 17509 3349 17543 3383
rect 20361 3349 20395 3383
rect 6377 3145 6411 3179
rect 8953 3145 8987 3179
rect 11805 3145 11839 3179
rect 12449 3145 12483 3179
rect 16681 3145 16715 3179
rect 17417 3145 17451 3179
rect 21373 3145 21407 3179
rect 22661 3145 22695 3179
rect 24593 3145 24627 3179
rect 8217 3077 8251 3111
rect 11621 3077 11655 3111
rect 13185 3077 13219 3111
rect 21281 3077 21315 3111
rect 6377 3009 6411 3043
rect 6837 3009 6871 3043
rect 12357 3009 12391 3043
rect 12909 3009 12943 3043
rect 13369 3009 13403 3043
rect 17325 3009 17359 3043
rect 21925 3009 21959 3043
rect 24501 3009 24535 3043
rect 25145 3009 25179 3043
rect 25881 3009 25915 3043
rect 6469 2941 6503 2975
rect 6653 2941 6687 2975
rect 8493 2941 8527 2975
rect 8585 2941 8619 2975
rect 11345 2941 11379 2975
rect 11437 2941 11471 2975
rect 11989 2941 12023 2975
rect 12633 2941 12667 2975
rect 12725 2941 12759 2975
rect 12817 2941 12851 2975
rect 13093 2941 13127 2975
rect 17969 2941 18003 2975
rect 18429 2941 18463 2975
rect 18705 2941 18739 2975
rect 19901 2941 19935 2975
rect 23213 2941 23247 2975
rect 23857 2941 23891 2975
rect 24041 2941 24075 2975
rect 24133 2941 24167 2975
rect 24225 2941 24259 2975
rect 25329 2941 25363 2975
rect 6745 2873 6779 2907
rect 7104 2873 7138 2907
rect 8921 2873 8955 2907
rect 9137 2873 9171 2907
rect 12081 2873 12115 2907
rect 20168 2873 20202 2907
rect 8769 2805 8803 2839
rect 12173 2805 12207 2839
rect 13369 2805 13403 2839
rect 18245 2805 18279 2839
rect 19349 2805 19383 2839
rect 7573 2601 7607 2635
rect 11345 2601 11379 2635
rect 11989 2601 12023 2635
rect 14841 2601 14875 2635
rect 19901 2601 19935 2635
rect 21281 2601 21315 2635
rect 23397 2601 23431 2635
rect 9965 2533 9999 2567
rect 12541 2533 12575 2567
rect 13521 2533 13555 2567
rect 13737 2533 13771 2567
rect 13829 2533 13863 2567
rect 18788 2533 18822 2567
rect 23121 2533 23155 2567
rect 26065 2533 26099 2567
rect 7481 2465 7515 2499
rect 7665 2465 7699 2499
rect 9781 2465 9815 2499
rect 10057 2465 10091 2499
rect 10241 2465 10275 2499
rect 10425 2465 10459 2499
rect 11069 2465 11103 2499
rect 11253 2465 11287 2499
rect 11529 2465 11563 2499
rect 11805 2465 11839 2499
rect 12173 2465 12207 2499
rect 12265 2465 12299 2499
rect 12357 2465 12391 2499
rect 14013 2465 14047 2499
rect 14105 2465 14139 2499
rect 14749 2465 14783 2499
rect 15025 2465 15059 2499
rect 15301 2465 15335 2499
rect 15393 2465 15427 2499
rect 15577 2465 15611 2499
rect 17141 2465 17175 2499
rect 17233 2465 17267 2499
rect 17325 2465 17359 2499
rect 17509 2465 17543 2499
rect 20637 2465 20671 2499
rect 21460 2465 21494 2499
rect 21557 2465 21591 2499
rect 21649 2465 21683 2499
rect 21832 2465 21866 2499
rect 21925 2465 21959 2499
rect 22196 2465 22230 2499
rect 22293 2465 22327 2499
rect 22385 2465 22419 2499
rect 22513 2465 22547 2499
rect 22661 2465 22695 2499
rect 22753 2465 22787 2499
rect 22901 2465 22935 2499
rect 23029 2465 23063 2499
rect 23218 2465 23252 2499
rect 24216 2465 24250 2499
rect 26433 2465 26467 2499
rect 10517 2397 10551 2431
rect 11161 2397 11195 2431
rect 11621 2397 11655 2431
rect 11713 2397 11747 2431
rect 13277 2397 13311 2431
rect 16681 2397 16715 2431
rect 17601 2397 17635 2431
rect 18245 2397 18279 2431
rect 18521 2397 18555 2431
rect 23949 2397 23983 2431
rect 25421 2397 25455 2431
rect 26985 2397 27019 2431
rect 12633 2329 12667 2363
rect 15761 2329 15795 2363
rect 25329 2329 25363 2363
rect 9597 2261 9631 2295
rect 10149 2261 10183 2295
rect 10425 2261 10459 2295
rect 10793 2261 10827 2295
rect 13369 2261 13403 2295
rect 13553 2261 13587 2295
rect 13829 2261 13863 2295
rect 15209 2261 15243 2295
rect 16129 2261 16163 2295
rect 16865 2261 16899 2295
rect 19993 2261 20027 2295
rect 22017 2261 22051 2295
rect 9689 2057 9723 2091
rect 10241 2057 10275 2091
rect 11253 2057 11287 2091
rect 14289 2057 14323 2091
rect 15577 2057 15611 2091
rect 18521 2057 18555 2091
rect 25973 2057 26007 2091
rect 10333 1989 10367 2023
rect 17049 1989 17083 2023
rect 21465 1989 21499 2023
rect 25237 1989 25271 2023
rect 10425 1921 10459 1955
rect 13369 1921 13403 1955
rect 15669 1921 15703 1955
rect 17785 1921 17819 1955
rect 20085 1921 20119 1955
rect 22201 1921 22235 1955
rect 23581 1921 23615 1955
rect 9413 1853 9447 1887
rect 9643 1819 9677 1853
rect 10150 1831 10184 1865
rect 10517 1853 10551 1887
rect 10701 1853 10735 1887
rect 10793 1853 10827 1887
rect 10885 1853 10919 1887
rect 11897 1853 11931 1887
rect 13113 1853 13147 1887
rect 13829 1853 13863 1887
rect 14105 1853 14139 1887
rect 14381 1853 14415 1887
rect 14473 1853 14507 1887
rect 14657 1853 14691 1887
rect 14933 1853 14967 1887
rect 15117 1853 15151 1887
rect 15209 1853 15243 1887
rect 15301 1853 15335 1887
rect 15936 1853 15970 1887
rect 17877 1853 17911 1887
rect 18061 1853 18095 1887
rect 18153 1853 18187 1887
rect 18245 1853 18279 1887
rect 18981 1853 19015 1887
rect 19073 1853 19107 1887
rect 19165 1853 19199 1887
rect 19349 1853 19383 1887
rect 21557 1853 21591 1887
rect 22845 1853 22879 1887
rect 23857 1853 23891 1887
rect 23950 1853 23984 1887
rect 24322 1853 24356 1887
rect 24593 1853 24627 1887
rect 24741 1853 24775 1887
rect 24869 1853 24903 1887
rect 24961 1853 24995 1887
rect 25058 1853 25092 1887
rect 25329 1853 25363 1887
rect 25513 1853 25547 1887
rect 25605 1853 25639 1887
rect 25697 1853 25731 1887
rect 26065 1853 26099 1887
rect 26249 1853 26283 1887
rect 26341 1853 26375 1887
rect 26433 1853 26467 1887
rect 9873 1785 9907 1819
rect 17141 1785 17175 1819
rect 20352 1785 20386 1819
rect 22293 1785 22327 1819
rect 24133 1785 24167 1819
rect 24225 1785 24259 1819
rect 9229 1717 9263 1751
rect 9505 1717 9539 1751
rect 11161 1717 11195 1751
rect 11989 1717 12023 1751
rect 13921 1717 13955 1751
rect 14841 1717 14875 1751
rect 18705 1717 18739 1751
rect 23029 1717 23063 1751
rect 24501 1717 24535 1751
rect 26709 1717 26743 1751
rect 10149 1513 10183 1547
rect 14105 1513 14139 1547
rect 20545 1513 20579 1547
rect 23305 1513 23339 1547
rect 24869 1513 24903 1547
rect 9036 1445 9070 1479
rect 16396 1445 16430 1479
rect 24532 1445 24566 1479
rect 25605 1445 25639 1479
rect 11244 1377 11278 1411
rect 12541 1377 12575 1411
rect 12641 1377 12675 1411
rect 12981 1377 13015 1411
rect 14657 1377 14691 1411
rect 14749 1377 14783 1411
rect 14933 1377 14967 1411
rect 16129 1377 16163 1411
rect 18817 1377 18851 1411
rect 19073 1377 19107 1411
rect 19165 1377 19199 1411
rect 19432 1377 19466 1411
rect 22192 1377 22226 1411
rect 26249 1377 26283 1411
rect 8769 1309 8803 1343
rect 10977 1309 11011 1343
rect 12725 1309 12759 1343
rect 21925 1309 21959 1343
rect 24777 1309 24811 1343
rect 25421 1309 25455 1343
rect 12357 1173 12391 1207
rect 15117 1173 15151 1207
rect 17509 1173 17543 1207
rect 17693 1173 17727 1207
rect 23397 1173 23431 1207
rect 12633 969 12667 1003
rect 18521 969 18555 1003
rect 19349 969 19383 1003
rect 20085 969 20119 1003
rect 22201 969 22235 1003
rect 23857 969 23891 1003
rect 25237 969 25271 1003
rect 17877 833 17911 867
rect 18705 833 18739 867
rect 23673 833 23707 867
rect 24409 833 24443 867
rect 12449 765 12483 799
rect 19441 765 19475 799
rect 19625 765 19659 799
rect 19717 765 19751 799
rect 19809 765 19843 799
rect 21557 765 21591 799
rect 21741 765 21775 799
rect 21833 765 21867 799
rect 21925 765 21959 799
rect 22293 765 22327 799
rect 22441 765 22475 799
rect 22569 765 22603 799
rect 22661 765 22695 799
rect 22799 765 22833 799
rect 23029 765 23063 799
rect 23213 765 23247 799
rect 23305 765 23339 799
rect 23397 765 23431 799
rect 24593 765 24627 799
rect 22937 629 22971 663
<< metal1 >>
rect 15470 17728 15476 17740
rect 9646 17700 15476 17728
rect 3602 17484 3608 17536
rect 3660 17524 3666 17536
rect 3970 17524 3976 17536
rect 3660 17496 3976 17524
rect 3660 17484 3666 17496
rect 3970 17484 3976 17496
rect 4028 17484 4034 17536
rect 5626 17484 5632 17536
rect 5684 17524 5690 17536
rect 9646 17524 9674 17700
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 10686 17620 10692 17672
rect 10744 17660 10750 17672
rect 18690 17660 18696 17672
rect 10744 17632 18696 17660
rect 10744 17620 10750 17632
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 9950 17552 9956 17604
rect 10008 17592 10014 17604
rect 16666 17592 16672 17604
rect 10008 17564 16672 17592
rect 10008 17552 10014 17564
rect 16666 17552 16672 17564
rect 16724 17552 16730 17604
rect 5684 17496 9674 17524
rect 5684 17484 5690 17496
rect 10318 17484 10324 17536
rect 10376 17524 10382 17536
rect 23198 17524 23204 17536
rect 10376 17496 23204 17524
rect 10376 17484 10382 17496
rect 23198 17484 23204 17496
rect 23256 17484 23262 17536
rect 23934 17484 23940 17536
rect 23992 17524 23998 17536
rect 24302 17524 24308 17536
rect 23992 17496 24308 17524
rect 23992 17484 23998 17496
rect 24302 17484 24308 17496
rect 24360 17484 24366 17536
rect 552 17434 27416 17456
rect 552 17382 3756 17434
rect 3808 17382 3820 17434
rect 3872 17382 3884 17434
rect 3936 17382 3948 17434
rect 4000 17382 4012 17434
rect 4064 17382 10472 17434
rect 10524 17382 10536 17434
rect 10588 17382 10600 17434
rect 10652 17382 10664 17434
rect 10716 17382 10728 17434
rect 10780 17382 17188 17434
rect 17240 17382 17252 17434
rect 17304 17382 17316 17434
rect 17368 17382 17380 17434
rect 17432 17382 17444 17434
rect 17496 17382 23904 17434
rect 23956 17382 23968 17434
rect 24020 17382 24032 17434
rect 24084 17382 24096 17434
rect 24148 17382 24160 17434
rect 24212 17382 27416 17434
rect 552 17360 27416 17382
rect 2130 17280 2136 17332
rect 2188 17280 2194 17332
rect 2682 17280 2688 17332
rect 2740 17320 2746 17332
rect 2777 17323 2835 17329
rect 2777 17320 2789 17323
rect 2740 17292 2789 17320
rect 2740 17280 2746 17292
rect 2777 17289 2789 17292
rect 2823 17289 2835 17323
rect 2777 17283 2835 17289
rect 3602 17280 3608 17332
rect 3660 17320 3666 17332
rect 4065 17323 4123 17329
rect 4065 17320 4077 17323
rect 3660 17292 4077 17320
rect 3660 17280 3666 17292
rect 4065 17289 4077 17292
rect 4111 17289 4123 17323
rect 4065 17283 4123 17289
rect 7282 17280 7288 17332
rect 7340 17280 7346 17332
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 7929 17323 7987 17329
rect 7929 17320 7941 17323
rect 7892 17292 7941 17320
rect 7892 17280 7898 17292
rect 7929 17289 7941 17292
rect 7975 17289 7987 17323
rect 7929 17283 7987 17289
rect 9122 17280 9128 17332
rect 9180 17320 9186 17332
rect 9309 17323 9367 17329
rect 9309 17320 9321 17323
rect 9180 17292 9321 17320
rect 9180 17280 9186 17292
rect 9309 17289 9321 17292
rect 9355 17289 9367 17323
rect 9309 17283 9367 17289
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 10137 17323 10195 17329
rect 10137 17320 10149 17323
rect 9824 17292 10149 17320
rect 9824 17280 9830 17292
rect 10137 17289 10149 17292
rect 10183 17289 10195 17323
rect 10137 17283 10195 17289
rect 12342 17280 12348 17332
rect 12400 17320 12406 17332
rect 12437 17323 12495 17329
rect 12437 17320 12449 17323
rect 12400 17292 12449 17320
rect 12400 17280 12406 17292
rect 12437 17289 12449 17292
rect 12483 17289 12495 17323
rect 12437 17283 12495 17289
rect 12897 17323 12955 17329
rect 12897 17289 12909 17323
rect 12943 17320 12955 17323
rect 12986 17320 12992 17332
rect 12943 17292 12992 17320
rect 12943 17289 12955 17292
rect 12897 17283 12955 17289
rect 12986 17280 12992 17292
rect 13044 17280 13050 17332
rect 18417 17323 18475 17329
rect 18417 17320 18429 17323
rect 16040 17292 18429 17320
rect 6730 17212 6736 17264
rect 6788 17252 6794 17264
rect 15930 17252 15936 17264
rect 6788 17224 15936 17252
rect 6788 17212 6794 17224
rect 15930 17212 15936 17224
rect 15988 17212 15994 17264
rect 3418 17144 3424 17196
rect 3476 17144 3482 17196
rect 4614 17144 4620 17196
rect 4672 17184 4678 17196
rect 4709 17187 4767 17193
rect 4709 17184 4721 17187
rect 4672 17156 4721 17184
rect 4672 17144 4678 17156
rect 4709 17153 4721 17156
rect 4755 17153 4767 17187
rect 4709 17147 4767 17153
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 5353 17187 5411 17193
rect 5353 17184 5365 17187
rect 5316 17156 5365 17184
rect 5316 17144 5322 17156
rect 5353 17153 5365 17156
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 7466 17144 7472 17196
rect 7524 17184 7530 17196
rect 9950 17184 9956 17196
rect 7524 17156 9956 17184
rect 7524 17144 7530 17156
rect 6546 17076 6552 17128
rect 6604 17116 6610 17128
rect 8864 17125 8892 17156
rect 9950 17144 9956 17156
rect 10008 17144 10014 17196
rect 14918 17144 14924 17196
rect 14976 17184 14982 17196
rect 15749 17187 15807 17193
rect 15749 17184 15761 17187
rect 14976 17156 15761 17184
rect 14976 17144 14982 17156
rect 15749 17153 15761 17156
rect 15795 17184 15807 17187
rect 16040 17184 16068 17292
rect 18417 17289 18429 17292
rect 18463 17289 18475 17323
rect 18417 17283 18475 17289
rect 16114 17212 16120 17264
rect 16172 17252 16178 17264
rect 17221 17255 17279 17261
rect 17221 17252 17233 17255
rect 16172 17224 17233 17252
rect 16172 17212 16178 17224
rect 17221 17221 17233 17224
rect 17267 17252 17279 17255
rect 19610 17252 19616 17264
rect 17267 17224 19616 17252
rect 17267 17221 17279 17224
rect 17221 17215 17279 17221
rect 19610 17212 19616 17224
rect 19668 17212 19674 17264
rect 24673 17255 24731 17261
rect 24673 17252 24685 17255
rect 23032 17224 24685 17252
rect 15795 17156 16068 17184
rect 15795 17153 15807 17156
rect 15749 17147 15807 17153
rect 16850 17144 16856 17196
rect 16908 17184 16914 17196
rect 16908 17156 17448 17184
rect 16908 17144 16914 17156
rect 8757 17119 8815 17125
rect 8757 17116 8769 17119
rect 6604 17088 8769 17116
rect 6604 17076 6610 17088
rect 8757 17085 8769 17088
rect 8803 17085 8815 17119
rect 8757 17079 8815 17085
rect 8849 17119 8907 17125
rect 8849 17085 8861 17119
rect 8895 17085 8907 17119
rect 8849 17079 8907 17085
rect 9217 17119 9275 17125
rect 9217 17085 9229 17119
rect 9263 17085 9275 17119
rect 9217 17079 9275 17085
rect 8772 17048 8800 17079
rect 9232 17048 9260 17079
rect 10318 17076 10324 17128
rect 10376 17076 10382 17128
rect 12066 17076 12072 17128
rect 12124 17076 12130 17128
rect 12253 17119 12311 17125
rect 12253 17085 12265 17119
rect 12299 17116 12311 17119
rect 12342 17116 12348 17128
rect 12299 17088 12348 17116
rect 12299 17085 12311 17088
rect 12253 17079 12311 17085
rect 12342 17076 12348 17088
rect 12400 17076 12406 17128
rect 12710 17076 12716 17128
rect 12768 17076 12774 17128
rect 16577 17119 16635 17125
rect 14384 17088 16528 17116
rect 9398 17048 9404 17060
rect 8772 17020 9168 17048
rect 9232 17020 9404 17048
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 6730 16980 6736 16992
rect 4212 16952 6736 16980
rect 4212 16940 4218 16952
rect 6730 16940 6736 16952
rect 6788 16940 6794 16992
rect 8938 16940 8944 16992
rect 8996 16940 9002 16992
rect 9140 16980 9168 17020
rect 9398 17008 9404 17020
rect 9456 17048 9462 17060
rect 14384 17048 14412 17088
rect 9456 17020 14412 17048
rect 9456 17008 9462 17020
rect 15470 17008 15476 17060
rect 15528 17008 15534 17060
rect 16500 17048 16528 17088
rect 16577 17085 16589 17119
rect 16623 17116 16635 17119
rect 16666 17116 16672 17128
rect 16623 17088 16672 17116
rect 16623 17085 16635 17088
rect 16577 17079 16635 17085
rect 16666 17076 16672 17088
rect 16724 17076 16730 17128
rect 17420 17125 17448 17156
rect 16761 17119 16819 17125
rect 16761 17085 16773 17119
rect 16807 17085 16819 17119
rect 16761 17079 16819 17085
rect 17037 17119 17095 17125
rect 17037 17085 17049 17119
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 17405 17119 17463 17125
rect 17405 17085 17417 17119
rect 17451 17085 17463 17119
rect 17405 17079 17463 17085
rect 16776 17048 16804 17079
rect 16500 17020 16804 17048
rect 17052 17048 17080 17079
rect 17586 17076 17592 17128
rect 17644 17116 17650 17128
rect 17865 17119 17923 17125
rect 17865 17116 17877 17119
rect 17644 17088 17877 17116
rect 17644 17076 17650 17088
rect 17865 17085 17877 17088
rect 17911 17085 17923 17119
rect 17865 17079 17923 17085
rect 18230 17076 18236 17128
rect 18288 17076 18294 17128
rect 19426 17076 19432 17128
rect 19484 17116 19490 17128
rect 19705 17119 19763 17125
rect 19705 17116 19717 17119
rect 19484 17088 19717 17116
rect 19484 17076 19490 17088
rect 19705 17085 19717 17088
rect 19751 17085 19763 17119
rect 19705 17079 19763 17085
rect 21634 17076 21640 17128
rect 21692 17076 21698 17128
rect 22002 17076 22008 17128
rect 22060 17116 22066 17128
rect 23032 17125 23060 17224
rect 24673 17221 24685 17224
rect 24719 17221 24731 17255
rect 24673 17215 24731 17221
rect 23290 17144 23296 17196
rect 23348 17184 23354 17196
rect 23348 17156 24072 17184
rect 23348 17144 23354 17156
rect 22281 17119 22339 17125
rect 22281 17116 22293 17119
rect 22060 17088 22293 17116
rect 22060 17076 22066 17088
rect 22281 17085 22293 17088
rect 22327 17085 22339 17119
rect 22281 17079 22339 17085
rect 23017 17119 23075 17125
rect 23017 17085 23029 17119
rect 23063 17085 23075 17119
rect 23017 17079 23075 17085
rect 23106 17076 23112 17128
rect 23164 17076 23170 17128
rect 24044 17125 24072 17156
rect 23477 17119 23535 17125
rect 23477 17085 23489 17119
rect 23523 17085 23535 17119
rect 23477 17079 23535 17085
rect 24029 17119 24087 17125
rect 24029 17085 24041 17119
rect 24075 17085 24087 17119
rect 24029 17079 24087 17085
rect 17052 17020 17724 17048
rect 16776 16992 16804 17020
rect 17696 16992 17724 17020
rect 22646 17008 22652 17060
rect 22704 17048 22710 17060
rect 23492 17048 23520 17079
rect 24302 17076 24308 17128
rect 24360 17076 24366 17128
rect 24578 17076 24584 17128
rect 24636 17116 24642 17128
rect 24857 17119 24915 17125
rect 24857 17116 24869 17119
rect 24636 17088 24869 17116
rect 24636 17076 24642 17088
rect 24857 17085 24869 17088
rect 24903 17085 24915 17119
rect 24857 17079 24915 17085
rect 25222 17076 25228 17128
rect 25280 17116 25286 17128
rect 25501 17119 25559 17125
rect 25501 17116 25513 17119
rect 25280 17088 25513 17116
rect 25280 17076 25286 17088
rect 25501 17085 25513 17088
rect 25547 17085 25559 17119
rect 25501 17079 25559 17085
rect 25866 17076 25872 17128
rect 25924 17116 25930 17128
rect 26145 17119 26203 17125
rect 26145 17116 26157 17119
rect 25924 17088 26157 17116
rect 25924 17076 25930 17088
rect 26145 17085 26157 17088
rect 26191 17085 26203 17119
rect 26145 17079 26203 17085
rect 26786 17076 26792 17128
rect 26844 17076 26850 17128
rect 22704 17020 23520 17048
rect 22704 17008 22710 17020
rect 23658 17008 23664 17060
rect 23716 17048 23722 17060
rect 23716 17020 24164 17048
rect 23716 17008 23722 17020
rect 9858 16980 9864 16992
rect 9140 16952 9864 16980
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 11882 16940 11888 16992
rect 11940 16940 11946 16992
rect 15102 16940 15108 16992
rect 15160 16940 15166 16992
rect 15565 16983 15623 16989
rect 15565 16949 15577 16983
rect 15611 16980 15623 16983
rect 15746 16980 15752 16992
rect 15611 16952 15752 16980
rect 15611 16949 15623 16952
rect 15565 16943 15623 16949
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 16666 16940 16672 16992
rect 16724 16940 16730 16992
rect 16758 16940 16764 16992
rect 16816 16940 16822 16992
rect 17494 16940 17500 16992
rect 17552 16980 17558 16992
rect 17589 16983 17647 16989
rect 17589 16980 17601 16983
rect 17552 16952 17601 16980
rect 17552 16940 17558 16952
rect 17589 16949 17601 16952
rect 17635 16949 17647 16983
rect 17589 16943 17647 16949
rect 17678 16940 17684 16992
rect 17736 16940 17742 16992
rect 19521 16983 19579 16989
rect 19521 16949 19533 16983
rect 19567 16980 19579 16983
rect 20162 16980 20168 16992
rect 19567 16952 20168 16980
rect 19567 16949 19579 16952
rect 19521 16943 19579 16949
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 21450 16940 21456 16992
rect 21508 16940 21514 16992
rect 22094 16940 22100 16992
rect 22152 16940 22158 16992
rect 22738 16940 22744 16992
rect 22796 16980 22802 16992
rect 22833 16983 22891 16989
rect 22833 16980 22845 16983
rect 22796 16952 22845 16980
rect 22796 16940 22802 16952
rect 22833 16949 22845 16952
rect 22879 16949 22891 16983
rect 22833 16943 22891 16949
rect 22922 16940 22928 16992
rect 22980 16980 22986 16992
rect 23293 16983 23351 16989
rect 23293 16980 23305 16983
rect 22980 16952 23305 16980
rect 22980 16940 22986 16952
rect 23293 16949 23305 16952
rect 23339 16949 23351 16983
rect 23293 16943 23351 16949
rect 23566 16940 23572 16992
rect 23624 16980 23630 16992
rect 24136 16989 24164 17020
rect 26602 17008 26608 17060
rect 26660 17008 26666 17060
rect 23845 16983 23903 16989
rect 23845 16980 23857 16983
rect 23624 16952 23857 16980
rect 23624 16940 23630 16952
rect 23845 16949 23857 16952
rect 23891 16949 23903 16983
rect 23845 16943 23903 16949
rect 24121 16983 24179 16989
rect 24121 16949 24133 16983
rect 24167 16949 24179 16983
rect 24121 16943 24179 16949
rect 25314 16940 25320 16992
rect 25372 16940 25378 16992
rect 25958 16940 25964 16992
rect 26016 16940 26022 16992
rect 552 16890 27576 16912
rect 552 16838 7114 16890
rect 7166 16838 7178 16890
rect 7230 16838 7242 16890
rect 7294 16838 7306 16890
rect 7358 16838 7370 16890
rect 7422 16838 13830 16890
rect 13882 16838 13894 16890
rect 13946 16838 13958 16890
rect 14010 16838 14022 16890
rect 14074 16838 14086 16890
rect 14138 16838 20546 16890
rect 20598 16838 20610 16890
rect 20662 16838 20674 16890
rect 20726 16838 20738 16890
rect 20790 16838 20802 16890
rect 20854 16838 27262 16890
rect 27314 16838 27326 16890
rect 27378 16838 27390 16890
rect 27442 16838 27454 16890
rect 27506 16838 27518 16890
rect 27570 16838 27576 16890
rect 552 16816 27576 16838
rect 750 16736 756 16788
rect 808 16776 814 16788
rect 1673 16779 1731 16785
rect 1673 16776 1685 16779
rect 808 16748 1685 16776
rect 808 16736 814 16748
rect 1673 16745 1685 16748
rect 1719 16745 1731 16779
rect 1673 16739 1731 16745
rect 2133 16779 2191 16785
rect 2133 16745 2145 16779
rect 2179 16745 2191 16779
rect 2133 16739 2191 16745
rect 1857 16643 1915 16649
rect 1857 16609 1869 16643
rect 1903 16640 1915 16643
rect 2148 16640 2176 16739
rect 5626 16736 5632 16788
rect 5684 16736 5690 16788
rect 5902 16736 5908 16788
rect 5960 16776 5966 16788
rect 6273 16779 6331 16785
rect 6273 16776 6285 16779
rect 5960 16748 6285 16776
rect 5960 16736 5966 16748
rect 6273 16745 6285 16748
rect 6319 16745 6331 16779
rect 6273 16739 6331 16745
rect 9398 16736 9404 16788
rect 9456 16736 9462 16788
rect 9858 16736 9864 16788
rect 9916 16736 9922 16788
rect 11054 16736 11060 16788
rect 11112 16776 11118 16788
rect 11149 16779 11207 16785
rect 11149 16776 11161 16779
rect 11112 16748 11161 16776
rect 11112 16736 11118 16748
rect 11149 16745 11161 16748
rect 11195 16745 11207 16779
rect 11149 16739 11207 16745
rect 11517 16779 11575 16785
rect 11517 16745 11529 16779
rect 11563 16776 11575 16779
rect 11698 16776 11704 16788
rect 11563 16748 11704 16776
rect 11563 16745 11575 16748
rect 11517 16739 11575 16745
rect 11698 16736 11704 16748
rect 11756 16736 11762 16788
rect 13449 16779 13507 16785
rect 13449 16745 13461 16779
rect 13495 16776 13507 16779
rect 13630 16776 13636 16788
rect 13495 16748 13636 16776
rect 13495 16745 13507 16748
rect 13449 16739 13507 16745
rect 13630 16736 13636 16748
rect 13688 16736 13694 16788
rect 13817 16779 13875 16785
rect 13817 16745 13829 16779
rect 13863 16776 13875 16779
rect 14090 16776 14096 16788
rect 13863 16748 14096 16776
rect 13863 16745 13875 16748
rect 13817 16739 13875 16745
rect 14090 16736 14096 16748
rect 14148 16736 14154 16788
rect 14200 16748 14872 16776
rect 4154 16708 4160 16720
rect 2332 16680 4160 16708
rect 2332 16649 2360 16680
rect 4154 16668 4160 16680
rect 4212 16668 4218 16720
rect 4264 16680 8064 16708
rect 4264 16649 4292 16680
rect 1903 16612 2176 16640
rect 2317 16643 2375 16649
rect 1903 16609 1915 16612
rect 1857 16603 1915 16609
rect 2317 16609 2329 16643
rect 2363 16609 2375 16643
rect 4249 16643 4307 16649
rect 4249 16640 4261 16643
rect 2317 16603 2375 16609
rect 4172 16612 4261 16640
rect 3234 16532 3240 16584
rect 3292 16572 3298 16584
rect 4172 16572 4200 16612
rect 4249 16609 4261 16612
rect 4295 16609 4307 16643
rect 4249 16603 4307 16609
rect 4516 16643 4574 16649
rect 4516 16609 4528 16643
rect 4562 16640 4574 16643
rect 4562 16612 5856 16640
rect 4562 16609 4574 16612
rect 4516 16603 4574 16609
rect 3292 16544 4200 16572
rect 3292 16532 3298 16544
rect 5828 16513 5856 16612
rect 5994 16600 6000 16652
rect 6052 16600 6058 16652
rect 6457 16643 6515 16649
rect 6457 16609 6469 16643
rect 6503 16640 6515 16643
rect 6549 16643 6607 16649
rect 6549 16640 6561 16643
rect 6503 16612 6561 16640
rect 6503 16609 6515 16612
rect 6457 16603 6515 16609
rect 6549 16609 6561 16612
rect 6595 16609 6607 16643
rect 6549 16603 6607 16609
rect 6730 16600 6736 16652
rect 6788 16600 6794 16652
rect 6822 16600 6828 16652
rect 6880 16640 6886 16652
rect 7009 16643 7067 16649
rect 7009 16640 7021 16643
rect 6880 16612 7021 16640
rect 6880 16600 6886 16612
rect 7009 16609 7021 16612
rect 7055 16609 7067 16643
rect 7466 16640 7472 16652
rect 7009 16603 7067 16609
rect 7116 16612 7472 16640
rect 6917 16575 6975 16581
rect 6917 16541 6929 16575
rect 6963 16572 6975 16575
rect 7116 16572 7144 16612
rect 7466 16600 7472 16612
rect 7524 16600 7530 16652
rect 8036 16584 8064 16680
rect 8288 16643 8346 16649
rect 8288 16609 8300 16643
rect 8334 16640 8346 16643
rect 8662 16640 8668 16652
rect 8334 16612 8668 16640
rect 8334 16609 8346 16612
rect 8288 16603 8346 16609
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 9416 16640 9444 16736
rect 9876 16708 9904 16736
rect 10137 16711 10195 16717
rect 10137 16708 10149 16711
rect 9876 16680 10149 16708
rect 10137 16677 10149 16680
rect 10183 16677 10195 16711
rect 10137 16671 10195 16677
rect 10226 16668 10232 16720
rect 10284 16708 10290 16720
rect 10284 16680 11836 16708
rect 10284 16668 10290 16680
rect 9493 16643 9551 16649
rect 9493 16640 9505 16643
rect 9416 16612 9505 16640
rect 9493 16609 9505 16612
rect 9539 16609 9551 16643
rect 9493 16603 9551 16609
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16640 10563 16643
rect 10551 16612 11284 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 6963 16544 7144 16572
rect 6963 16541 6975 16544
rect 6917 16535 6975 16541
rect 8018 16532 8024 16584
rect 8076 16532 8082 16584
rect 11256 16572 11284 16612
rect 11330 16600 11336 16652
rect 11388 16600 11394 16652
rect 11698 16600 11704 16652
rect 11756 16600 11762 16652
rect 11808 16649 11836 16680
rect 11882 16668 11888 16720
rect 11940 16708 11946 16720
rect 12038 16711 12096 16717
rect 12038 16708 12050 16711
rect 11940 16680 12050 16708
rect 11940 16668 11946 16680
rect 12038 16677 12050 16680
rect 12084 16677 12096 16711
rect 14200 16708 14228 16748
rect 14642 16708 14648 16720
rect 12038 16671 12096 16677
rect 12406 16680 14228 16708
rect 14292 16680 14648 16708
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16609 11851 16643
rect 12406 16640 12434 16680
rect 11793 16603 11851 16609
rect 11900 16612 12434 16640
rect 13633 16643 13691 16649
rect 11900 16572 11928 16612
rect 13633 16609 13645 16643
rect 13679 16640 13691 16643
rect 13906 16640 13912 16652
rect 13679 16612 13912 16640
rect 13679 16609 13691 16612
rect 13633 16603 13691 16609
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 14001 16643 14059 16649
rect 14001 16609 14013 16643
rect 14047 16640 14059 16643
rect 14182 16640 14188 16652
rect 14047 16612 14188 16640
rect 14047 16609 14059 16612
rect 14001 16603 14059 16609
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 11256 16544 11928 16572
rect 14292 16513 14320 16680
rect 14642 16668 14648 16680
rect 14700 16668 14706 16720
rect 14844 16708 14872 16748
rect 15102 16736 15108 16788
rect 15160 16776 15166 16788
rect 15197 16779 15255 16785
rect 15197 16776 15209 16779
rect 15160 16748 15209 16776
rect 15160 16736 15166 16748
rect 15197 16745 15209 16748
rect 15243 16745 15255 16779
rect 15197 16739 15255 16745
rect 15562 16736 15568 16788
rect 15620 16776 15626 16788
rect 16301 16779 16359 16785
rect 16301 16776 16313 16779
rect 15620 16748 16313 16776
rect 15620 16736 15626 16748
rect 16301 16745 16313 16748
rect 16347 16745 16359 16779
rect 16942 16776 16948 16788
rect 16301 16739 16359 16745
rect 16408 16748 16948 16776
rect 16408 16708 16436 16748
rect 16942 16736 16948 16748
rect 17000 16776 17006 16788
rect 17310 16776 17316 16788
rect 17000 16748 17316 16776
rect 17000 16736 17006 16748
rect 17310 16736 17316 16748
rect 17368 16736 17374 16788
rect 17494 16736 17500 16788
rect 17552 16736 17558 16788
rect 19705 16779 19763 16785
rect 19705 16776 19717 16779
rect 17788 16748 19717 16776
rect 14844 16680 15608 16708
rect 14461 16643 14519 16649
rect 14461 16609 14473 16643
rect 14507 16640 14519 16643
rect 14507 16612 14780 16640
rect 14507 16609 14519 16612
rect 14461 16603 14519 16609
rect 14752 16513 14780 16612
rect 15102 16600 15108 16652
rect 15160 16600 15166 16652
rect 15580 16649 15608 16680
rect 15948 16680 16436 16708
rect 15565 16643 15623 16649
rect 15565 16609 15577 16643
rect 15611 16609 15623 16643
rect 15565 16603 15623 16609
rect 15654 16600 15660 16652
rect 15712 16640 15718 16652
rect 15948 16649 15976 16680
rect 16758 16668 16764 16720
rect 16816 16668 16822 16720
rect 17221 16711 17279 16717
rect 17221 16677 17233 16711
rect 17267 16708 17279 16711
rect 17405 16711 17463 16717
rect 17405 16708 17417 16711
rect 17267 16680 17417 16708
rect 17267 16677 17279 16680
rect 17221 16671 17279 16677
rect 17405 16677 17417 16680
rect 17451 16708 17463 16711
rect 17678 16708 17684 16720
rect 17451 16680 17684 16708
rect 17451 16677 17463 16680
rect 17405 16671 17463 16677
rect 15749 16643 15807 16649
rect 15749 16640 15761 16643
rect 15712 16612 15761 16640
rect 15712 16600 15718 16612
rect 15749 16609 15761 16612
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16609 15991 16643
rect 15933 16603 15991 16609
rect 16114 16600 16120 16652
rect 16172 16600 16178 16652
rect 16574 16600 16580 16652
rect 16632 16640 16638 16652
rect 17236 16640 17264 16671
rect 17678 16668 17684 16680
rect 17736 16668 17742 16720
rect 16632 16612 17264 16640
rect 16632 16600 16638 16612
rect 15286 16532 15292 16584
rect 15344 16532 15350 16584
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16572 16911 16575
rect 16899 16544 17080 16572
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 5813 16507 5871 16513
rect 5813 16473 5825 16507
rect 5859 16473 5871 16507
rect 5813 16467 5871 16473
rect 14277 16507 14335 16513
rect 14277 16473 14289 16507
rect 14323 16473 14335 16507
rect 14277 16467 14335 16473
rect 14737 16507 14795 16513
rect 14737 16473 14749 16507
rect 14783 16473 14795 16507
rect 17052 16504 17080 16544
rect 17310 16532 17316 16584
rect 17368 16572 17374 16584
rect 17589 16575 17647 16581
rect 17589 16572 17601 16575
rect 17368 16544 17601 16572
rect 17368 16532 17374 16544
rect 17589 16541 17601 16544
rect 17635 16572 17647 16575
rect 17788 16572 17816 16748
rect 19705 16745 19717 16748
rect 19751 16745 19763 16779
rect 19705 16739 19763 16745
rect 23474 16736 23480 16788
rect 23532 16776 23538 16788
rect 24673 16779 24731 16785
rect 24673 16776 24685 16779
rect 23532 16748 24685 16776
rect 23532 16736 23538 16748
rect 24673 16745 24685 16748
rect 24719 16745 24731 16779
rect 24673 16739 24731 16745
rect 19610 16668 19616 16720
rect 19668 16708 19674 16720
rect 19668 16680 21312 16708
rect 19668 16668 19674 16680
rect 18506 16600 18512 16652
rect 18564 16640 18570 16652
rect 19254 16643 19312 16649
rect 19254 16640 19266 16643
rect 18564 16612 19266 16640
rect 18564 16600 18570 16612
rect 19254 16609 19266 16612
rect 19300 16609 19312 16643
rect 19254 16603 19312 16609
rect 20806 16600 20812 16652
rect 20864 16649 20870 16652
rect 20864 16603 20876 16649
rect 20864 16600 20870 16603
rect 17635 16544 17816 16572
rect 17635 16541 17647 16544
rect 17589 16535 17647 16541
rect 19518 16532 19524 16584
rect 19576 16532 19582 16584
rect 21082 16532 21088 16584
rect 21140 16532 21146 16584
rect 21284 16581 21312 16680
rect 22278 16668 22284 16720
rect 22336 16708 22342 16720
rect 23017 16711 23075 16717
rect 23017 16708 23029 16711
rect 22336 16680 23029 16708
rect 22336 16668 22342 16680
rect 23017 16677 23029 16680
rect 23063 16677 23075 16711
rect 25314 16708 25320 16720
rect 23017 16671 23075 16677
rect 23676 16680 25320 16708
rect 21450 16600 21456 16652
rect 21508 16600 21514 16652
rect 21634 16600 21640 16652
rect 21692 16600 21698 16652
rect 21910 16600 21916 16652
rect 21968 16600 21974 16652
rect 22094 16600 22100 16652
rect 22152 16600 22158 16652
rect 22462 16600 22468 16652
rect 22520 16600 22526 16652
rect 22649 16643 22707 16649
rect 22649 16609 22661 16643
rect 22695 16640 22707 16643
rect 22922 16640 22928 16652
rect 22695 16612 22928 16640
rect 22695 16609 22707 16612
rect 22649 16603 22707 16609
rect 22922 16600 22928 16612
rect 22980 16600 22986 16652
rect 23201 16643 23259 16649
rect 23201 16609 23213 16643
rect 23247 16640 23259 16643
rect 23566 16640 23572 16652
rect 23247 16612 23572 16640
rect 23247 16609 23259 16612
rect 23201 16603 23259 16609
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 23676 16649 23704 16680
rect 25314 16668 25320 16680
rect 25372 16668 25378 16720
rect 23661 16643 23719 16649
rect 23661 16609 23673 16643
rect 23707 16609 23719 16643
rect 23661 16603 23719 16609
rect 23750 16600 23756 16652
rect 23808 16640 23814 16652
rect 24029 16643 24087 16649
rect 24029 16640 24041 16643
rect 23808 16612 24041 16640
rect 23808 16600 23814 16612
rect 24029 16609 24041 16612
rect 24075 16609 24087 16643
rect 24029 16603 24087 16609
rect 24397 16643 24455 16649
rect 24397 16609 24409 16643
rect 24443 16640 24455 16643
rect 24670 16640 24676 16652
rect 24443 16612 24676 16640
rect 24443 16609 24455 16612
rect 24397 16603 24455 16609
rect 24670 16600 24676 16612
rect 24728 16600 24734 16652
rect 24949 16643 25007 16649
rect 24949 16609 24961 16643
rect 24995 16640 25007 16643
rect 25038 16640 25044 16652
rect 24995 16612 25044 16640
rect 24995 16609 25007 16612
rect 24949 16603 25007 16609
rect 25038 16600 25044 16612
rect 25096 16600 25102 16652
rect 21269 16575 21327 16581
rect 21269 16541 21281 16575
rect 21315 16572 21327 16575
rect 22281 16575 22339 16581
rect 22281 16572 22293 16575
rect 21315 16544 22293 16572
rect 21315 16541 21327 16544
rect 21269 16535 21327 16541
rect 22281 16541 22293 16544
rect 22327 16572 22339 16575
rect 22833 16575 22891 16581
rect 22833 16572 22845 16575
rect 22327 16544 22845 16572
rect 22327 16541 22339 16544
rect 22281 16535 22339 16541
rect 22833 16541 22845 16544
rect 22879 16572 22891 16575
rect 23014 16572 23020 16584
rect 22879 16544 23020 16572
rect 22879 16541 22891 16544
rect 22833 16535 22891 16541
rect 23014 16532 23020 16544
rect 23072 16572 23078 16584
rect 23385 16575 23443 16581
rect 23385 16572 23397 16575
rect 23072 16544 23397 16572
rect 23072 16532 23078 16544
rect 23385 16541 23397 16544
rect 23431 16572 23443 16575
rect 23477 16575 23535 16581
rect 23477 16572 23489 16575
rect 23431 16544 23489 16572
rect 23431 16541 23443 16544
rect 23385 16535 23443 16541
rect 23477 16541 23489 16544
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 17126 16504 17132 16516
rect 17052 16476 17132 16504
rect 14737 16467 14795 16473
rect 17126 16464 17132 16476
rect 17184 16504 17190 16516
rect 17184 16476 17724 16504
rect 17184 16464 17190 16476
rect 17696 16448 17724 16476
rect 17770 16464 17776 16516
rect 17828 16504 17834 16516
rect 18141 16507 18199 16513
rect 18141 16504 18153 16507
rect 17828 16476 18153 16504
rect 17828 16464 17834 16476
rect 18141 16473 18153 16476
rect 18187 16473 18199 16507
rect 18141 16467 18199 16473
rect 7558 16396 7564 16448
rect 7616 16436 7622 16448
rect 7653 16439 7711 16445
rect 7653 16436 7665 16439
rect 7616 16408 7665 16436
rect 7616 16396 7622 16408
rect 7653 16405 7665 16408
rect 7699 16405 7711 16439
rect 7653 16399 7711 16405
rect 9861 16439 9919 16445
rect 9861 16405 9873 16439
rect 9907 16436 9919 16439
rect 9950 16436 9956 16448
rect 9907 16408 9956 16436
rect 9907 16405 9919 16408
rect 9861 16399 9919 16405
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 10042 16396 10048 16448
rect 10100 16396 10106 16448
rect 11606 16396 11612 16448
rect 11664 16436 11670 16448
rect 13173 16439 13231 16445
rect 13173 16436 13185 16439
rect 11664 16408 13185 16436
rect 11664 16396 11670 16408
rect 13173 16405 13185 16408
rect 13219 16436 13231 16439
rect 13538 16436 13544 16448
rect 13219 16408 13544 16436
rect 13219 16405 13231 16408
rect 13173 16399 13231 16405
rect 13538 16396 13544 16408
rect 13596 16396 13602 16448
rect 16577 16439 16635 16445
rect 16577 16405 16589 16439
rect 16623 16436 16635 16439
rect 16758 16436 16764 16448
rect 16623 16408 16764 16436
rect 16623 16405 16635 16408
rect 16577 16399 16635 16405
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 17678 16396 17684 16448
rect 17736 16396 17742 16448
rect 17954 16396 17960 16448
rect 18012 16396 18018 16448
rect 23845 16439 23903 16445
rect 23845 16405 23857 16439
rect 23891 16436 23903 16439
rect 24578 16436 24584 16448
rect 23891 16408 24584 16436
rect 23891 16405 23903 16408
rect 23845 16399 23903 16405
rect 24578 16396 24584 16408
rect 24636 16396 24642 16448
rect 552 16346 27416 16368
rect 552 16294 3756 16346
rect 3808 16294 3820 16346
rect 3872 16294 3884 16346
rect 3936 16294 3948 16346
rect 4000 16294 4012 16346
rect 4064 16294 10472 16346
rect 10524 16294 10536 16346
rect 10588 16294 10600 16346
rect 10652 16294 10664 16346
rect 10716 16294 10728 16346
rect 10780 16294 17188 16346
rect 17240 16294 17252 16346
rect 17304 16294 17316 16346
rect 17368 16294 17380 16346
rect 17432 16294 17444 16346
rect 17496 16294 23904 16346
rect 23956 16294 23968 16346
rect 24020 16294 24032 16346
rect 24084 16294 24096 16346
rect 24148 16294 24160 16346
rect 24212 16294 27416 16346
rect 552 16272 27416 16294
rect 5534 16192 5540 16244
rect 5592 16232 5598 16244
rect 6457 16235 6515 16241
rect 6457 16232 6469 16235
rect 5592 16204 6469 16232
rect 5592 16192 5598 16204
rect 6457 16201 6469 16204
rect 6503 16232 6515 16235
rect 6822 16232 6828 16244
rect 6503 16204 6828 16232
rect 6503 16201 6515 16204
rect 6457 16195 6515 16201
rect 6822 16192 6828 16204
rect 6880 16192 6886 16244
rect 8110 16232 8116 16244
rect 6932 16204 8116 16232
rect 4617 16167 4675 16173
rect 4617 16133 4629 16167
rect 4663 16164 4675 16167
rect 4798 16164 4804 16176
rect 4663 16136 4804 16164
rect 4663 16133 4675 16136
rect 4617 16127 4675 16133
rect 4798 16124 4804 16136
rect 4856 16164 4862 16176
rect 6638 16164 6644 16176
rect 4856 16136 6644 16164
rect 4856 16124 4862 16136
rect 6638 16124 6644 16136
rect 6696 16164 6702 16176
rect 6932 16164 6960 16204
rect 8110 16192 8116 16204
rect 8168 16192 8174 16244
rect 8662 16192 8668 16244
rect 8720 16192 8726 16244
rect 8938 16192 8944 16244
rect 8996 16232 9002 16244
rect 9033 16235 9091 16241
rect 9033 16232 9045 16235
rect 8996 16204 9045 16232
rect 8996 16192 9002 16204
rect 9033 16201 9045 16204
rect 9079 16201 9091 16235
rect 9033 16195 9091 16201
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 12345 16235 12403 16241
rect 12345 16232 12357 16235
rect 11756 16204 12357 16232
rect 11756 16192 11762 16204
rect 12345 16201 12357 16204
rect 12391 16201 12403 16235
rect 12345 16195 12403 16201
rect 13906 16192 13912 16244
rect 13964 16192 13970 16244
rect 18506 16192 18512 16244
rect 18564 16192 18570 16244
rect 20349 16235 20407 16241
rect 20349 16201 20361 16235
rect 20395 16232 20407 16235
rect 20806 16232 20812 16244
rect 20395 16204 20812 16232
rect 20395 16201 20407 16204
rect 20349 16195 20407 16201
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 23566 16232 23572 16244
rect 22112 16204 23572 16232
rect 6696 16136 6960 16164
rect 16577 16167 16635 16173
rect 6696 16124 6702 16136
rect 16577 16133 16589 16167
rect 16623 16164 16635 16167
rect 16666 16164 16672 16176
rect 16623 16136 16672 16164
rect 16623 16133 16635 16136
rect 16577 16127 16635 16133
rect 16666 16124 16672 16136
rect 16724 16124 16730 16176
rect 17773 16167 17831 16173
rect 17773 16133 17785 16167
rect 17819 16133 17831 16167
rect 17773 16127 17831 16133
rect 19981 16167 20039 16173
rect 19981 16133 19993 16167
rect 20027 16133 20039 16167
rect 19981 16127 20039 16133
rect 3234 16056 3240 16108
rect 3292 16056 3298 16108
rect 7837 16099 7895 16105
rect 5460 16068 6868 16096
rect 2869 16031 2927 16037
rect 2869 15997 2881 16031
rect 2915 16028 2927 16031
rect 3326 16028 3332 16040
rect 2915 16000 3332 16028
rect 2915 15997 2927 16000
rect 2869 15991 2927 15997
rect 3326 15988 3332 16000
rect 3384 15988 3390 16040
rect 5261 16031 5319 16037
rect 5261 15997 5273 16031
rect 5307 15997 5319 16031
rect 5261 15991 5319 15997
rect 3482 15963 3540 15969
rect 3482 15960 3494 15963
rect 3068 15932 3494 15960
rect 3068 15901 3096 15932
rect 3482 15929 3494 15932
rect 3528 15929 3540 15963
rect 5276 15960 5304 15991
rect 5350 15988 5356 16040
rect 5408 15988 5414 16040
rect 5460 16037 5488 16068
rect 5445 16031 5503 16037
rect 5445 15997 5457 16031
rect 5491 15997 5503 16031
rect 5445 15991 5503 15997
rect 5626 15988 5632 16040
rect 5684 15988 5690 16040
rect 6270 15988 6276 16040
rect 6328 15988 6334 16040
rect 6840 16028 6868 16068
rect 7837 16065 7849 16099
rect 7883 16096 7895 16099
rect 8018 16096 8024 16108
rect 7883 16068 8024 16096
rect 7883 16065 7895 16068
rect 7837 16059 7895 16065
rect 8018 16056 8024 16068
rect 8076 16056 8082 16108
rect 8754 16056 8760 16108
rect 8812 16096 8818 16108
rect 8812 16068 9168 16096
rect 8812 16056 8818 16068
rect 8294 16028 8300 16040
rect 6840 16000 8300 16028
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 9140 16037 9168 16068
rect 9674 16056 9680 16108
rect 9732 16096 9738 16108
rect 10226 16096 10232 16108
rect 9732 16068 10232 16096
rect 9732 16056 9738 16068
rect 10226 16056 10232 16068
rect 10284 16056 10290 16108
rect 11974 16056 11980 16108
rect 12032 16096 12038 16108
rect 12989 16099 13047 16105
rect 12032 16068 12112 16096
rect 12032 16056 12038 16068
rect 8849 16031 8907 16037
rect 8849 15997 8861 16031
rect 8895 15997 8907 16031
rect 8849 15991 8907 15997
rect 9125 16031 9183 16037
rect 9125 15997 9137 16031
rect 9171 15997 9183 16031
rect 9125 15991 9183 15997
rect 5721 15963 5779 15969
rect 5721 15960 5733 15963
rect 5276 15932 5733 15960
rect 3482 15923 3540 15929
rect 5721 15929 5733 15932
rect 5767 15929 5779 15963
rect 5721 15923 5779 15929
rect 7466 15920 7472 15972
rect 7524 15960 7530 15972
rect 7570 15963 7628 15969
rect 7570 15960 7582 15963
rect 7524 15932 7582 15960
rect 7524 15920 7530 15932
rect 7570 15929 7582 15932
rect 7616 15929 7628 15963
rect 8864 15960 8892 15991
rect 11606 15988 11612 16040
rect 11664 16028 11670 16040
rect 12084 16037 12112 16068
rect 12989 16065 13001 16099
rect 13035 16096 13047 16099
rect 13078 16096 13084 16108
rect 13035 16068 13084 16096
rect 13035 16065 13047 16068
rect 12989 16059 13047 16065
rect 13078 16056 13084 16068
rect 13136 16096 13142 16108
rect 14461 16099 14519 16105
rect 14461 16096 14473 16099
rect 13136 16068 14473 16096
rect 13136 16056 13142 16068
rect 14461 16065 14473 16068
rect 14507 16096 14519 16099
rect 15286 16096 15292 16108
rect 14507 16068 15292 16096
rect 14507 16065 14519 16068
rect 14461 16059 14519 16065
rect 15286 16056 15292 16068
rect 15344 16096 15350 16108
rect 15344 16068 15424 16096
rect 15344 16056 15350 16068
rect 15396 16037 15424 16068
rect 15746 16056 15752 16108
rect 15804 16096 15810 16108
rect 16761 16099 16819 16105
rect 15804 16068 16712 16096
rect 15804 16056 15810 16068
rect 11701 16031 11759 16037
rect 11701 16028 11713 16031
rect 11664 16000 11713 16028
rect 11664 15988 11670 16000
rect 11701 15997 11713 16000
rect 11747 15997 11759 16031
rect 11701 15991 11759 15997
rect 12069 16031 12127 16037
rect 12069 15997 12081 16031
rect 12115 15997 12127 16031
rect 12069 15991 12127 15997
rect 15381 16031 15439 16037
rect 15381 15997 15393 16031
rect 15427 15997 15439 16031
rect 15381 15991 15439 15997
rect 16301 16031 16359 16037
rect 16301 15997 16313 16031
rect 16347 16028 16359 16031
rect 16485 16031 16543 16037
rect 16485 16028 16497 16031
rect 16347 16000 16497 16028
rect 16347 15997 16359 16000
rect 16301 15991 16359 15997
rect 16485 15997 16497 16000
rect 16531 16028 16543 16031
rect 16574 16028 16580 16040
rect 16531 16000 16580 16028
rect 16531 15997 16543 16000
rect 16485 15991 16543 15997
rect 16574 15988 16580 16000
rect 16632 15988 16638 16040
rect 16684 16028 16712 16068
rect 16761 16065 16773 16099
rect 16807 16096 16819 16099
rect 16942 16096 16948 16108
rect 16807 16068 16948 16096
rect 16807 16065 16819 16068
rect 16761 16059 16819 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 17034 16056 17040 16108
rect 17092 16096 17098 16108
rect 17788 16096 17816 16127
rect 17092 16068 17540 16096
rect 17788 16068 18092 16096
rect 17092 16056 17098 16068
rect 16850 16028 16856 16040
rect 16684 16000 16856 16028
rect 16850 15988 16856 16000
rect 16908 16028 16914 16040
rect 17221 16031 17279 16037
rect 17221 16028 17233 16031
rect 16908 16000 17233 16028
rect 16908 15988 16914 16000
rect 17221 15997 17233 16000
rect 17267 16028 17279 16031
rect 17310 16028 17316 16040
rect 17267 16000 17316 16028
rect 17267 15997 17279 16000
rect 17221 15991 17279 15997
rect 17310 15988 17316 16000
rect 17368 15988 17374 16040
rect 17512 16037 17540 16068
rect 17497 16031 17555 16037
rect 17497 15997 17509 16031
rect 17543 15997 17555 16031
rect 17497 15991 17555 15997
rect 9306 15960 9312 15972
rect 8864 15932 9312 15960
rect 7570 15923 7628 15929
rect 9306 15920 9312 15932
rect 9364 15920 9370 15972
rect 10318 15920 10324 15972
rect 10376 15960 10382 15972
rect 10474 15963 10532 15969
rect 10474 15960 10486 15963
rect 10376 15932 10486 15960
rect 10376 15920 10382 15932
rect 10474 15929 10486 15932
rect 10520 15929 10532 15963
rect 10474 15923 10532 15929
rect 11514 15920 11520 15972
rect 11572 15960 11578 15972
rect 11885 15963 11943 15969
rect 11885 15960 11897 15963
rect 11572 15932 11897 15960
rect 11572 15920 11578 15932
rect 11885 15929 11897 15932
rect 11931 15929 11943 15963
rect 11885 15923 11943 15929
rect 11974 15920 11980 15972
rect 12032 15920 12038 15972
rect 12158 15920 12164 15972
rect 12216 15960 12222 15972
rect 12713 15963 12771 15969
rect 12713 15960 12725 15963
rect 12216 15932 12725 15960
rect 12216 15920 12222 15932
rect 12713 15929 12725 15932
rect 12759 15929 12771 15963
rect 12713 15923 12771 15929
rect 15010 15920 15016 15972
rect 15068 15920 15074 15972
rect 17405 15963 17463 15969
rect 17405 15929 17417 15963
rect 17451 15929 17463 15963
rect 17512 15960 17540 15991
rect 17586 15988 17592 16040
rect 17644 15988 17650 16040
rect 17770 15988 17776 16040
rect 17828 16028 17834 16040
rect 18064 16037 18092 16068
rect 18138 16056 18144 16108
rect 18196 16096 18202 16108
rect 19996 16096 20024 16127
rect 18196 16068 19748 16096
rect 19996 16068 20392 16096
rect 18196 16056 18202 16068
rect 17865 16031 17923 16037
rect 17865 16028 17877 16031
rect 17828 16000 17877 16028
rect 17828 15988 17834 16000
rect 17865 15997 17877 16000
rect 17911 15997 17923 16031
rect 17865 15991 17923 15997
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 18233 16031 18291 16037
rect 18233 15997 18245 16031
rect 18279 16028 18291 16031
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 18279 16000 18337 16028
rect 18279 15997 18291 16000
rect 18233 15991 18291 15997
rect 18325 15997 18337 16000
rect 18371 15997 18383 16031
rect 18325 15991 18383 15997
rect 19610 15988 19616 16040
rect 19668 15988 19674 16040
rect 18874 15960 18880 15972
rect 17512 15932 18880 15960
rect 17405 15923 17463 15929
rect 3053 15895 3111 15901
rect 3053 15861 3065 15895
rect 3099 15861 3111 15895
rect 3053 15855 3111 15861
rect 4985 15895 5043 15901
rect 4985 15861 4997 15895
rect 5031 15892 5043 15895
rect 5902 15892 5908 15904
rect 5031 15864 5908 15892
rect 5031 15861 5043 15864
rect 4985 15855 5043 15861
rect 5902 15852 5908 15864
rect 5960 15852 5966 15904
rect 11609 15895 11667 15901
rect 11609 15861 11621 15895
rect 11655 15892 11667 15895
rect 11992 15892 12020 15920
rect 11655 15864 12020 15892
rect 11655 15861 11667 15864
rect 11609 15855 11667 15861
rect 12250 15852 12256 15904
rect 12308 15852 12314 15904
rect 12805 15895 12863 15901
rect 12805 15861 12817 15895
rect 12851 15892 12863 15895
rect 13170 15892 13176 15904
rect 12851 15864 13176 15892
rect 12851 15861 12863 15864
rect 12805 15855 12863 15861
rect 13170 15852 13176 15864
rect 13228 15852 13234 15904
rect 13722 15852 13728 15904
rect 13780 15892 13786 15904
rect 14277 15895 14335 15901
rect 14277 15892 14289 15895
rect 13780 15864 14289 15892
rect 13780 15852 13786 15864
rect 14277 15861 14289 15864
rect 14323 15861 14335 15895
rect 14277 15855 14335 15861
rect 14369 15895 14427 15901
rect 14369 15861 14381 15895
rect 14415 15892 14427 15895
rect 14458 15892 14464 15904
rect 14415 15864 14464 15892
rect 14415 15861 14427 15864
rect 14369 15855 14427 15861
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 16206 15852 16212 15904
rect 16264 15852 16270 15904
rect 16942 15852 16948 15904
rect 17000 15892 17006 15904
rect 17420 15892 17448 15923
rect 18874 15920 18880 15932
rect 18932 15920 18938 15972
rect 19334 15920 19340 15972
rect 19392 15960 19398 15972
rect 19521 15963 19579 15969
rect 19521 15960 19533 15963
rect 19392 15932 19533 15960
rect 19392 15920 19398 15932
rect 19521 15929 19533 15932
rect 19567 15929 19579 15963
rect 19720 15960 19748 16068
rect 20364 16037 20392 16068
rect 19889 16031 19947 16037
rect 19889 15997 19901 16031
rect 19935 16028 19947 16031
rect 20257 16031 20315 16037
rect 20257 16028 20269 16031
rect 19935 16000 20269 16028
rect 19935 15997 19947 16000
rect 19889 15991 19947 15997
rect 20257 15997 20269 16000
rect 20303 15997 20315 16031
rect 20257 15991 20315 15997
rect 20349 16031 20407 16037
rect 20349 15997 20361 16031
rect 20395 15997 20407 16031
rect 20349 15991 20407 15997
rect 19981 15963 20039 15969
rect 19981 15960 19993 15963
rect 19720 15932 19993 15960
rect 19521 15923 19579 15929
rect 19981 15929 19993 15932
rect 20027 15929 20039 15963
rect 20272 15960 20300 15991
rect 20438 15988 20444 16040
rect 20496 16028 20502 16040
rect 22112 16038 22140 16204
rect 23566 16192 23572 16204
rect 23624 16192 23630 16244
rect 25958 16164 25964 16176
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 20496 16000 20545 16028
rect 20496 15988 20502 16000
rect 20533 15997 20545 16000
rect 20579 16028 20591 16031
rect 22066 16028 22140 16038
rect 20579 16010 22140 16028
rect 22756 16136 25964 16164
rect 20579 16000 22094 16010
rect 20579 15997 20591 16000
rect 20533 15991 20591 15997
rect 22756 15960 22784 16136
rect 25958 16124 25964 16136
rect 26016 16124 26022 16176
rect 23658 16096 23664 16108
rect 22940 16068 23664 16096
rect 22940 16037 22968 16068
rect 23658 16056 23664 16068
rect 23716 16056 23722 16108
rect 22925 16031 22983 16037
rect 22925 15997 22937 16031
rect 22971 15997 22983 16031
rect 22925 15991 22983 15997
rect 23014 15988 23020 16040
rect 23072 15988 23078 16040
rect 23106 15988 23112 16040
rect 23164 16028 23170 16040
rect 24029 16031 24087 16037
rect 24029 16028 24041 16031
rect 23164 16000 24041 16028
rect 23164 15988 23170 16000
rect 24029 15997 24041 16000
rect 24075 16028 24087 16031
rect 26602 16028 26608 16040
rect 24075 16000 26608 16028
rect 24075 15997 24087 16000
rect 24029 15991 24087 15997
rect 26602 15988 26608 16000
rect 26660 15988 26666 16040
rect 20272 15932 22784 15960
rect 19981 15923 20039 15929
rect 17000 15864 17448 15892
rect 17000 15852 17006 15864
rect 17862 15852 17868 15904
rect 17920 15892 17926 15904
rect 20165 15895 20223 15901
rect 20165 15892 20177 15895
rect 17920 15864 20177 15892
rect 17920 15852 17926 15864
rect 20165 15861 20177 15864
rect 20211 15892 20223 15895
rect 21266 15892 21272 15904
rect 20211 15864 21272 15892
rect 20211 15861 20223 15864
rect 20165 15855 20223 15861
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 22738 15852 22744 15904
rect 22796 15852 22802 15904
rect 23658 15852 23664 15904
rect 23716 15892 23722 15904
rect 23937 15895 23995 15901
rect 23937 15892 23949 15895
rect 23716 15864 23949 15892
rect 23716 15852 23722 15864
rect 23937 15861 23949 15864
rect 23983 15861 23995 15895
rect 23937 15855 23995 15861
rect 552 15802 27576 15824
rect 552 15750 7114 15802
rect 7166 15750 7178 15802
rect 7230 15750 7242 15802
rect 7294 15750 7306 15802
rect 7358 15750 7370 15802
rect 7422 15750 13830 15802
rect 13882 15750 13894 15802
rect 13946 15750 13958 15802
rect 14010 15750 14022 15802
rect 14074 15750 14086 15802
rect 14138 15750 20546 15802
rect 20598 15750 20610 15802
rect 20662 15750 20674 15802
rect 20726 15750 20738 15802
rect 20790 15750 20802 15802
rect 20854 15750 27262 15802
rect 27314 15750 27326 15802
rect 27378 15750 27390 15802
rect 27442 15750 27454 15802
rect 27506 15750 27518 15802
rect 27570 15750 27576 15802
rect 552 15728 27576 15750
rect 3326 15648 3332 15700
rect 3384 15648 3390 15700
rect 6270 15688 6276 15700
rect 4540 15660 6276 15688
rect 4540 15629 4568 15660
rect 6270 15648 6276 15660
rect 6328 15688 6334 15700
rect 7193 15691 7251 15697
rect 7193 15688 7205 15691
rect 6328 15660 7205 15688
rect 6328 15648 6334 15660
rect 7193 15657 7205 15660
rect 7239 15657 7251 15691
rect 7193 15651 7251 15657
rect 7285 15691 7343 15697
rect 7285 15657 7297 15691
rect 7331 15688 7343 15691
rect 7466 15688 7472 15700
rect 7331 15660 7472 15688
rect 7331 15657 7343 15660
rect 7285 15651 7343 15657
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 10042 15648 10048 15700
rect 10100 15688 10106 15700
rect 11333 15691 11391 15697
rect 11333 15688 11345 15691
rect 10100 15660 11345 15688
rect 10100 15648 10106 15660
rect 11333 15657 11345 15660
rect 11379 15657 11391 15691
rect 11333 15651 11391 15657
rect 13170 15648 13176 15700
rect 13228 15648 13234 15700
rect 13538 15648 13544 15700
rect 13596 15648 13602 15700
rect 14458 15648 14464 15700
rect 14516 15648 14522 15700
rect 14921 15691 14979 15697
rect 14921 15657 14933 15691
rect 14967 15688 14979 15691
rect 15930 15688 15936 15700
rect 14967 15660 15936 15688
rect 14967 15657 14979 15660
rect 14921 15651 14979 15657
rect 15930 15648 15936 15660
rect 15988 15648 15994 15700
rect 19613 15691 19671 15697
rect 19613 15657 19625 15691
rect 19659 15657 19671 15691
rect 23106 15688 23112 15700
rect 19613 15651 19671 15657
rect 20088 15660 23112 15688
rect 4525 15623 4583 15629
rect 4525 15589 4537 15623
rect 4571 15589 4583 15623
rect 4525 15583 4583 15589
rect 4617 15623 4675 15629
rect 4617 15589 4629 15623
rect 4663 15620 4675 15623
rect 4982 15620 4988 15632
rect 4663 15592 4988 15620
rect 4663 15589 4675 15592
rect 4617 15583 4675 15589
rect 4982 15580 4988 15592
rect 5040 15580 5046 15632
rect 5169 15623 5227 15629
rect 5169 15589 5181 15623
rect 5215 15620 5227 15623
rect 5534 15620 5540 15632
rect 5215 15592 5540 15620
rect 5215 15589 5227 15592
rect 5169 15583 5227 15589
rect 5534 15580 5540 15592
rect 5592 15580 5598 15632
rect 8018 15620 8024 15632
rect 5828 15592 8024 15620
rect 3513 15555 3571 15561
rect 3513 15521 3525 15555
rect 3559 15552 3571 15555
rect 3559 15524 4292 15552
rect 3559 15521 3571 15524
rect 3513 15515 3571 15521
rect 3602 15444 3608 15496
rect 3660 15484 3666 15496
rect 3697 15487 3755 15493
rect 3697 15484 3709 15487
rect 3660 15456 3709 15484
rect 3660 15444 3666 15456
rect 3697 15453 3709 15456
rect 3743 15453 3755 15487
rect 3697 15447 3755 15453
rect 4264 15425 4292 15524
rect 4430 15512 4436 15564
rect 4488 15512 4494 15564
rect 4798 15512 4804 15564
rect 4856 15512 4862 15564
rect 5077 15555 5135 15561
rect 5077 15521 5089 15555
rect 5123 15521 5135 15555
rect 5077 15515 5135 15521
rect 5261 15555 5319 15561
rect 5261 15521 5273 15555
rect 5307 15521 5319 15555
rect 5261 15515 5319 15521
rect 4448 15484 4476 15512
rect 5092 15484 5120 15515
rect 4448 15456 5120 15484
rect 4249 15419 4307 15425
rect 4249 15385 4261 15419
rect 4295 15385 4307 15419
rect 4249 15379 4307 15385
rect 4982 15376 4988 15428
rect 5040 15416 5046 15428
rect 5276 15416 5304 15515
rect 5442 15512 5448 15564
rect 5500 15512 5506 15564
rect 5828 15561 5856 15592
rect 8018 15580 8024 15592
rect 8076 15580 8082 15632
rect 8110 15580 8116 15632
rect 8168 15620 8174 15632
rect 14829 15623 14887 15629
rect 14829 15620 14841 15623
rect 8168 15592 14841 15620
rect 8168 15580 8174 15592
rect 14829 15589 14841 15592
rect 14875 15589 14887 15623
rect 14829 15583 14887 15589
rect 15286 15580 15292 15632
rect 15344 15580 15350 15632
rect 16393 15623 16451 15629
rect 16393 15589 16405 15623
rect 16439 15620 16451 15623
rect 17862 15620 17868 15632
rect 16439 15592 17868 15620
rect 16439 15589 16451 15592
rect 16393 15583 16451 15589
rect 17862 15580 17868 15592
rect 17920 15580 17926 15632
rect 17957 15623 18015 15629
rect 17957 15589 17969 15623
rect 18003 15620 18015 15623
rect 19628 15620 19656 15651
rect 19950 15623 20008 15629
rect 19950 15620 19962 15623
rect 18003 15592 19564 15620
rect 19628 15592 19962 15620
rect 18003 15589 18015 15592
rect 17957 15583 18015 15589
rect 5813 15555 5871 15561
rect 5813 15521 5825 15555
rect 5859 15521 5871 15555
rect 5813 15515 5871 15521
rect 5902 15512 5908 15564
rect 5960 15552 5966 15564
rect 6069 15555 6127 15561
rect 6069 15552 6081 15555
rect 5960 15524 6081 15552
rect 5960 15512 5966 15524
rect 6069 15521 6081 15524
rect 6115 15521 6127 15555
rect 6069 15515 6127 15521
rect 7558 15512 7564 15564
rect 7616 15512 7622 15564
rect 7653 15555 7711 15561
rect 7653 15521 7665 15555
rect 7699 15521 7711 15555
rect 7653 15515 7711 15521
rect 7745 15555 7803 15561
rect 7745 15521 7757 15555
rect 7791 15521 7803 15555
rect 7745 15515 7803 15521
rect 5040 15388 5304 15416
rect 5040 15376 5046 15388
rect 4798 15308 4804 15360
rect 4856 15348 4862 15360
rect 4893 15351 4951 15357
rect 4893 15348 4905 15351
rect 4856 15320 4905 15348
rect 4856 15308 4862 15320
rect 4893 15317 4905 15320
rect 4939 15317 4951 15351
rect 4893 15311 4951 15317
rect 5350 15308 5356 15360
rect 5408 15348 5414 15360
rect 7668 15348 7696 15515
rect 7760 15484 7788 15515
rect 7926 15512 7932 15564
rect 7984 15512 7990 15564
rect 11790 15512 11796 15564
rect 11848 15512 11854 15564
rect 11974 15512 11980 15564
rect 12032 15552 12038 15564
rect 12621 15555 12679 15561
rect 12621 15552 12633 15555
rect 12032 15524 12633 15552
rect 12032 15512 12038 15524
rect 12621 15521 12633 15524
rect 12667 15521 12679 15555
rect 12621 15515 12679 15521
rect 12802 15512 12808 15564
rect 12860 15552 12866 15564
rect 12860 15524 15148 15552
rect 12860 15512 12866 15524
rect 9401 15487 9459 15493
rect 9401 15484 9413 15487
rect 7760 15456 9413 15484
rect 9401 15453 9413 15456
rect 9447 15453 9459 15487
rect 9401 15447 9459 15453
rect 9582 15444 9588 15496
rect 9640 15444 9646 15496
rect 9677 15487 9735 15493
rect 9677 15453 9689 15487
rect 9723 15484 9735 15487
rect 11238 15484 11244 15496
rect 9723 15456 11244 15484
rect 9723 15453 9735 15456
rect 9677 15447 9735 15453
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 11701 15487 11759 15493
rect 11701 15453 11713 15487
rect 11747 15484 11759 15487
rect 12158 15484 12164 15496
rect 11747 15456 12164 15484
rect 11747 15453 11759 15456
rect 11701 15447 11759 15453
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13817 15487 13875 15493
rect 13817 15453 13829 15487
rect 13863 15484 13875 15487
rect 14090 15484 14096 15496
rect 13863 15456 14096 15484
rect 13863 15453 13875 15456
rect 13817 15447 13875 15453
rect 10962 15376 10968 15428
rect 11020 15416 11026 15428
rect 12069 15419 12127 15425
rect 12069 15416 12081 15419
rect 11020 15388 12081 15416
rect 11020 15376 11026 15388
rect 12069 15385 12081 15388
rect 12115 15385 12127 15419
rect 13648 15416 13676 15447
rect 14090 15444 14096 15456
rect 14148 15484 14154 15496
rect 14918 15484 14924 15496
rect 14148 15456 14924 15484
rect 14148 15444 14154 15456
rect 14918 15444 14924 15456
rect 14976 15484 14982 15496
rect 15013 15487 15071 15493
rect 15013 15484 15025 15487
rect 14976 15456 15025 15484
rect 14976 15444 14982 15456
rect 15013 15453 15025 15456
rect 15059 15453 15071 15487
rect 15120 15484 15148 15524
rect 15654 15512 15660 15564
rect 15712 15552 15718 15564
rect 16117 15555 16175 15561
rect 16117 15552 16129 15555
rect 15712 15524 16129 15552
rect 15712 15512 15718 15524
rect 16117 15521 16129 15524
rect 16163 15552 16175 15555
rect 16206 15552 16212 15564
rect 16163 15524 16212 15552
rect 16163 15521 16175 15524
rect 16117 15515 16175 15521
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 16758 15512 16764 15564
rect 16816 15512 16822 15564
rect 17770 15512 17776 15564
rect 17828 15512 17834 15564
rect 18598 15512 18604 15564
rect 18656 15512 18662 15564
rect 18785 15555 18843 15561
rect 18785 15521 18797 15555
rect 18831 15552 18843 15555
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 18831 15524 19441 15552
rect 18831 15521 18843 15524
rect 18785 15515 18843 15521
rect 19429 15521 19441 15524
rect 19475 15521 19487 15555
rect 19536 15552 19564 15592
rect 19950 15589 19962 15592
rect 19996 15589 20008 15623
rect 19950 15583 20008 15589
rect 20088 15552 20116 15660
rect 23106 15648 23112 15660
rect 23164 15648 23170 15700
rect 23198 15648 23204 15700
rect 23256 15648 23262 15700
rect 25222 15620 25228 15632
rect 21836 15592 25228 15620
rect 19536 15524 20116 15552
rect 19429 15515 19487 15521
rect 21082 15512 21088 15564
rect 21140 15552 21146 15564
rect 21836 15561 21864 15592
rect 22094 15561 22100 15564
rect 21821 15555 21879 15561
rect 21821 15552 21833 15555
rect 21140 15524 21833 15552
rect 21140 15512 21146 15524
rect 21821 15521 21833 15524
rect 21867 15521 21879 15555
rect 21821 15515 21879 15521
rect 22088 15515 22100 15561
rect 22094 15512 22100 15515
rect 22152 15512 22158 15564
rect 23198 15512 23204 15564
rect 23256 15552 23262 15564
rect 24044 15561 24072 15592
rect 25222 15580 25228 15592
rect 25280 15580 25286 15632
rect 23845 15555 23903 15561
rect 23845 15552 23857 15555
rect 23256 15524 23857 15552
rect 23256 15512 23262 15524
rect 23845 15521 23857 15524
rect 23891 15521 23903 15555
rect 23845 15515 23903 15521
rect 24029 15555 24087 15561
rect 24029 15521 24041 15555
rect 24075 15521 24087 15555
rect 24029 15515 24087 15521
rect 24296 15555 24354 15561
rect 24296 15521 24308 15555
rect 24342 15552 24354 15555
rect 24762 15552 24768 15564
rect 24342 15524 24768 15552
rect 24342 15521 24354 15524
rect 24296 15515 24354 15521
rect 24762 15512 24768 15524
rect 24820 15512 24826 15564
rect 17788 15484 17816 15512
rect 15120 15456 17816 15484
rect 15013 15447 15071 15453
rect 18230 15444 18236 15496
rect 18288 15484 18294 15496
rect 18417 15487 18475 15493
rect 18417 15484 18429 15487
rect 18288 15456 18429 15484
rect 18288 15444 18294 15456
rect 18417 15453 18429 15456
rect 18463 15453 18475 15487
rect 18417 15447 18475 15453
rect 19518 15444 19524 15496
rect 19576 15484 19582 15496
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 19576 15456 19717 15484
rect 19576 15444 19582 15456
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 17034 15416 17040 15428
rect 13648 15388 17040 15416
rect 12069 15379 12127 15385
rect 17034 15376 17040 15388
rect 17092 15416 17098 15428
rect 19058 15416 19064 15428
rect 17092 15388 19064 15416
rect 17092 15376 17098 15388
rect 19058 15376 19064 15388
rect 19116 15376 19122 15428
rect 22830 15376 22836 15428
rect 22888 15416 22894 15428
rect 23293 15419 23351 15425
rect 23293 15416 23305 15419
rect 22888 15388 23305 15416
rect 22888 15376 22894 15388
rect 23293 15385 23305 15388
rect 23339 15385 23351 15419
rect 23293 15379 23351 15385
rect 8754 15348 8760 15360
rect 5408 15320 8760 15348
rect 5408 15308 5414 15320
rect 8754 15308 8760 15320
rect 8812 15308 8818 15360
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 11977 15351 12035 15357
rect 11977 15348 11989 15351
rect 11204 15320 11989 15348
rect 11204 15308 11210 15320
rect 11977 15317 11989 15320
rect 12023 15317 12035 15351
rect 11977 15311 12035 15317
rect 16390 15308 16396 15360
rect 16448 15348 16454 15360
rect 16945 15351 17003 15357
rect 16945 15348 16957 15351
rect 16448 15320 16957 15348
rect 16448 15308 16454 15320
rect 16945 15317 16957 15320
rect 16991 15317 17003 15351
rect 16945 15311 17003 15317
rect 19886 15308 19892 15360
rect 19944 15348 19950 15360
rect 20438 15348 20444 15360
rect 19944 15320 20444 15348
rect 19944 15308 19950 15320
rect 20438 15308 20444 15320
rect 20496 15308 20502 15360
rect 21082 15308 21088 15360
rect 21140 15308 21146 15360
rect 25038 15308 25044 15360
rect 25096 15348 25102 15360
rect 25409 15351 25467 15357
rect 25409 15348 25421 15351
rect 25096 15320 25421 15348
rect 25096 15308 25102 15320
rect 25409 15317 25421 15320
rect 25455 15317 25467 15351
rect 25409 15311 25467 15317
rect 552 15258 27416 15280
rect 552 15206 3756 15258
rect 3808 15206 3820 15258
rect 3872 15206 3884 15258
rect 3936 15206 3948 15258
rect 4000 15206 4012 15258
rect 4064 15206 10472 15258
rect 10524 15206 10536 15258
rect 10588 15206 10600 15258
rect 10652 15206 10664 15258
rect 10716 15206 10728 15258
rect 10780 15206 17188 15258
rect 17240 15206 17252 15258
rect 17304 15206 17316 15258
rect 17368 15206 17380 15258
rect 17432 15206 17444 15258
rect 17496 15206 23904 15258
rect 23956 15206 23968 15258
rect 24020 15206 24032 15258
rect 24084 15206 24096 15258
rect 24148 15206 24160 15258
rect 24212 15206 27416 15258
rect 552 15184 27416 15206
rect 4985 15147 5043 15153
rect 4985 15113 4997 15147
rect 5031 15144 5043 15147
rect 5994 15144 6000 15156
rect 5031 15116 6000 15144
rect 5031 15113 5043 15116
rect 4985 15107 5043 15113
rect 5994 15104 6000 15116
rect 6052 15104 6058 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 9401 15147 9459 15153
rect 9401 15144 9413 15147
rect 8352 15116 9413 15144
rect 8352 15104 8358 15116
rect 9401 15113 9413 15116
rect 9447 15113 9459 15147
rect 9401 15107 9459 15113
rect 10318 15104 10324 15156
rect 10376 15144 10382 15156
rect 10689 15147 10747 15153
rect 10689 15144 10701 15147
rect 10376 15116 10701 15144
rect 10376 15104 10382 15116
rect 10689 15113 10701 15116
rect 10735 15113 10747 15147
rect 10689 15107 10747 15113
rect 12621 15147 12679 15153
rect 12621 15113 12633 15147
rect 12667 15144 12679 15147
rect 12710 15144 12716 15156
rect 12667 15116 12716 15144
rect 12667 15113 12679 15116
rect 12621 15107 12679 15113
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 12986 15104 12992 15156
rect 13044 15144 13050 15156
rect 14921 15147 14979 15153
rect 14921 15144 14933 15147
rect 13044 15116 14933 15144
rect 13044 15104 13050 15116
rect 14921 15113 14933 15116
rect 14967 15113 14979 15147
rect 14921 15107 14979 15113
rect 17681 15147 17739 15153
rect 17681 15113 17693 15147
rect 17727 15144 17739 15147
rect 18598 15144 18604 15156
rect 17727 15116 18604 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 18598 15104 18604 15116
rect 18656 15104 18662 15156
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 23750 15144 23756 15156
rect 18748 15116 23756 15144
rect 18748 15104 18754 15116
rect 23750 15104 23756 15116
rect 23808 15104 23814 15156
rect 24762 15104 24768 15156
rect 24820 15104 24826 15156
rect 6454 15076 6460 15088
rect 5920 15048 6460 15076
rect 5813 15011 5871 15017
rect 5813 15008 5825 15011
rect 5368 14980 5825 15008
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4617 14943 4675 14949
rect 4617 14940 4629 14943
rect 4120 14912 4629 14940
rect 4120 14900 4126 14912
rect 4617 14909 4629 14912
rect 4663 14909 4675 14943
rect 4617 14903 4675 14909
rect 4798 14900 4804 14952
rect 4856 14900 4862 14952
rect 5368 14949 5396 14980
rect 5813 14977 5825 14980
rect 5859 14977 5871 15011
rect 5813 14971 5871 14977
rect 5353 14943 5411 14949
rect 5353 14909 5365 14943
rect 5399 14909 5411 14943
rect 5353 14903 5411 14909
rect 5442 14900 5448 14952
rect 5500 14900 5506 14952
rect 5537 14943 5595 14949
rect 5537 14909 5549 14943
rect 5583 14909 5595 14943
rect 5537 14903 5595 14909
rect 5074 14832 5080 14884
rect 5132 14832 5138 14884
rect 5552 14804 5580 14903
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 5721 14943 5779 14949
rect 5721 14940 5733 14943
rect 5684 14912 5733 14940
rect 5684 14900 5690 14912
rect 5721 14909 5733 14912
rect 5767 14940 5779 14943
rect 5920 14940 5948 15048
rect 6454 15036 6460 15048
rect 6512 15076 6518 15088
rect 7926 15076 7932 15088
rect 6512 15048 7932 15076
rect 6512 15036 6518 15048
rect 7926 15036 7932 15048
rect 7984 15076 7990 15088
rect 9030 15076 9036 15088
rect 7984 15048 9036 15076
rect 7984 15036 7990 15048
rect 9030 15036 9036 15048
rect 9088 15076 9094 15088
rect 11698 15076 11704 15088
rect 9088 15048 11704 15076
rect 9088 15036 9094 15048
rect 11698 15036 11704 15048
rect 11756 15036 11762 15088
rect 13722 15076 13728 15088
rect 12360 15048 13728 15076
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 15008 9735 15011
rect 12360 15008 12388 15048
rect 13722 15036 13728 15048
rect 13780 15076 13786 15088
rect 15562 15076 15568 15088
rect 13780 15048 15568 15076
rect 13780 15036 13786 15048
rect 15562 15036 15568 15048
rect 15620 15076 15626 15088
rect 16298 15076 16304 15088
rect 15620 15048 16304 15076
rect 15620 15036 15626 15048
rect 16298 15036 16304 15048
rect 16356 15036 16362 15088
rect 16390 15036 16396 15088
rect 16448 15076 16454 15088
rect 16448 15048 17448 15076
rect 16448 15036 16454 15048
rect 9723 14980 12388 15008
rect 9723 14977 9735 14980
rect 9677 14971 9735 14977
rect 13170 14968 13176 15020
rect 13228 14968 13234 15020
rect 13814 14968 13820 15020
rect 13872 15008 13878 15020
rect 14090 15008 14096 15020
rect 13872 14980 14096 15008
rect 13872 14968 13878 14980
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 14458 15008 14464 15020
rect 14384 14980 14464 15008
rect 5767 14912 5948 14940
rect 5767 14909 5779 14912
rect 5721 14903 5779 14909
rect 6362 14900 6368 14952
rect 6420 14900 6426 14952
rect 8938 14900 8944 14952
rect 8996 14940 9002 14952
rect 9217 14943 9275 14949
rect 9217 14940 9229 14943
rect 8996 14912 9229 14940
rect 8996 14900 9002 14912
rect 9217 14909 9229 14912
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 9582 14900 9588 14952
rect 9640 14900 9646 14952
rect 10042 14900 10048 14952
rect 10100 14940 10106 14952
rect 10137 14943 10195 14949
rect 10137 14940 10149 14943
rect 10100 14912 10149 14940
rect 10100 14900 10106 14912
rect 10137 14909 10149 14912
rect 10183 14909 10195 14943
rect 10137 14903 10195 14909
rect 10962 14900 10968 14952
rect 11020 14900 11026 14952
rect 11057 14943 11115 14949
rect 11057 14909 11069 14943
rect 11103 14909 11115 14943
rect 11057 14903 11115 14909
rect 8570 14804 8576 14816
rect 5552 14776 8576 14804
rect 8570 14764 8576 14776
rect 8628 14764 8634 14816
rect 8662 14764 8668 14816
rect 8720 14764 8726 14816
rect 8754 14764 8760 14816
rect 8812 14804 8818 14816
rect 10321 14807 10379 14813
rect 10321 14804 10333 14807
rect 8812 14776 10333 14804
rect 8812 14764 8818 14776
rect 10321 14773 10333 14776
rect 10367 14804 10379 14807
rect 11072 14804 11100 14903
rect 11146 14900 11152 14952
rect 11204 14900 11210 14952
rect 11333 14943 11391 14949
rect 11333 14909 11345 14943
rect 11379 14940 11391 14943
rect 11698 14940 11704 14952
rect 11379 14912 11704 14940
rect 11379 14909 11391 14912
rect 11333 14903 11391 14909
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 12066 14900 12072 14952
rect 12124 14900 12130 14952
rect 12250 14900 12256 14952
rect 12308 14900 12314 14952
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 12802 14940 12808 14952
rect 12492 14912 12808 14940
rect 12492 14900 12498 14912
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 12989 14943 13047 14949
rect 12989 14909 13001 14943
rect 13035 14940 13047 14943
rect 14384 14940 14412 14980
rect 14458 14968 14464 14980
rect 14516 15008 14522 15020
rect 17218 15008 17224 15020
rect 14516 14980 17224 15008
rect 14516 14968 14522 14980
rect 17218 14968 17224 14980
rect 17276 14968 17282 15020
rect 17420 15008 17448 15048
rect 18138 15036 18144 15088
rect 18196 15036 18202 15088
rect 19702 15036 19708 15088
rect 19760 15076 19766 15088
rect 20073 15079 20131 15085
rect 20073 15076 20085 15079
rect 19760 15048 20085 15076
rect 19760 15036 19766 15048
rect 20073 15045 20085 15048
rect 20119 15045 20131 15079
rect 20073 15039 20131 15045
rect 24305 15079 24363 15085
rect 24305 15045 24317 15079
rect 24351 15076 24363 15079
rect 25406 15076 25412 15088
rect 24351 15048 25412 15076
rect 24351 15045 24363 15048
rect 24305 15039 24363 15045
rect 25406 15036 25412 15048
rect 25464 15036 25470 15088
rect 17586 15008 17592 15020
rect 17420 14980 17592 15008
rect 13035 14912 14412 14940
rect 15105 14943 15163 14949
rect 13035 14909 13047 14912
rect 12989 14903 13047 14909
rect 15105 14909 15117 14943
rect 15151 14940 15163 14943
rect 15654 14940 15660 14952
rect 15151 14912 15660 14940
rect 15151 14909 15163 14912
rect 15105 14903 15163 14909
rect 11422 14832 11428 14884
rect 11480 14872 11486 14884
rect 13004 14872 13032 14903
rect 15654 14900 15660 14912
rect 15712 14900 15718 14952
rect 15930 14900 15936 14952
rect 15988 14940 15994 14952
rect 16025 14943 16083 14949
rect 16025 14940 16037 14943
rect 15988 14912 16037 14940
rect 15988 14900 15994 14912
rect 16025 14909 16037 14912
rect 16071 14909 16083 14943
rect 16025 14903 16083 14909
rect 16298 14900 16304 14952
rect 16356 14900 16362 14952
rect 16390 14900 16396 14952
rect 16448 14900 16454 14952
rect 17034 14900 17040 14952
rect 17092 14940 17098 14952
rect 17512 14949 17540 14980
rect 17586 14968 17592 14980
rect 17644 14968 17650 15020
rect 24486 15008 24492 15020
rect 24320 14980 24492 15008
rect 17129 14943 17187 14949
rect 17129 14940 17141 14943
rect 17092 14912 17141 14940
rect 17092 14900 17098 14912
rect 17129 14909 17141 14912
rect 17175 14909 17187 14943
rect 17129 14903 17187 14909
rect 17497 14943 17555 14949
rect 17497 14909 17509 14943
rect 17543 14909 17555 14943
rect 17497 14903 17555 14909
rect 18322 14900 18328 14952
rect 18380 14900 18386 14952
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14940 18751 14943
rect 19518 14940 19524 14952
rect 18739 14912 19524 14940
rect 18739 14909 18751 14912
rect 18693 14903 18751 14909
rect 19518 14900 19524 14912
rect 19576 14900 19582 14952
rect 24026 14900 24032 14952
rect 24084 14900 24090 14952
rect 24320 14949 24348 14980
rect 24486 14968 24492 14980
rect 24544 15008 24550 15020
rect 25041 15011 25099 15017
rect 25041 15008 25053 15011
rect 24544 14980 25053 15008
rect 24544 14968 24550 14980
rect 25041 14977 25053 14980
rect 25087 14977 25099 15011
rect 25041 14971 25099 14977
rect 24305 14943 24363 14949
rect 24305 14909 24317 14943
rect 24351 14909 24363 14943
rect 24854 14940 24860 14952
rect 24305 14903 24363 14909
rect 24504 14912 24860 14940
rect 11480 14844 13032 14872
rect 11480 14832 11486 14844
rect 13906 14832 13912 14884
rect 13964 14832 13970 14884
rect 16209 14875 16267 14881
rect 16209 14841 16221 14875
rect 16255 14872 16267 14875
rect 16942 14872 16948 14884
rect 16255 14844 16948 14872
rect 16255 14841 16267 14844
rect 16209 14835 16267 14841
rect 16942 14832 16948 14844
rect 17000 14872 17006 14884
rect 17313 14875 17371 14881
rect 17313 14872 17325 14875
rect 17000 14844 17325 14872
rect 17000 14832 17006 14844
rect 17313 14841 17325 14844
rect 17359 14841 17371 14875
rect 17313 14835 17371 14841
rect 10367 14776 11100 14804
rect 13081 14807 13139 14813
rect 10367 14773 10379 14776
rect 10321 14767 10379 14773
rect 13081 14773 13093 14807
rect 13127 14804 13139 14807
rect 13541 14807 13599 14813
rect 13541 14804 13553 14807
rect 13127 14776 13553 14804
rect 13127 14773 13139 14776
rect 13081 14767 13139 14773
rect 13541 14773 13553 14776
rect 13587 14773 13599 14807
rect 13541 14767 13599 14773
rect 14001 14807 14059 14813
rect 14001 14773 14013 14807
rect 14047 14804 14059 14807
rect 16022 14804 16028 14816
rect 14047 14776 16028 14804
rect 14047 14773 14059 14776
rect 14001 14767 14059 14773
rect 16022 14764 16028 14776
rect 16080 14764 16086 14816
rect 16577 14807 16635 14813
rect 16577 14773 16589 14807
rect 16623 14804 16635 14807
rect 17126 14804 17132 14816
rect 16623 14776 17132 14804
rect 16623 14773 16635 14776
rect 16577 14767 16635 14773
rect 17126 14764 17132 14776
rect 17184 14764 17190 14816
rect 17328 14804 17356 14835
rect 17402 14832 17408 14884
rect 17460 14832 17466 14884
rect 17865 14875 17923 14881
rect 17865 14841 17877 14875
rect 17911 14841 17923 14875
rect 18949 14875 19007 14881
rect 18949 14872 18961 14875
rect 17865 14835 17923 14841
rect 18892 14844 18961 14872
rect 17770 14804 17776 14816
rect 17328 14776 17776 14804
rect 17770 14764 17776 14776
rect 17828 14804 17834 14816
rect 17880 14804 17908 14835
rect 17828 14776 17908 14804
rect 18509 14807 18567 14813
rect 17828 14764 17834 14776
rect 18509 14773 18521 14807
rect 18555 14804 18567 14807
rect 18892 14804 18920 14844
rect 18949 14841 18961 14844
rect 18995 14841 19007 14875
rect 18949 14835 19007 14841
rect 24121 14875 24179 14881
rect 24121 14841 24133 14875
rect 24167 14872 24179 14875
rect 24504 14872 24532 14912
rect 24854 14900 24860 14912
rect 24912 14900 24918 14952
rect 24946 14900 24952 14952
rect 25004 14900 25010 14952
rect 25593 14943 25651 14949
rect 25593 14909 25605 14943
rect 25639 14909 25651 14943
rect 25593 14903 25651 14909
rect 24167 14844 24532 14872
rect 24581 14875 24639 14881
rect 24167 14841 24179 14844
rect 24121 14835 24179 14841
rect 24581 14841 24593 14875
rect 24627 14841 24639 14875
rect 24581 14835 24639 14841
rect 18555 14776 18920 14804
rect 18555 14773 18567 14776
rect 18509 14767 18567 14773
rect 19058 14764 19064 14816
rect 19116 14804 19122 14816
rect 21082 14804 21088 14816
rect 19116 14776 21088 14804
rect 19116 14764 19122 14776
rect 21082 14764 21088 14776
rect 21140 14804 21146 14816
rect 21450 14804 21456 14816
rect 21140 14776 21456 14804
rect 21140 14764 21146 14776
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 23934 14764 23940 14816
rect 23992 14804 23998 14816
rect 24394 14804 24400 14816
rect 23992 14776 24400 14804
rect 23992 14764 23998 14776
rect 24394 14764 24400 14776
rect 24452 14804 24458 14816
rect 24489 14807 24547 14813
rect 24489 14804 24501 14807
rect 24452 14776 24501 14804
rect 24452 14764 24458 14776
rect 24489 14773 24501 14776
rect 24535 14773 24547 14807
rect 24596 14804 24624 14835
rect 24670 14832 24676 14884
rect 24728 14872 24734 14884
rect 25608 14872 25636 14903
rect 24728 14844 25636 14872
rect 24728 14832 24734 14844
rect 25038 14804 25044 14816
rect 24596 14776 25044 14804
rect 24489 14767 24547 14773
rect 25038 14764 25044 14776
rect 25096 14764 25102 14816
rect 552 14714 27576 14736
rect 552 14662 7114 14714
rect 7166 14662 7178 14714
rect 7230 14662 7242 14714
rect 7294 14662 7306 14714
rect 7358 14662 7370 14714
rect 7422 14662 13830 14714
rect 13882 14662 13894 14714
rect 13946 14662 13958 14714
rect 14010 14662 14022 14714
rect 14074 14662 14086 14714
rect 14138 14662 20546 14714
rect 20598 14662 20610 14714
rect 20662 14662 20674 14714
rect 20726 14662 20738 14714
rect 20790 14662 20802 14714
rect 20854 14662 27262 14714
rect 27314 14662 27326 14714
rect 27378 14662 27390 14714
rect 27442 14662 27454 14714
rect 27506 14662 27518 14714
rect 27570 14662 27576 14714
rect 552 14640 27576 14662
rect 3697 14603 3755 14609
rect 3697 14569 3709 14603
rect 3743 14600 3755 14603
rect 4522 14600 4528 14612
rect 3743 14572 4528 14600
rect 3743 14569 3755 14572
rect 3697 14563 3755 14569
rect 4522 14560 4528 14572
rect 4580 14560 4586 14612
rect 6362 14600 6368 14612
rect 4632 14572 6368 14600
rect 4632 14541 4660 14572
rect 6362 14560 6368 14572
rect 6420 14600 6426 14612
rect 7193 14603 7251 14609
rect 7193 14600 7205 14603
rect 6420 14572 7205 14600
rect 6420 14560 6426 14572
rect 7193 14569 7205 14572
rect 7239 14569 7251 14603
rect 7193 14563 7251 14569
rect 8938 14560 8944 14612
rect 8996 14600 9002 14612
rect 9398 14600 9404 14612
rect 8996 14572 9404 14600
rect 8996 14560 9002 14572
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 9769 14603 9827 14609
rect 9769 14569 9781 14603
rect 9815 14600 9827 14603
rect 9950 14600 9956 14612
rect 9815 14572 9956 14600
rect 9815 14569 9827 14572
rect 9769 14563 9827 14569
rect 9950 14560 9956 14572
rect 10008 14600 10014 14612
rect 10318 14600 10324 14612
rect 10008 14572 10324 14600
rect 10008 14560 10014 14572
rect 10318 14560 10324 14572
rect 10376 14600 10382 14612
rect 10689 14603 10747 14609
rect 10689 14600 10701 14603
rect 10376 14572 10701 14600
rect 10376 14560 10382 14572
rect 10689 14569 10701 14572
rect 10735 14569 10747 14603
rect 10689 14563 10747 14569
rect 12342 14560 12348 14612
rect 12400 14560 12406 14612
rect 12805 14603 12863 14609
rect 12805 14569 12817 14603
rect 12851 14600 12863 14603
rect 13173 14603 13231 14609
rect 13173 14600 13185 14603
rect 12851 14572 13185 14600
rect 12851 14569 12863 14572
rect 12805 14563 12863 14569
rect 13173 14569 13185 14572
rect 13219 14569 13231 14603
rect 13173 14563 13231 14569
rect 14182 14560 14188 14612
rect 14240 14600 14246 14612
rect 14553 14603 14611 14609
rect 14553 14600 14565 14603
rect 14240 14572 14565 14600
rect 14240 14560 14246 14572
rect 14553 14569 14565 14572
rect 14599 14569 14611 14603
rect 14553 14563 14611 14569
rect 17313 14603 17371 14609
rect 17313 14569 17325 14603
rect 17359 14600 17371 14603
rect 18322 14600 18328 14612
rect 17359 14572 18328 14600
rect 17359 14569 17371 14572
rect 17313 14563 17371 14569
rect 18322 14560 18328 14572
rect 18380 14560 18386 14612
rect 19337 14603 19395 14609
rect 19337 14569 19349 14603
rect 19383 14600 19395 14603
rect 21821 14603 21879 14609
rect 19383 14572 19748 14600
rect 19383 14569 19395 14572
rect 19337 14563 19395 14569
rect 4617 14535 4675 14541
rect 4617 14501 4629 14535
rect 4663 14501 4675 14535
rect 4617 14495 4675 14501
rect 4709 14535 4767 14541
rect 4709 14501 4721 14535
rect 4755 14532 4767 14535
rect 4982 14532 4988 14544
rect 4755 14504 4988 14532
rect 4755 14501 4767 14504
rect 4709 14495 4767 14501
rect 4982 14492 4988 14504
rect 5040 14492 5046 14544
rect 6914 14532 6920 14544
rect 5828 14504 6920 14532
rect 2590 14473 2596 14476
rect 2584 14427 2596 14473
rect 2590 14424 2596 14427
rect 2648 14424 2654 14476
rect 3973 14467 4031 14473
rect 3973 14433 3985 14467
rect 4019 14464 4031 14467
rect 4019 14436 4384 14464
rect 4019 14433 4031 14436
rect 3973 14427 4031 14433
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14365 2375 14399
rect 2317 14359 2375 14365
rect 2332 14260 2360 14359
rect 4062 14356 4068 14408
rect 4120 14396 4126 14408
rect 4157 14399 4215 14405
rect 4157 14396 4169 14399
rect 4120 14368 4169 14396
rect 4120 14356 4126 14368
rect 4157 14365 4169 14368
rect 4203 14365 4215 14399
rect 4157 14359 4215 14365
rect 3326 14288 3332 14340
rect 3384 14328 3390 14340
rect 3789 14331 3847 14337
rect 3789 14328 3801 14331
rect 3384 14300 3801 14328
rect 3384 14288 3390 14300
rect 3789 14297 3801 14300
rect 3835 14297 3847 14331
rect 3789 14291 3847 14297
rect 2498 14260 2504 14272
rect 2332 14232 2504 14260
rect 2498 14220 2504 14232
rect 2556 14220 2562 14272
rect 3602 14220 3608 14272
rect 3660 14260 3666 14272
rect 4172 14260 4200 14359
rect 4356 14337 4384 14436
rect 4430 14424 4436 14476
rect 4488 14464 4494 14476
rect 4525 14467 4583 14473
rect 4525 14464 4537 14467
rect 4488 14436 4537 14464
rect 4488 14424 4494 14436
rect 4525 14433 4537 14436
rect 4571 14433 4583 14467
rect 4525 14427 4583 14433
rect 4890 14424 4896 14476
rect 4948 14424 4954 14476
rect 5258 14424 5264 14476
rect 5316 14464 5322 14476
rect 5828 14473 5856 14504
rect 6914 14492 6920 14504
rect 6972 14532 6978 14544
rect 8018 14532 8024 14544
rect 6972 14504 8024 14532
rect 6972 14492 6978 14504
rect 7576 14473 7604 14504
rect 8018 14492 8024 14504
rect 8076 14492 8082 14544
rect 8570 14492 8576 14544
rect 8628 14532 8634 14544
rect 10045 14535 10103 14541
rect 10045 14532 10057 14535
rect 8628 14504 10057 14532
rect 8628 14492 8634 14504
rect 10045 14501 10057 14504
rect 10091 14501 10103 14535
rect 10045 14495 10103 14501
rect 10134 14492 10140 14544
rect 10192 14532 10198 14544
rect 13541 14535 13599 14541
rect 13541 14532 13553 14535
rect 10192 14504 13553 14532
rect 10192 14492 10198 14504
rect 13541 14501 13553 14504
rect 13587 14501 13599 14535
rect 13541 14495 13599 14501
rect 17678 14492 17684 14544
rect 17736 14532 17742 14544
rect 19426 14532 19432 14544
rect 17736 14504 19432 14532
rect 17736 14492 17742 14504
rect 19426 14492 19432 14504
rect 19484 14492 19490 14544
rect 19720 14532 19748 14572
rect 21821 14569 21833 14603
rect 21867 14600 21879 14603
rect 22094 14600 22100 14612
rect 21867 14572 22100 14600
rect 21867 14569 21879 14572
rect 21821 14563 21879 14569
rect 22094 14560 22100 14572
rect 22152 14560 22158 14612
rect 23109 14603 23167 14609
rect 23109 14600 23121 14603
rect 22204 14572 23121 14600
rect 19777 14535 19835 14541
rect 19777 14532 19789 14535
rect 19720 14504 19789 14532
rect 19777 14501 19789 14504
rect 19823 14501 19835 14535
rect 22204 14532 22232 14572
rect 23109 14569 23121 14572
rect 23155 14569 23167 14603
rect 23109 14563 23167 14569
rect 24581 14603 24639 14609
rect 24581 14569 24593 14603
rect 24627 14600 24639 14603
rect 24946 14600 24952 14612
rect 24627 14572 24952 14600
rect 24627 14569 24639 14572
rect 24581 14563 24639 14569
rect 24946 14560 24952 14572
rect 25004 14560 25010 14612
rect 22557 14535 22615 14541
rect 22557 14532 22569 14535
rect 19777 14495 19835 14501
rect 22112 14504 22232 14532
rect 22296 14504 22569 14532
rect 5813 14467 5871 14473
rect 5813 14464 5825 14467
rect 5316 14436 5825 14464
rect 5316 14424 5322 14436
rect 5813 14433 5825 14436
rect 5859 14433 5871 14467
rect 6069 14467 6127 14473
rect 6069 14464 6081 14467
rect 5813 14427 5871 14433
rect 5920 14436 6081 14464
rect 5074 14356 5080 14408
rect 5132 14396 5138 14408
rect 5920 14396 5948 14436
rect 6069 14433 6081 14436
rect 6115 14433 6127 14467
rect 6069 14427 6127 14433
rect 7561 14467 7619 14473
rect 7561 14433 7573 14467
rect 7607 14433 7619 14467
rect 7561 14427 7619 14433
rect 7828 14467 7886 14473
rect 7828 14433 7840 14467
rect 7874 14464 7886 14467
rect 8386 14464 8392 14476
rect 7874 14436 8392 14464
rect 7874 14433 7886 14436
rect 7828 14427 7886 14433
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 9401 14467 9459 14473
rect 9401 14433 9413 14467
rect 9447 14464 9459 14467
rect 12713 14467 12771 14473
rect 12713 14464 12725 14467
rect 9447 14436 12725 14464
rect 9447 14433 9459 14436
rect 9401 14427 9459 14433
rect 12713 14433 12725 14436
rect 12759 14464 12771 14467
rect 14921 14467 14979 14473
rect 14921 14464 14933 14467
rect 12759 14436 13492 14464
rect 12759 14433 12771 14436
rect 12713 14427 12771 14433
rect 5132 14368 5948 14396
rect 9309 14399 9367 14405
rect 5132 14356 5138 14368
rect 9309 14365 9321 14399
rect 9355 14396 9367 14399
rect 9582 14396 9588 14408
rect 9355 14368 9588 14396
rect 9355 14365 9367 14368
rect 9309 14359 9367 14365
rect 9582 14356 9588 14368
rect 9640 14396 9646 14408
rect 10226 14396 10232 14408
rect 9640 14368 10232 14396
rect 9640 14356 9646 14368
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 11422 14396 11428 14408
rect 10367 14368 11428 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 11422 14356 11428 14368
rect 11480 14356 11486 14408
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 12897 14399 12955 14405
rect 12897 14396 12909 14399
rect 11848 14368 12909 14396
rect 11848 14356 11854 14368
rect 12897 14365 12909 14368
rect 12943 14396 12955 14399
rect 13170 14396 13176 14408
rect 12943 14368 13176 14396
rect 12943 14365 12955 14368
rect 12897 14359 12955 14365
rect 13170 14356 13176 14368
rect 13228 14356 13234 14408
rect 4341 14331 4399 14337
rect 4341 14297 4353 14331
rect 4387 14297 4399 14331
rect 4341 14291 4399 14297
rect 8496 14300 9240 14328
rect 7834 14260 7840 14272
rect 3660 14232 7840 14260
rect 3660 14220 3666 14232
rect 7834 14220 7840 14232
rect 7892 14260 7898 14272
rect 8496 14260 8524 14300
rect 7892 14232 8524 14260
rect 7892 14220 7898 14232
rect 8846 14220 8852 14272
rect 8904 14260 8910 14272
rect 9125 14263 9183 14269
rect 9125 14260 9137 14263
rect 8904 14232 9137 14260
rect 8904 14220 8910 14232
rect 9125 14229 9137 14232
rect 9171 14229 9183 14263
rect 9212 14260 9240 14300
rect 12434 14260 12440 14272
rect 9212 14232 12440 14260
rect 9125 14223 9183 14229
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 13464 14260 13492 14436
rect 13556 14436 14933 14464
rect 13556 14408 13584 14436
rect 14921 14433 14933 14436
rect 14967 14433 14979 14467
rect 14921 14427 14979 14433
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 16114 14464 16120 14476
rect 15252 14436 16120 14464
rect 15252 14424 15258 14436
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 17126 14424 17132 14476
rect 17184 14424 17190 14476
rect 17218 14424 17224 14476
rect 17276 14464 17282 14476
rect 17862 14464 17868 14476
rect 17276 14436 17868 14464
rect 17276 14424 17282 14436
rect 17862 14424 17868 14436
rect 17920 14424 17926 14476
rect 18230 14424 18236 14476
rect 18288 14424 18294 14476
rect 18322 14424 18328 14476
rect 18380 14424 18386 14476
rect 18509 14467 18567 14473
rect 18509 14433 18521 14467
rect 18555 14464 18567 14467
rect 19153 14467 19211 14473
rect 19153 14464 19165 14467
rect 18555 14436 19165 14464
rect 18555 14433 18567 14436
rect 18509 14427 18567 14433
rect 19153 14433 19165 14436
rect 19199 14433 19211 14467
rect 21174 14464 21180 14476
rect 19153 14427 19211 14433
rect 19444 14436 21180 14464
rect 13538 14356 13544 14408
rect 13596 14356 13602 14408
rect 13633 14399 13691 14405
rect 13633 14365 13645 14399
rect 13679 14365 13691 14399
rect 13633 14359 13691 14365
rect 13648 14328 13676 14359
rect 13722 14356 13728 14408
rect 13780 14356 13786 14408
rect 14734 14356 14740 14408
rect 14792 14396 14798 14408
rect 15013 14399 15071 14405
rect 15013 14396 15025 14399
rect 14792 14368 15025 14396
rect 14792 14356 14798 14368
rect 15013 14365 15025 14368
rect 15059 14365 15071 14399
rect 15013 14359 15071 14365
rect 15102 14356 15108 14408
rect 15160 14356 15166 14408
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14396 17003 14399
rect 18248 14396 18276 14424
rect 16991 14368 18276 14396
rect 16991 14365 17003 14368
rect 16945 14359 17003 14365
rect 16850 14328 16856 14340
rect 13648 14300 16856 14328
rect 16850 14288 16856 14300
rect 16908 14328 16914 14340
rect 19444 14328 19472 14436
rect 21174 14424 21180 14436
rect 21232 14424 21238 14476
rect 22112 14473 22140 14504
rect 22097 14467 22155 14473
rect 22097 14433 22109 14467
rect 22143 14433 22155 14467
rect 22097 14427 22155 14433
rect 22186 14424 22192 14476
rect 22244 14424 22250 14476
rect 22296 14473 22324 14504
rect 22557 14501 22569 14504
rect 22603 14501 22615 14535
rect 22557 14495 22615 14501
rect 22925 14535 22983 14541
rect 22925 14501 22937 14535
rect 22971 14532 22983 14535
rect 23934 14532 23940 14544
rect 22971 14504 23940 14532
rect 22971 14501 22983 14504
rect 22925 14495 22983 14501
rect 22281 14467 22339 14473
rect 22281 14433 22293 14467
rect 22327 14433 22339 14467
rect 22281 14427 22339 14433
rect 22370 14424 22376 14476
rect 22428 14464 22434 14476
rect 22465 14467 22523 14473
rect 22465 14464 22477 14467
rect 22428 14436 22477 14464
rect 22428 14424 22434 14436
rect 22465 14433 22477 14436
rect 22511 14433 22523 14467
rect 22465 14427 22523 14433
rect 22741 14467 22799 14473
rect 22741 14433 22753 14467
rect 22787 14464 22799 14467
rect 22830 14464 22836 14476
rect 22787 14436 22836 14464
rect 22787 14433 22799 14436
rect 22741 14427 22799 14433
rect 22830 14424 22836 14436
rect 22888 14424 22894 14476
rect 23124 14473 23152 14504
rect 23934 14492 23940 14504
rect 23992 14492 23998 14544
rect 25222 14492 25228 14544
rect 25280 14532 25286 14544
rect 25280 14504 26280 14532
rect 25280 14492 25286 14504
rect 23017 14467 23075 14473
rect 23017 14433 23029 14467
rect 23063 14433 23075 14467
rect 23017 14427 23075 14433
rect 23109 14467 23167 14473
rect 23109 14433 23121 14467
rect 23155 14433 23167 14467
rect 23109 14427 23167 14433
rect 19518 14356 19524 14408
rect 19576 14356 19582 14408
rect 16908 14300 19472 14328
rect 16908 14288 16914 14300
rect 14642 14260 14648 14272
rect 13464 14232 14648 14260
rect 14642 14220 14648 14232
rect 14700 14260 14706 14272
rect 15838 14260 15844 14272
rect 14700 14232 15844 14260
rect 14700 14220 14706 14232
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 15930 14220 15936 14272
rect 15988 14260 15994 14272
rect 19426 14260 19432 14272
rect 15988 14232 19432 14260
rect 15988 14220 15994 14232
rect 19426 14220 19432 14232
rect 19484 14220 19490 14272
rect 19536 14260 19564 14356
rect 23032 14328 23060 14427
rect 23290 14424 23296 14476
rect 23348 14424 23354 14476
rect 24397 14467 24455 14473
rect 24397 14433 24409 14467
rect 24443 14462 24455 14467
rect 24486 14462 24492 14476
rect 24443 14434 24492 14462
rect 24443 14433 24455 14434
rect 24397 14427 24455 14433
rect 24486 14424 24492 14434
rect 24544 14424 24550 14476
rect 25498 14424 25504 14476
rect 25556 14464 25562 14476
rect 26252 14473 26280 14504
rect 25970 14467 26028 14473
rect 25970 14464 25982 14467
rect 25556 14436 25982 14464
rect 25556 14424 25562 14436
rect 25970 14433 25982 14436
rect 26016 14433 26028 14467
rect 25970 14427 26028 14433
rect 26237 14467 26295 14473
rect 26237 14433 26249 14467
rect 26283 14433 26295 14467
rect 26237 14427 26295 14433
rect 24026 14356 24032 14408
rect 24084 14396 24090 14408
rect 24305 14399 24363 14405
rect 24305 14396 24317 14399
rect 24084 14368 24317 14396
rect 24084 14356 24090 14368
rect 24305 14365 24317 14368
rect 24351 14365 24363 14399
rect 24305 14359 24363 14365
rect 23290 14328 23296 14340
rect 23032 14300 23296 14328
rect 23290 14288 23296 14300
rect 23348 14288 23354 14340
rect 19794 14260 19800 14272
rect 19536 14232 19800 14260
rect 19794 14220 19800 14232
rect 19852 14220 19858 14272
rect 20898 14220 20904 14272
rect 20956 14220 20962 14272
rect 23658 14220 23664 14272
rect 23716 14260 23722 14272
rect 24029 14263 24087 14269
rect 24029 14260 24041 14263
rect 23716 14232 24041 14260
rect 23716 14220 23722 14232
rect 24029 14229 24041 14232
rect 24075 14229 24087 14263
rect 24320 14260 24348 14359
rect 24670 14288 24676 14340
rect 24728 14328 24734 14340
rect 24857 14331 24915 14337
rect 24857 14328 24869 14331
rect 24728 14300 24869 14328
rect 24728 14288 24734 14300
rect 24857 14297 24869 14300
rect 24903 14297 24915 14331
rect 24857 14291 24915 14297
rect 25590 14260 25596 14272
rect 24320 14232 25596 14260
rect 24029 14223 24087 14229
rect 25590 14220 25596 14232
rect 25648 14220 25654 14272
rect 552 14170 27416 14192
rect 552 14118 3756 14170
rect 3808 14118 3820 14170
rect 3872 14118 3884 14170
rect 3936 14118 3948 14170
rect 4000 14118 4012 14170
rect 4064 14118 10472 14170
rect 10524 14118 10536 14170
rect 10588 14118 10600 14170
rect 10652 14118 10664 14170
rect 10716 14118 10728 14170
rect 10780 14118 17188 14170
rect 17240 14118 17252 14170
rect 17304 14118 17316 14170
rect 17368 14118 17380 14170
rect 17432 14118 17444 14170
rect 17496 14118 23904 14170
rect 23956 14118 23968 14170
rect 24020 14118 24032 14170
rect 24084 14118 24096 14170
rect 24148 14118 24160 14170
rect 24212 14118 27416 14170
rect 552 14096 27416 14118
rect 2590 14016 2596 14068
rect 2648 14056 2654 14068
rect 2777 14059 2835 14065
rect 2777 14056 2789 14059
rect 2648 14028 2789 14056
rect 2648 14016 2654 14028
rect 2777 14025 2789 14028
rect 2823 14025 2835 14059
rect 2777 14019 2835 14025
rect 4982 14016 4988 14068
rect 5040 14056 5046 14068
rect 9490 14056 9496 14068
rect 5040 14028 9496 14056
rect 5040 14016 5046 14028
rect 9490 14016 9496 14028
rect 9548 14056 9554 14068
rect 9548 14028 10088 14056
rect 9548 14016 9554 14028
rect 3881 13991 3939 13997
rect 3881 13957 3893 13991
rect 3927 13988 3939 13991
rect 4246 13988 4252 14000
rect 3927 13960 4252 13988
rect 3927 13957 3939 13960
rect 3881 13951 3939 13957
rect 4246 13948 4252 13960
rect 4304 13948 4310 14000
rect 8386 13948 8392 14000
rect 8444 13948 8450 14000
rect 9122 13948 9128 14000
rect 9180 13948 9186 14000
rect 9950 13988 9956 14000
rect 9324 13960 9956 13988
rect 2498 13880 2504 13932
rect 2556 13920 2562 13932
rect 2556 13892 4292 13920
rect 2556 13880 2562 13892
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13852 3019 13855
rect 3326 13852 3332 13864
rect 3007 13824 3332 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 4264 13852 4292 13892
rect 5258 13880 5264 13932
rect 5316 13880 5322 13932
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 5500 13892 5764 13920
rect 5500 13880 5506 13892
rect 5276 13852 5304 13880
rect 5736 13864 5764 13892
rect 4264 13824 5304 13852
rect 5626 13812 5632 13864
rect 5684 13812 5690 13864
rect 5718 13812 5724 13864
rect 5776 13812 5782 13864
rect 5810 13812 5816 13864
rect 5868 13812 5874 13864
rect 5997 13855 6055 13861
rect 5997 13821 6009 13855
rect 6043 13852 6055 13855
rect 6454 13852 6460 13864
rect 6043 13824 6460 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 7834 13812 7840 13864
rect 7892 13812 7898 13864
rect 8018 13812 8024 13864
rect 8076 13812 8082 13864
rect 8662 13812 8668 13864
rect 8720 13812 8726 13864
rect 8754 13812 8760 13864
rect 8812 13812 8818 13864
rect 8846 13812 8852 13864
rect 8904 13812 8910 13864
rect 9030 13812 9036 13864
rect 9088 13812 9094 13864
rect 9324 13861 9352 13960
rect 9950 13948 9956 13960
rect 10008 13948 10014 14000
rect 10060 13988 10088 14028
rect 11330 14016 11336 14068
rect 11388 14056 11394 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11388 14028 11989 14056
rect 11388 14016 11394 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 11977 14019 12035 14025
rect 12618 14016 12624 14068
rect 12676 14016 12682 14068
rect 14734 14016 14740 14068
rect 14792 14016 14798 14068
rect 14918 14016 14924 14068
rect 14976 14056 14982 14068
rect 14976 14028 15332 14056
rect 14976 14016 14982 14028
rect 11514 13988 11520 14000
rect 10060 13960 11520 13988
rect 11514 13948 11520 13960
rect 11572 13988 11578 14000
rect 12636 13988 12664 14016
rect 11572 13960 12664 13988
rect 14645 13991 14703 13997
rect 11572 13948 11578 13960
rect 14645 13957 14657 13991
rect 14691 13988 14703 13991
rect 15194 13988 15200 14000
rect 14691 13960 15200 13988
rect 14691 13957 14703 13960
rect 14645 13951 14703 13957
rect 15194 13948 15200 13960
rect 15252 13948 15258 14000
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 9769 13923 9827 13929
rect 9769 13920 9781 13923
rect 9640 13892 9781 13920
rect 9640 13880 9646 13892
rect 9769 13889 9781 13892
rect 9815 13889 9827 13923
rect 9769 13883 9827 13889
rect 10042 13880 10048 13932
rect 10100 13880 10106 13932
rect 10318 13880 10324 13932
rect 10376 13920 10382 13932
rect 10413 13923 10471 13929
rect 10413 13920 10425 13923
rect 10376 13892 10425 13920
rect 10376 13880 10382 13892
rect 10413 13889 10425 13892
rect 10459 13889 10471 13923
rect 12621 13923 12679 13929
rect 10413 13883 10471 13889
rect 11348 13892 11928 13920
rect 9309 13855 9367 13861
rect 9309 13821 9321 13855
rect 9355 13821 9367 13855
rect 9309 13815 9367 13821
rect 9398 13812 9404 13864
rect 9456 13812 9462 13864
rect 9490 13812 9496 13864
rect 9548 13812 9554 13864
rect 9677 13855 9735 13861
rect 9677 13821 9689 13855
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 9953 13855 10011 13861
rect 9953 13821 9965 13855
rect 9999 13852 10011 13855
rect 10226 13852 10232 13864
rect 9999 13824 10232 13852
rect 9999 13821 10011 13824
rect 9953 13815 10011 13821
rect 5016 13787 5074 13793
rect 5016 13753 5028 13787
rect 5062 13784 5074 13787
rect 5353 13787 5411 13793
rect 5353 13784 5365 13787
rect 5062 13756 5365 13784
rect 5062 13753 5074 13756
rect 5016 13747 5074 13753
rect 5353 13753 5365 13756
rect 5399 13753 5411 13787
rect 5353 13747 5411 13753
rect 8202 13744 8208 13796
rect 8260 13744 8266 13796
rect 9692 13784 9720 13815
rect 10226 13812 10232 13824
rect 10284 13812 10290 13864
rect 10134 13784 10140 13796
rect 9692 13756 10140 13784
rect 10134 13744 10140 13756
rect 10192 13744 10198 13796
rect 10428 13784 10456 13883
rect 11241 13787 11299 13793
rect 11241 13784 11253 13787
rect 10428 13756 11253 13784
rect 11241 13753 11253 13756
rect 11287 13753 11299 13787
rect 11241 13747 11299 13753
rect 4706 13676 4712 13728
rect 4764 13716 4770 13728
rect 11348 13716 11376 13892
rect 11609 13855 11667 13861
rect 11609 13821 11621 13855
rect 11655 13821 11667 13855
rect 11609 13815 11667 13821
rect 11701 13855 11759 13861
rect 11701 13821 11713 13855
rect 11747 13852 11759 13855
rect 11790 13852 11796 13864
rect 11747 13824 11796 13852
rect 11747 13821 11759 13824
rect 11701 13815 11759 13821
rect 11624 13784 11652 13815
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 11900 13852 11928 13892
rect 12621 13889 12633 13923
rect 12667 13920 12679 13923
rect 12986 13920 12992 13932
rect 12667 13892 12992 13920
rect 12667 13889 12679 13892
rect 12621 13883 12679 13889
rect 12986 13880 12992 13892
rect 13044 13880 13050 13932
rect 13262 13880 13268 13932
rect 13320 13920 13326 13932
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 13320 13892 14013 13920
rect 13320 13880 13326 13892
rect 14001 13889 14013 13892
rect 14047 13920 14059 13923
rect 15102 13920 15108 13932
rect 14047 13892 15108 13920
rect 14047 13889 14059 13892
rect 14001 13883 14059 13889
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 15304 13929 15332 14028
rect 16298 14016 16304 14068
rect 16356 14056 16362 14068
rect 17126 14056 17132 14068
rect 16356 14028 17132 14056
rect 16356 14016 16362 14028
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 18141 14059 18199 14065
rect 17420 14028 18092 14056
rect 16390 13948 16396 14000
rect 16448 13988 16454 14000
rect 17310 13988 17316 14000
rect 16448 13960 17316 13988
rect 16448 13948 16454 13960
rect 17310 13948 17316 13960
rect 17368 13948 17374 14000
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13920 15347 13923
rect 15335 13892 15792 13920
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 11900 13824 15148 13852
rect 15120 13793 15148 13824
rect 15105 13787 15163 13793
rect 11624 13756 12020 13784
rect 4764 13688 11376 13716
rect 4764 13676 4770 13688
rect 11422 13676 11428 13728
rect 11480 13716 11486 13728
rect 11885 13719 11943 13725
rect 11885 13716 11897 13719
rect 11480 13688 11897 13716
rect 11480 13676 11486 13688
rect 11885 13685 11897 13688
rect 11931 13685 11943 13719
rect 11992 13716 12020 13756
rect 15105 13753 15117 13787
rect 15151 13753 15163 13787
rect 15764 13784 15792 13892
rect 16022 13880 16028 13932
rect 16080 13920 16086 13932
rect 17420 13920 17448 14028
rect 17497 13991 17555 13997
rect 17497 13957 17509 13991
rect 17543 13957 17555 13991
rect 18064 13988 18092 14028
rect 18141 14025 18153 14059
rect 18187 14056 18199 14059
rect 18322 14056 18328 14068
rect 18187 14028 18328 14056
rect 18187 14025 18199 14028
rect 18141 14019 18199 14025
rect 18322 14016 18328 14028
rect 18380 14016 18386 14068
rect 20898 14056 20904 14068
rect 19444 14028 20904 14056
rect 19444 13988 19472 14028
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 21174 14016 21180 14068
rect 21232 14016 21238 14068
rect 22370 14016 22376 14068
rect 22428 14016 22434 14068
rect 23474 14016 23480 14068
rect 23532 14056 23538 14068
rect 23845 14059 23903 14065
rect 23845 14056 23857 14059
rect 23532 14028 23857 14056
rect 23532 14016 23538 14028
rect 23845 14025 23857 14028
rect 23891 14056 23903 14059
rect 24026 14056 24032 14068
rect 23891 14028 24032 14056
rect 23891 14025 23903 14028
rect 23845 14019 23903 14025
rect 24026 14016 24032 14028
rect 24084 14016 24090 14068
rect 24320 14028 25360 14056
rect 18064 13960 19472 13988
rect 19521 13991 19579 13997
rect 17497 13951 17555 13957
rect 19521 13957 19533 13991
rect 19567 13957 19579 13991
rect 22388 13988 22416 14016
rect 24320 13988 24348 14028
rect 22388 13960 24348 13988
rect 19521 13951 19579 13957
rect 16080 13892 17448 13920
rect 17512 13920 17540 13951
rect 19536 13920 19564 13951
rect 17512 13892 18920 13920
rect 19536 13892 19932 13920
rect 16080 13880 16086 13892
rect 15838 13812 15844 13864
rect 15896 13852 15902 13864
rect 15896 13824 16804 13852
rect 15896 13812 15902 13824
rect 16666 13784 16672 13796
rect 15764 13756 16672 13784
rect 15105 13747 15163 13753
rect 16666 13744 16672 13756
rect 16724 13744 16730 13796
rect 16776 13784 16804 13824
rect 16850 13812 16856 13864
rect 16908 13852 16914 13864
rect 16945 13855 17003 13861
rect 16945 13852 16957 13855
rect 16908 13824 16957 13852
rect 16908 13812 16914 13824
rect 16945 13821 16957 13824
rect 16991 13821 17003 13855
rect 17221 13855 17279 13861
rect 17221 13852 17233 13855
rect 16945 13815 17003 13821
rect 17052 13824 17233 13852
rect 17052 13784 17080 13824
rect 17221 13821 17233 13824
rect 17267 13821 17279 13855
rect 17221 13815 17279 13821
rect 17310 13812 17316 13864
rect 17368 13812 17374 13864
rect 17420 13852 17448 13892
rect 17589 13855 17647 13861
rect 17589 13852 17601 13855
rect 17420 13824 17601 13852
rect 17589 13821 17601 13824
rect 17635 13821 17647 13855
rect 17957 13855 18015 13861
rect 17957 13852 17969 13855
rect 17589 13815 17647 13821
rect 17696 13824 17969 13852
rect 16776 13756 17080 13784
rect 17126 13744 17132 13796
rect 17184 13744 17190 13796
rect 17328 13784 17356 13812
rect 17696 13784 17724 13824
rect 17957 13821 17969 13824
rect 18003 13821 18015 13855
rect 17957 13815 18015 13821
rect 18230 13812 18236 13864
rect 18288 13852 18294 13864
rect 18690 13852 18696 13864
rect 18288 13824 18696 13852
rect 18288 13812 18294 13824
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 18892 13861 18920 13892
rect 18877 13855 18935 13861
rect 18877 13821 18889 13855
rect 18923 13821 18935 13855
rect 18877 13815 18935 13821
rect 19061 13855 19119 13861
rect 19061 13821 19073 13855
rect 19107 13852 19119 13855
rect 19337 13855 19395 13861
rect 19337 13852 19349 13855
rect 19107 13824 19349 13852
rect 19107 13821 19119 13824
rect 19061 13815 19119 13821
rect 19337 13821 19349 13824
rect 19383 13821 19395 13855
rect 19337 13815 19395 13821
rect 19794 13812 19800 13864
rect 19852 13812 19858 13864
rect 19904 13852 19932 13892
rect 21358 13880 21364 13932
rect 21416 13920 21422 13932
rect 21910 13920 21916 13932
rect 21416 13892 21916 13920
rect 21416 13880 21422 13892
rect 21910 13880 21916 13892
rect 21968 13880 21974 13932
rect 22370 13880 22376 13932
rect 22428 13880 22434 13932
rect 25222 13880 25228 13932
rect 25280 13880 25286 13932
rect 25332 13920 25360 14028
rect 25406 14016 25412 14068
rect 25464 14016 25470 14068
rect 25498 14016 25504 14068
rect 25556 14016 25562 14068
rect 25590 14016 25596 14068
rect 25648 14056 25654 14068
rect 25685 14059 25743 14065
rect 25685 14056 25697 14059
rect 25648 14028 25697 14056
rect 25648 14016 25654 14028
rect 25685 14025 25697 14028
rect 25731 14025 25743 14059
rect 25685 14019 25743 14025
rect 25593 13923 25651 13929
rect 25593 13920 25605 13923
rect 25332 13892 25605 13920
rect 25593 13889 25605 13892
rect 25639 13920 25651 13923
rect 25774 13920 25780 13932
rect 25639 13892 25780 13920
rect 25639 13889 25651 13892
rect 25593 13883 25651 13889
rect 25774 13880 25780 13892
rect 25832 13880 25838 13932
rect 20053 13855 20111 13861
rect 20053 13852 20065 13855
rect 19904 13824 20065 13852
rect 20053 13821 20065 13824
rect 20099 13821 20111 13855
rect 20053 13815 20111 13821
rect 21266 13812 21272 13864
rect 21324 13812 21330 13864
rect 21450 13812 21456 13864
rect 21508 13812 21514 13864
rect 21542 13812 21548 13864
rect 21600 13852 21606 13864
rect 21821 13855 21879 13861
rect 21821 13852 21833 13855
rect 21600 13824 21833 13852
rect 21600 13812 21606 13824
rect 21821 13821 21833 13824
rect 21867 13821 21879 13855
rect 21821 13815 21879 13821
rect 23290 13812 23296 13864
rect 23348 13852 23354 13864
rect 23348 13824 25084 13852
rect 23348 13812 23354 13824
rect 17328 13756 17724 13784
rect 17770 13744 17776 13796
rect 17828 13744 17834 13796
rect 17862 13744 17868 13796
rect 17920 13744 17926 13796
rect 24854 13744 24860 13796
rect 24912 13784 24918 13796
rect 24958 13787 25016 13793
rect 24958 13784 24970 13787
rect 24912 13756 24970 13784
rect 24912 13744 24918 13756
rect 24958 13753 24970 13756
rect 25004 13753 25016 13787
rect 25056 13784 25084 13824
rect 25130 13812 25136 13864
rect 25188 13852 25194 13864
rect 25317 13855 25375 13861
rect 25317 13852 25329 13855
rect 25188 13824 25329 13852
rect 25188 13812 25194 13824
rect 25317 13821 25329 13824
rect 25363 13821 25375 13855
rect 25317 13815 25375 13821
rect 25406 13812 25412 13864
rect 25464 13852 25470 13864
rect 25685 13855 25743 13861
rect 25685 13852 25697 13855
rect 25464 13824 25697 13852
rect 25464 13812 25470 13824
rect 25685 13821 25697 13824
rect 25731 13821 25743 13855
rect 25685 13815 25743 13821
rect 25866 13812 25872 13864
rect 25924 13812 25930 13864
rect 25590 13784 25596 13796
rect 25056 13756 25596 13784
rect 24958 13747 25016 13753
rect 25590 13744 25596 13756
rect 25648 13744 25654 13796
rect 12250 13716 12256 13728
rect 11992 13688 12256 13716
rect 11885 13679 11943 13685
rect 12250 13676 12256 13688
rect 12308 13716 12314 13728
rect 12345 13719 12403 13725
rect 12345 13716 12357 13719
rect 12308 13688 12357 13716
rect 12308 13676 12314 13688
rect 12345 13685 12357 13688
rect 12391 13685 12403 13719
rect 12345 13679 12403 13685
rect 12434 13676 12440 13728
rect 12492 13676 12498 13728
rect 14182 13676 14188 13728
rect 14240 13676 14246 13728
rect 14277 13719 14335 13725
rect 14277 13685 14289 13719
rect 14323 13716 14335 13719
rect 14366 13716 14372 13728
rect 14323 13688 14372 13716
rect 14323 13685 14335 13688
rect 14277 13679 14335 13685
rect 14366 13676 14372 13688
rect 14424 13676 14430 13728
rect 15197 13719 15255 13725
rect 15197 13685 15209 13719
rect 15243 13716 15255 13719
rect 16114 13716 16120 13728
rect 15243 13688 16120 13716
rect 15243 13685 15255 13688
rect 15197 13679 15255 13685
rect 16114 13676 16120 13688
rect 16172 13676 16178 13728
rect 17144 13716 17172 13744
rect 17788 13716 17816 13744
rect 17144 13688 17816 13716
rect 552 13626 27576 13648
rect 552 13574 7114 13626
rect 7166 13574 7178 13626
rect 7230 13574 7242 13626
rect 7294 13574 7306 13626
rect 7358 13574 7370 13626
rect 7422 13574 13830 13626
rect 13882 13574 13894 13626
rect 13946 13574 13958 13626
rect 14010 13574 14022 13626
rect 14074 13574 14086 13626
rect 14138 13574 20546 13626
rect 20598 13574 20610 13626
rect 20662 13574 20674 13626
rect 20726 13574 20738 13626
rect 20790 13574 20802 13626
rect 20854 13574 27262 13626
rect 27314 13574 27326 13626
rect 27378 13574 27390 13626
rect 27442 13574 27454 13626
rect 27506 13574 27518 13626
rect 27570 13574 27576 13626
rect 552 13552 27576 13574
rect 5445 13515 5503 13521
rect 5445 13481 5457 13515
rect 5491 13512 5503 13515
rect 5626 13512 5632 13524
rect 5491 13484 5632 13512
rect 5491 13481 5503 13484
rect 5445 13475 5503 13481
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 8941 13515 8999 13521
rect 8941 13481 8953 13515
rect 8987 13512 8999 13515
rect 9858 13512 9864 13524
rect 8987 13484 9864 13512
rect 8987 13481 8999 13484
rect 8941 13475 8999 13481
rect 9858 13472 9864 13484
rect 9916 13512 9922 13524
rect 10134 13512 10140 13524
rect 9916 13484 10140 13512
rect 9916 13472 9922 13484
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 13081 13515 13139 13521
rect 13081 13512 13093 13515
rect 12492 13484 13093 13512
rect 12492 13472 12498 13484
rect 13081 13481 13093 13484
rect 13127 13481 13139 13515
rect 13081 13475 13139 13481
rect 13446 13472 13452 13524
rect 13504 13472 13510 13524
rect 14182 13472 14188 13524
rect 14240 13512 14246 13524
rect 14553 13515 14611 13521
rect 14553 13512 14565 13515
rect 14240 13484 14565 13512
rect 14240 13472 14246 13484
rect 14553 13481 14565 13484
rect 14599 13481 14611 13515
rect 14553 13475 14611 13481
rect 24305 13515 24363 13521
rect 24305 13481 24317 13515
rect 24351 13512 24363 13515
rect 24854 13512 24860 13524
rect 24351 13484 24860 13512
rect 24351 13481 24363 13484
rect 24305 13475 24363 13481
rect 24854 13472 24860 13484
rect 24912 13472 24918 13524
rect 25225 13515 25283 13521
rect 25225 13481 25237 13515
rect 25271 13512 25283 13515
rect 25866 13512 25872 13524
rect 25271 13484 25872 13512
rect 25271 13481 25283 13484
rect 25225 13475 25283 13481
rect 25866 13472 25872 13484
rect 25924 13472 25930 13524
rect 4246 13404 4252 13456
rect 4304 13444 4310 13456
rect 4433 13447 4491 13453
rect 4433 13444 4445 13447
rect 4304 13416 4445 13444
rect 4304 13404 4310 13416
rect 4433 13413 4445 13416
rect 4479 13444 4491 13447
rect 9674 13444 9680 13456
rect 4479 13416 4844 13444
rect 4479 13413 4491 13416
rect 4433 13407 4491 13413
rect 4341 13379 4399 13385
rect 4341 13345 4353 13379
rect 4387 13376 4399 13379
rect 4525 13379 4583 13385
rect 4387 13348 4476 13376
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 4448 13320 4476 13348
rect 4525 13345 4537 13379
rect 4571 13345 4583 13379
rect 4525 13339 4583 13345
rect 4430 13268 4436 13320
rect 4488 13268 4494 13320
rect 4540 13308 4568 13339
rect 4706 13336 4712 13388
rect 4764 13336 4770 13388
rect 4816 13385 4844 13416
rect 7576 13416 9680 13444
rect 7576 13385 7604 13416
rect 9674 13404 9680 13416
rect 9732 13404 9738 13456
rect 9950 13404 9956 13456
rect 10008 13444 10014 13456
rect 11882 13444 11888 13456
rect 10008 13416 11888 13444
rect 10008 13404 10014 13416
rect 11882 13404 11888 13416
rect 11940 13444 11946 13456
rect 12713 13447 12771 13453
rect 11940 13416 12572 13444
rect 11940 13404 11946 13416
rect 4801 13379 4859 13385
rect 4801 13345 4813 13379
rect 4847 13345 4859 13379
rect 4801 13339 4859 13345
rect 7561 13379 7619 13385
rect 7561 13345 7573 13379
rect 7607 13345 7619 13379
rect 7561 13339 7619 13345
rect 7828 13379 7886 13385
rect 7828 13345 7840 13379
rect 7874 13376 7886 13379
rect 8386 13376 8392 13388
rect 7874 13348 8392 13376
rect 7874 13345 7886 13348
rect 7828 13339 7886 13345
rect 8386 13336 8392 13348
rect 8444 13336 8450 13388
rect 9217 13379 9275 13385
rect 9217 13345 9229 13379
rect 9263 13376 9275 13379
rect 10226 13376 10232 13388
rect 9263 13348 10232 13376
rect 9263 13345 9275 13348
rect 9217 13339 9275 13345
rect 10226 13336 10232 13348
rect 10284 13336 10290 13388
rect 11054 13336 11060 13388
rect 11112 13376 11118 13388
rect 11221 13379 11279 13385
rect 11221 13376 11233 13379
rect 11112 13348 11233 13376
rect 11112 13336 11118 13348
rect 11221 13345 11233 13348
rect 11267 13345 11279 13379
rect 11221 13339 11279 13345
rect 12434 13336 12440 13388
rect 12492 13336 12498 13388
rect 4890 13308 4896 13320
rect 4540 13280 4896 13308
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 4982 13268 4988 13320
rect 5040 13308 5046 13320
rect 6365 13311 6423 13317
rect 6365 13308 6377 13311
rect 5040 13280 6377 13308
rect 5040 13268 5046 13280
rect 6365 13277 6377 13280
rect 6411 13277 6423 13311
rect 6365 13271 6423 13277
rect 8754 13268 8760 13320
rect 8812 13308 8818 13320
rect 9309 13311 9367 13317
rect 8812 13280 9260 13308
rect 8812 13268 8818 13280
rect 9033 13243 9091 13249
rect 9033 13240 9045 13243
rect 8496 13212 9045 13240
rect 4154 13132 4160 13184
rect 4212 13132 4218 13184
rect 5813 13175 5871 13181
rect 5813 13141 5825 13175
rect 5859 13172 5871 13175
rect 6086 13172 6092 13184
rect 5859 13144 6092 13172
rect 5859 13141 5871 13144
rect 5813 13135 5871 13141
rect 6086 13132 6092 13144
rect 6144 13132 6150 13184
rect 7926 13132 7932 13184
rect 7984 13172 7990 13184
rect 8496 13172 8524 13212
rect 9033 13209 9045 13212
rect 9079 13209 9091 13243
rect 9232 13240 9260 13280
rect 9309 13277 9321 13311
rect 9355 13308 9367 13311
rect 9398 13308 9404 13320
rect 9355 13280 9404 13308
rect 9355 13277 9367 13280
rect 9309 13271 9367 13277
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 9692 13240 9720 13271
rect 10962 13268 10968 13320
rect 11020 13268 11026 13320
rect 12544 13308 12572 13416
rect 12713 13413 12725 13447
rect 12759 13444 12771 13447
rect 12759 13416 12940 13444
rect 12759 13413 12771 13416
rect 12713 13407 12771 13413
rect 12618 13336 12624 13388
rect 12676 13336 12682 13388
rect 12805 13379 12863 13385
rect 12805 13345 12817 13379
rect 12851 13345 12863 13379
rect 12805 13339 12863 13345
rect 12820 13308 12848 13339
rect 12544 13280 12848 13308
rect 9232 13212 9720 13240
rect 9033 13203 9091 13209
rect 7984 13144 8524 13172
rect 9692 13172 9720 13212
rect 12342 13200 12348 13252
rect 12400 13240 12406 13252
rect 12912 13240 12940 13416
rect 13538 13404 13544 13456
rect 13596 13444 13602 13456
rect 13596 13416 16252 13444
rect 13596 13404 13602 13416
rect 14921 13379 14979 13385
rect 14921 13345 14933 13379
rect 14967 13376 14979 13379
rect 15194 13376 15200 13388
rect 14967 13348 15200 13376
rect 14967 13345 14979 13348
rect 14921 13339 14979 13345
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 16114 13336 16120 13388
rect 16172 13336 16178 13388
rect 16224 13376 16252 13416
rect 16298 13404 16304 13456
rect 16356 13404 16362 13456
rect 16666 13404 16672 13456
rect 16724 13444 16730 13456
rect 16724 13416 17540 13444
rect 16724 13404 16730 13416
rect 16393 13379 16451 13385
rect 16393 13376 16405 13379
rect 16224 13348 16405 13376
rect 16393 13345 16405 13348
rect 16439 13345 16451 13379
rect 16393 13339 16451 13345
rect 16482 13336 16488 13388
rect 16540 13336 16546 13388
rect 17512 13385 17540 13416
rect 21542 13404 21548 13456
rect 21600 13404 21606 13456
rect 25593 13447 25651 13453
rect 25593 13444 25605 13447
rect 24780 13416 25605 13444
rect 16945 13379 17003 13385
rect 16945 13345 16957 13379
rect 16991 13345 17003 13379
rect 16945 13339 17003 13345
rect 17497 13379 17555 13385
rect 17497 13345 17509 13379
rect 17543 13345 17555 13379
rect 17497 13339 17555 13345
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13277 13599 13311
rect 13541 13271 13599 13277
rect 12400 13212 12940 13240
rect 13556 13240 13584 13271
rect 13722 13268 13728 13320
rect 13780 13268 13786 13320
rect 14550 13268 14556 13320
rect 14608 13308 14614 13320
rect 15013 13311 15071 13317
rect 15013 13308 15025 13311
rect 14608 13280 15025 13308
rect 14608 13268 14614 13280
rect 15013 13277 15025 13280
rect 15059 13277 15071 13311
rect 15013 13271 15071 13277
rect 15102 13268 15108 13320
rect 15160 13268 15166 13320
rect 16574 13240 16580 13252
rect 13556 13212 16580 13240
rect 12400 13200 12406 13212
rect 16574 13200 16580 13212
rect 16632 13200 16638 13252
rect 16669 13243 16727 13249
rect 16669 13209 16681 13243
rect 16715 13240 16727 13243
rect 16960 13240 16988 13339
rect 20898 13336 20904 13388
rect 20956 13376 20962 13388
rect 21453 13379 21511 13385
rect 21453 13376 21465 13379
rect 20956 13348 21465 13376
rect 20956 13336 20962 13348
rect 21453 13345 21465 13348
rect 21499 13345 21511 13379
rect 21560 13376 21588 13404
rect 21821 13379 21879 13385
rect 21821 13376 21833 13379
rect 21560 13348 21833 13376
rect 21453 13339 21511 13345
rect 21821 13345 21833 13348
rect 21867 13345 21879 13379
rect 21821 13339 21879 13345
rect 24026 13336 24032 13388
rect 24084 13336 24090 13388
rect 24780 13385 24808 13416
rect 25593 13413 25605 13416
rect 25639 13413 25651 13447
rect 25593 13407 25651 13413
rect 24765 13379 24823 13385
rect 24765 13345 24777 13379
rect 24811 13345 24823 13379
rect 24765 13339 24823 13345
rect 25038 13336 25044 13388
rect 25096 13336 25102 13388
rect 25133 13379 25191 13385
rect 25133 13345 25145 13379
rect 25179 13345 25191 13379
rect 25133 13339 25191 13345
rect 17129 13311 17187 13317
rect 17129 13277 17141 13311
rect 17175 13277 17187 13311
rect 17129 13271 17187 13277
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13308 17831 13311
rect 17862 13308 17868 13320
rect 17819 13280 17868 13308
rect 17819 13277 17831 13280
rect 17773 13271 17831 13277
rect 16715 13212 16988 13240
rect 17144 13240 17172 13271
rect 17862 13268 17868 13280
rect 17920 13268 17926 13320
rect 21266 13268 21272 13320
rect 21324 13308 21330 13320
rect 21545 13311 21603 13317
rect 21545 13308 21557 13311
rect 21324 13280 21557 13308
rect 21324 13268 21330 13280
rect 21545 13277 21557 13280
rect 21591 13277 21603 13311
rect 21545 13271 21603 13277
rect 21729 13311 21787 13317
rect 21729 13277 21741 13311
rect 21775 13308 21787 13311
rect 22278 13308 22284 13320
rect 21775 13280 22284 13308
rect 21775 13277 21787 13280
rect 21729 13271 21787 13277
rect 18690 13240 18696 13252
rect 17144 13212 18696 13240
rect 16715 13209 16727 13212
rect 16669 13203 16727 13209
rect 18690 13200 18696 13212
rect 18748 13200 18754 13252
rect 21082 13200 21088 13252
rect 21140 13240 21146 13252
rect 21744 13240 21772 13271
rect 22278 13268 22284 13280
rect 22336 13268 22342 13320
rect 22465 13311 22523 13317
rect 22465 13277 22477 13311
rect 22511 13308 22523 13311
rect 22554 13308 22560 13320
rect 22511 13280 22560 13308
rect 22511 13277 22523 13280
rect 22465 13271 22523 13277
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 23750 13268 23756 13320
rect 23808 13308 23814 13320
rect 23845 13311 23903 13317
rect 23845 13308 23857 13311
rect 23808 13280 23857 13308
rect 23808 13268 23814 13280
rect 23845 13277 23857 13280
rect 23891 13277 23903 13311
rect 23845 13271 23903 13277
rect 23937 13311 23995 13317
rect 23937 13277 23949 13311
rect 23983 13277 23995 13311
rect 23937 13271 23995 13277
rect 24121 13311 24179 13317
rect 24121 13277 24133 13311
rect 24167 13308 24179 13311
rect 24302 13308 24308 13320
rect 24167 13280 24308 13308
rect 24167 13277 24179 13280
rect 24121 13271 24179 13277
rect 21140 13212 21772 13240
rect 23952 13240 23980 13271
rect 24302 13268 24308 13280
rect 24360 13268 24366 13320
rect 24946 13268 24952 13320
rect 25004 13308 25010 13320
rect 25148 13308 25176 13339
rect 25406 13336 25412 13388
rect 25464 13336 25470 13388
rect 25608 13376 25636 13407
rect 25685 13379 25743 13385
rect 25685 13376 25697 13379
rect 25608 13348 25697 13376
rect 25685 13345 25697 13348
rect 25731 13345 25743 13379
rect 25685 13339 25743 13345
rect 25774 13336 25780 13388
rect 25832 13376 25838 13388
rect 25869 13379 25927 13385
rect 25869 13376 25881 13379
rect 25832 13348 25881 13376
rect 25832 13336 25838 13348
rect 25869 13345 25881 13348
rect 25915 13345 25927 13379
rect 25869 13339 25927 13345
rect 25314 13308 25320 13320
rect 25004 13280 25320 13308
rect 25004 13268 25010 13280
rect 25314 13268 25320 13280
rect 25372 13268 25378 13320
rect 25866 13240 25872 13252
rect 23952 13212 25872 13240
rect 21140 13200 21146 13212
rect 25866 13200 25872 13212
rect 25924 13200 25930 13252
rect 11330 13172 11336 13184
rect 9692 13144 11336 13172
rect 7984 13132 7990 13144
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 12710 13132 12716 13184
rect 12768 13172 12774 13184
rect 12989 13175 13047 13181
rect 12989 13172 13001 13175
rect 12768 13144 13001 13172
rect 12768 13132 12774 13144
rect 12989 13141 13001 13144
rect 13035 13141 13047 13175
rect 12989 13135 13047 13141
rect 15930 13132 15936 13184
rect 15988 13172 15994 13184
rect 16761 13175 16819 13181
rect 16761 13172 16773 13175
rect 15988 13144 16773 13172
rect 15988 13132 15994 13144
rect 16761 13141 16773 13144
rect 16807 13141 16819 13175
rect 16761 13135 16819 13141
rect 24581 13175 24639 13181
rect 24581 13141 24593 13175
rect 24627 13172 24639 13175
rect 24762 13172 24768 13184
rect 24627 13144 24768 13172
rect 24627 13141 24639 13144
rect 24581 13135 24639 13141
rect 24762 13132 24768 13144
rect 24820 13132 24826 13184
rect 24946 13132 24952 13184
rect 25004 13132 25010 13184
rect 25774 13132 25780 13184
rect 25832 13132 25838 13184
rect 552 13082 27416 13104
rect 552 13030 3756 13082
rect 3808 13030 3820 13082
rect 3872 13030 3884 13082
rect 3936 13030 3948 13082
rect 4000 13030 4012 13082
rect 4064 13030 10472 13082
rect 10524 13030 10536 13082
rect 10588 13030 10600 13082
rect 10652 13030 10664 13082
rect 10716 13030 10728 13082
rect 10780 13030 17188 13082
rect 17240 13030 17252 13082
rect 17304 13030 17316 13082
rect 17368 13030 17380 13082
rect 17432 13030 17444 13082
rect 17496 13030 23904 13082
rect 23956 13030 23968 13082
rect 24020 13030 24032 13082
rect 24084 13030 24096 13082
rect 24148 13030 24160 13082
rect 24212 13030 27416 13082
rect 552 13008 27416 13030
rect 4982 12928 4988 12980
rect 5040 12928 5046 12980
rect 6914 12928 6920 12980
rect 6972 12928 6978 12980
rect 8386 12928 8392 12980
rect 8444 12928 8450 12980
rect 10965 12971 11023 12977
rect 10965 12937 10977 12971
rect 11011 12968 11023 12971
rect 11054 12968 11060 12980
rect 11011 12940 11060 12968
rect 11011 12937 11023 12940
rect 10965 12931 11023 12937
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 13446 12968 13452 12980
rect 12492 12940 13452 12968
rect 12492 12928 12498 12940
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 17589 12971 17647 12977
rect 17589 12968 17601 12971
rect 16172 12940 17601 12968
rect 16172 12928 16178 12940
rect 17589 12937 17601 12940
rect 17635 12968 17647 12971
rect 17678 12968 17684 12980
rect 17635 12940 17684 12968
rect 17635 12937 17647 12940
rect 17589 12931 17647 12937
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 20438 12968 20444 12980
rect 17788 12940 20444 12968
rect 3697 12835 3755 12841
rect 3697 12832 3709 12835
rect 3068 12804 3709 12832
rect 3068 12773 3096 12804
rect 3697 12801 3709 12804
rect 3743 12801 3755 12835
rect 4154 12832 4160 12844
rect 3697 12795 3755 12801
rect 3896 12804 4160 12832
rect 3053 12767 3111 12773
rect 3053 12733 3065 12767
rect 3099 12733 3111 12767
rect 3053 12727 3111 12733
rect 3421 12767 3479 12773
rect 3421 12733 3433 12767
rect 3467 12733 3479 12767
rect 3421 12727 3479 12733
rect 3436 12696 3464 12727
rect 3602 12724 3608 12776
rect 3660 12724 3666 12776
rect 3896 12773 3924 12804
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 5000 12832 5028 12928
rect 4540 12804 5028 12832
rect 6365 12835 6423 12841
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12733 3939 12767
rect 3881 12727 3939 12733
rect 3970 12724 3976 12776
rect 4028 12724 4034 12776
rect 4430 12724 4436 12776
rect 4488 12724 4494 12776
rect 4540 12773 4568 12804
rect 6365 12801 6377 12835
rect 6411 12832 6423 12835
rect 6932 12832 6960 12928
rect 15194 12900 15200 12912
rect 6411 12804 6960 12832
rect 7392 12872 15200 12900
rect 6411 12801 6423 12804
rect 6365 12795 6423 12801
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12733 4583 12767
rect 4525 12727 4583 12733
rect 4801 12767 4859 12773
rect 4801 12733 4813 12767
rect 4847 12764 4859 12767
rect 5350 12764 5356 12776
rect 4847 12736 5356 12764
rect 4847 12733 4859 12736
rect 4801 12727 4859 12733
rect 5350 12724 5356 12736
rect 5408 12764 5414 12776
rect 7392 12764 7420 12872
rect 15194 12860 15200 12872
rect 15252 12860 15258 12912
rect 17494 12860 17500 12912
rect 17552 12900 17558 12912
rect 17788 12900 17816 12940
rect 20438 12928 20444 12940
rect 20496 12968 20502 12980
rect 20533 12971 20591 12977
rect 20533 12968 20545 12971
rect 20496 12940 20545 12968
rect 20496 12928 20502 12940
rect 20533 12937 20545 12940
rect 20579 12937 20591 12971
rect 20533 12931 20591 12937
rect 23750 12928 23756 12980
rect 23808 12968 23814 12980
rect 23937 12971 23995 12977
rect 23937 12968 23949 12971
rect 23808 12940 23949 12968
rect 23808 12928 23814 12940
rect 23937 12937 23949 12940
rect 23983 12937 23995 12971
rect 23937 12931 23995 12937
rect 24121 12971 24179 12977
rect 24121 12937 24133 12971
rect 24167 12937 24179 12971
rect 24121 12931 24179 12937
rect 17552 12872 17816 12900
rect 18233 12903 18291 12909
rect 17552 12860 17558 12872
rect 18233 12869 18245 12903
rect 18279 12900 18291 12903
rect 18598 12900 18604 12912
rect 18279 12872 18604 12900
rect 18279 12869 18291 12872
rect 18233 12863 18291 12869
rect 18598 12860 18604 12872
rect 18656 12860 18662 12912
rect 18708 12872 19196 12900
rect 8202 12792 8208 12844
rect 8260 12792 8266 12844
rect 9398 12792 9404 12844
rect 9456 12832 9462 12844
rect 9456 12804 12020 12832
rect 9456 12792 9462 12804
rect 5408 12736 7420 12764
rect 8220 12764 8248 12792
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 8220 12736 8585 12764
rect 5408 12724 5414 12736
rect 8573 12733 8585 12736
rect 8619 12733 8631 12767
rect 8573 12727 8631 12733
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 4617 12699 4675 12705
rect 3436 12668 4292 12696
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 2869 12631 2927 12637
rect 2869 12628 2881 12631
rect 2832 12600 2881 12628
rect 2832 12588 2838 12600
rect 2869 12597 2881 12600
rect 2915 12597 2927 12631
rect 2869 12591 2927 12597
rect 3234 12588 3240 12640
rect 3292 12588 3298 12640
rect 4264 12637 4292 12668
rect 4617 12665 4629 12699
rect 4663 12696 4675 12699
rect 4890 12696 4896 12708
rect 4663 12668 4896 12696
rect 4663 12665 4675 12668
rect 4617 12659 4675 12665
rect 4890 12656 4896 12668
rect 4948 12656 4954 12708
rect 5810 12656 5816 12708
rect 5868 12696 5874 12708
rect 6098 12699 6156 12705
rect 6098 12696 6110 12699
rect 5868 12668 6110 12696
rect 5868 12656 5874 12668
rect 6098 12665 6110 12668
rect 6144 12665 6156 12699
rect 6098 12659 6156 12665
rect 8202 12656 8208 12708
rect 8260 12656 8266 12708
rect 4249 12631 4307 12637
rect 4249 12597 4261 12631
rect 4295 12597 4307 12631
rect 9508 12628 9536 12727
rect 9582 12724 9588 12776
rect 9640 12764 9646 12776
rect 9784 12773 9812 12804
rect 9677 12767 9735 12773
rect 9677 12764 9689 12767
rect 9640 12736 9689 12764
rect 9640 12724 9646 12736
rect 9677 12733 9689 12736
rect 9723 12733 9735 12767
rect 9677 12727 9735 12733
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12733 9827 12767
rect 9769 12727 9827 12733
rect 9861 12767 9919 12773
rect 9861 12733 9873 12767
rect 9907 12764 9919 12767
rect 9950 12764 9956 12776
rect 9907 12736 9956 12764
rect 9907 12733 9919 12736
rect 9861 12727 9919 12733
rect 9950 12724 9956 12736
rect 10008 12724 10014 12776
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 10060 12736 10333 12764
rect 9950 12628 9956 12640
rect 9508 12600 9956 12628
rect 4249 12591 4307 12597
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10060 12637 10088 12736
rect 10321 12733 10333 12736
rect 10367 12733 10379 12767
rect 10321 12727 10379 12733
rect 10502 12724 10508 12776
rect 10560 12724 10566 12776
rect 11241 12767 11299 12773
rect 11241 12733 11253 12767
rect 11287 12733 11299 12767
rect 11241 12727 11299 12733
rect 11256 12696 11284 12727
rect 11330 12724 11336 12776
rect 11388 12724 11394 12776
rect 11422 12724 11428 12776
rect 11480 12724 11486 12776
rect 11609 12767 11667 12773
rect 11609 12733 11621 12767
rect 11655 12764 11667 12767
rect 11698 12764 11704 12776
rect 11655 12736 11704 12764
rect 11655 12733 11667 12736
rect 11609 12727 11667 12733
rect 11698 12724 11704 12736
rect 11756 12724 11762 12776
rect 11793 12699 11851 12705
rect 11793 12696 11805 12699
rect 11256 12668 11805 12696
rect 11793 12665 11805 12668
rect 11839 12665 11851 12699
rect 11992 12696 12020 12804
rect 12342 12792 12348 12844
rect 12400 12792 12406 12844
rect 12526 12792 12532 12844
rect 12584 12792 12590 12844
rect 16209 12835 16267 12841
rect 16209 12801 16221 12835
rect 16255 12832 16267 12835
rect 18708 12832 18736 12872
rect 19168 12841 19196 12872
rect 23474 12860 23480 12912
rect 23532 12900 23538 12912
rect 24136 12900 24164 12931
rect 24946 12928 24952 12980
rect 25004 12968 25010 12980
rect 25133 12971 25191 12977
rect 25133 12968 25145 12971
rect 25004 12940 25145 12968
rect 25004 12928 25010 12940
rect 25133 12937 25145 12940
rect 25179 12937 25191 12971
rect 25133 12931 25191 12937
rect 23532 12872 24164 12900
rect 23532 12860 23538 12872
rect 25038 12860 25044 12912
rect 25096 12900 25102 12912
rect 25406 12900 25412 12912
rect 25096 12872 25412 12900
rect 25096 12860 25102 12872
rect 25406 12860 25412 12872
rect 25464 12860 25470 12912
rect 16255 12804 16344 12832
rect 16255 12801 16267 12804
rect 16209 12795 16267 12801
rect 16316 12776 16344 12804
rect 17604 12804 18736 12832
rect 19153 12835 19211 12841
rect 12710 12724 12716 12776
rect 12768 12724 12774 12776
rect 12897 12767 12955 12773
rect 12897 12733 12909 12767
rect 12943 12764 12955 12767
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12943 12736 13001 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 12989 12733 13001 12736
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 15102 12764 15108 12776
rect 14875 12736 15108 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 15930 12724 15936 12776
rect 15988 12724 15994 12776
rect 16298 12724 16304 12776
rect 16356 12764 16362 12776
rect 17604 12764 17632 12804
rect 19153 12801 19165 12835
rect 19199 12801 19211 12835
rect 19153 12795 19211 12801
rect 16356 12736 17632 12764
rect 17681 12767 17739 12773
rect 16356 12724 16362 12736
rect 17681 12733 17693 12767
rect 17727 12733 17739 12767
rect 17681 12727 17739 12733
rect 14366 12696 14372 12708
rect 11992 12668 14372 12696
rect 11793 12659 11851 12665
rect 14366 12656 14372 12668
rect 14424 12656 14430 12708
rect 16465 12699 16523 12705
rect 16465 12665 16477 12699
rect 16511 12665 16523 12699
rect 16465 12659 16523 12665
rect 10045 12631 10103 12637
rect 10045 12597 10057 12631
rect 10091 12597 10103 12631
rect 10045 12591 10103 12597
rect 10134 12588 10140 12640
rect 10192 12588 10198 12640
rect 10226 12588 10232 12640
rect 10284 12628 10290 12640
rect 12986 12628 12992 12640
rect 10284 12600 12992 12628
rect 10284 12588 10290 12600
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 13173 12631 13231 12637
rect 13173 12597 13185 12631
rect 13219 12628 13231 12631
rect 13446 12628 13452 12640
rect 13219 12600 13452 12628
rect 13219 12597 13231 12600
rect 13173 12591 13231 12597
rect 13446 12588 13452 12600
rect 13504 12588 13510 12640
rect 14182 12588 14188 12640
rect 14240 12628 14246 12640
rect 14737 12631 14795 12637
rect 14737 12628 14749 12631
rect 14240 12600 14749 12628
rect 14240 12588 14246 12600
rect 14737 12597 14749 12600
rect 14783 12597 14795 12631
rect 14737 12591 14795 12597
rect 16117 12631 16175 12637
rect 16117 12597 16129 12631
rect 16163 12628 16175 12631
rect 16469 12628 16497 12659
rect 16574 12656 16580 12708
rect 16632 12696 16638 12708
rect 17494 12696 17500 12708
rect 16632 12668 17500 12696
rect 16632 12656 16638 12668
rect 17494 12656 17500 12668
rect 17552 12696 17558 12708
rect 17696 12696 17724 12727
rect 17770 12724 17776 12776
rect 17828 12764 17834 12776
rect 17865 12767 17923 12773
rect 17865 12764 17877 12767
rect 17828 12736 17877 12764
rect 17828 12724 17834 12736
rect 17865 12733 17877 12736
rect 17911 12733 17923 12767
rect 17865 12727 17923 12733
rect 18046 12724 18052 12776
rect 18104 12724 18110 12776
rect 18230 12724 18236 12776
rect 18288 12764 18294 12776
rect 18690 12764 18696 12776
rect 18288 12736 18696 12764
rect 18288 12724 18294 12736
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 18782 12724 18788 12776
rect 18840 12764 18846 12776
rect 18877 12767 18935 12773
rect 18877 12764 18889 12767
rect 18840 12736 18889 12764
rect 18840 12724 18846 12736
rect 18877 12733 18889 12736
rect 18923 12733 18935 12767
rect 19168 12764 19196 12795
rect 20990 12792 20996 12844
rect 21048 12832 21054 12844
rect 21266 12832 21272 12844
rect 21048 12804 21272 12832
rect 21048 12792 21054 12804
rect 21266 12792 21272 12804
rect 21324 12792 21330 12844
rect 21450 12792 21456 12844
rect 21508 12832 21514 12844
rect 22462 12832 22468 12844
rect 21508 12804 22468 12832
rect 21508 12792 21514 12804
rect 22462 12792 22468 12804
rect 22520 12792 22526 12844
rect 23569 12835 23627 12841
rect 23569 12801 23581 12835
rect 23615 12832 23627 12835
rect 25130 12832 25136 12844
rect 23615 12804 25136 12832
rect 23615 12801 23627 12804
rect 23569 12795 23627 12801
rect 25130 12792 25136 12804
rect 25188 12792 25194 12844
rect 25222 12792 25228 12844
rect 25280 12832 25286 12844
rect 25501 12835 25559 12841
rect 25501 12832 25513 12835
rect 25280 12804 25513 12832
rect 25280 12792 25286 12804
rect 25501 12801 25513 12804
rect 25547 12801 25559 12835
rect 25501 12795 25559 12801
rect 19794 12764 19800 12776
rect 19168 12736 19800 12764
rect 18877 12727 18935 12733
rect 19794 12724 19800 12736
rect 19852 12764 19858 12776
rect 19978 12764 19984 12776
rect 19852 12736 19984 12764
rect 19852 12724 19858 12736
rect 19978 12724 19984 12736
rect 20036 12724 20042 12776
rect 21174 12724 21180 12776
rect 21232 12724 21238 12776
rect 21542 12724 21548 12776
rect 21600 12724 21606 12776
rect 23477 12767 23535 12773
rect 23477 12764 23489 12767
rect 22066 12736 23489 12764
rect 17552 12668 17724 12696
rect 17957 12699 18015 12705
rect 17552 12656 17558 12668
rect 17957 12665 17969 12699
rect 18003 12696 18015 12699
rect 18138 12696 18144 12708
rect 18003 12668 18144 12696
rect 18003 12665 18015 12668
rect 17957 12659 18015 12665
rect 18138 12656 18144 12668
rect 18196 12656 18202 12708
rect 19426 12705 19432 12708
rect 18248 12668 19196 12696
rect 16163 12600 16497 12628
rect 16163 12597 16175 12600
rect 16117 12591 16175 12597
rect 16942 12588 16948 12640
rect 17000 12628 17006 12640
rect 18248 12628 18276 12668
rect 17000 12600 18276 12628
rect 17000 12588 17006 12600
rect 18966 12588 18972 12640
rect 19024 12628 19030 12640
rect 19061 12631 19119 12637
rect 19061 12628 19073 12631
rect 19024 12600 19073 12628
rect 19024 12588 19030 12600
rect 19061 12597 19073 12600
rect 19107 12597 19119 12631
rect 19168 12628 19196 12668
rect 19420 12659 19432 12705
rect 19426 12656 19432 12659
rect 19484 12656 19490 12708
rect 22066 12628 22094 12736
rect 23477 12733 23489 12736
rect 23523 12733 23535 12767
rect 23477 12727 23535 12733
rect 23661 12767 23719 12773
rect 23661 12733 23673 12767
rect 23707 12764 23719 12767
rect 23750 12764 23756 12776
rect 23707 12736 23756 12764
rect 23707 12733 23719 12736
rect 23661 12727 23719 12733
rect 23750 12724 23756 12736
rect 23808 12764 23814 12776
rect 24489 12767 24547 12773
rect 24489 12764 24501 12767
rect 23808 12736 24501 12764
rect 23808 12724 23814 12736
rect 24489 12733 24501 12736
rect 24535 12764 24547 12767
rect 25317 12767 25375 12773
rect 25317 12764 25329 12767
rect 24535 12736 25329 12764
rect 24535 12733 24547 12736
rect 24489 12727 24547 12733
rect 25317 12733 25329 12736
rect 25363 12733 25375 12767
rect 25317 12727 25375 12733
rect 25406 12724 25412 12776
rect 25464 12724 25470 12776
rect 25774 12773 25780 12776
rect 25768 12764 25780 12773
rect 25735 12736 25780 12764
rect 25768 12727 25780 12736
rect 25774 12724 25780 12727
rect 25832 12724 25838 12776
rect 22189 12699 22247 12705
rect 22189 12665 22201 12699
rect 22235 12696 22247 12699
rect 23290 12696 23296 12708
rect 22235 12668 23296 12696
rect 22235 12665 22247 12668
rect 22189 12659 22247 12665
rect 23290 12656 23296 12668
rect 23348 12656 23354 12708
rect 24305 12699 24363 12705
rect 24305 12665 24317 12699
rect 24351 12696 24363 12699
rect 24394 12696 24400 12708
rect 24351 12668 24400 12696
rect 24351 12665 24363 12668
rect 24305 12659 24363 12665
rect 24394 12656 24400 12668
rect 24452 12656 24458 12708
rect 25133 12699 25191 12705
rect 25133 12665 25145 12699
rect 25179 12696 25191 12699
rect 25590 12696 25596 12708
rect 25179 12668 25596 12696
rect 25179 12665 25191 12668
rect 25133 12659 25191 12665
rect 25590 12656 25596 12668
rect 25648 12656 25654 12708
rect 19168 12600 22094 12628
rect 19061 12591 19119 12597
rect 23658 12588 23664 12640
rect 23716 12628 23722 12640
rect 24095 12631 24153 12637
rect 24095 12628 24107 12631
rect 23716 12600 24107 12628
rect 23716 12588 23722 12600
rect 24095 12597 24107 12600
rect 24141 12597 24153 12631
rect 24095 12591 24153 12597
rect 25038 12588 25044 12640
rect 25096 12588 25102 12640
rect 25314 12588 25320 12640
rect 25372 12628 25378 12640
rect 25866 12628 25872 12640
rect 25372 12600 25872 12628
rect 25372 12588 25378 12600
rect 25866 12588 25872 12600
rect 25924 12588 25930 12640
rect 26878 12588 26884 12640
rect 26936 12588 26942 12640
rect 552 12538 27576 12560
rect 552 12486 7114 12538
rect 7166 12486 7178 12538
rect 7230 12486 7242 12538
rect 7294 12486 7306 12538
rect 7358 12486 7370 12538
rect 7422 12486 13830 12538
rect 13882 12486 13894 12538
rect 13946 12486 13958 12538
rect 14010 12486 14022 12538
rect 14074 12486 14086 12538
rect 14138 12486 20546 12538
rect 20598 12486 20610 12538
rect 20662 12486 20674 12538
rect 20726 12486 20738 12538
rect 20790 12486 20802 12538
rect 20854 12486 27262 12538
rect 27314 12486 27326 12538
rect 27378 12486 27390 12538
rect 27442 12486 27454 12538
rect 27506 12486 27518 12538
rect 27570 12486 27576 12538
rect 552 12464 27576 12486
rect 5350 12384 5356 12436
rect 5408 12384 5414 12436
rect 5810 12384 5816 12436
rect 5868 12384 5874 12436
rect 8849 12427 8907 12433
rect 8849 12393 8861 12427
rect 8895 12393 8907 12427
rect 8849 12387 8907 12393
rect 2516 12328 4016 12356
rect 2516 12232 2544 12328
rect 2774 12297 2780 12300
rect 2768 12251 2780 12297
rect 2832 12288 2838 12300
rect 3988 12297 4016 12328
rect 5718 12316 5724 12368
rect 5776 12356 5782 12368
rect 7926 12356 7932 12368
rect 5776 12328 6224 12356
rect 5776 12316 5782 12328
rect 4246 12297 4252 12300
rect 3973 12291 4031 12297
rect 2832 12260 2868 12288
rect 2774 12248 2780 12251
rect 2832 12248 2838 12260
rect 3973 12257 3985 12291
rect 4019 12257 4031 12291
rect 3973 12251 4031 12257
rect 4240 12251 4252 12297
rect 4246 12248 4252 12251
rect 4304 12248 4310 12300
rect 6086 12248 6092 12300
rect 6144 12248 6150 12300
rect 6196 12297 6224 12328
rect 6288 12328 7932 12356
rect 6288 12297 6316 12328
rect 7926 12316 7932 12328
rect 7984 12316 7990 12368
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12257 6239 12291
rect 6181 12251 6239 12257
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12257 6331 12291
rect 6273 12251 6331 12257
rect 6454 12248 6460 12300
rect 6512 12248 6518 12300
rect 7834 12248 7840 12300
rect 7892 12248 7898 12300
rect 8018 12248 8024 12300
rect 8076 12248 8082 12300
rect 8389 12291 8447 12297
rect 8389 12257 8401 12291
rect 8435 12288 8447 12291
rect 8478 12288 8484 12300
rect 8435 12260 8484 12288
rect 8435 12257 8447 12260
rect 8389 12251 8447 12257
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 8665 12291 8723 12297
rect 8665 12257 8677 12291
rect 8711 12257 8723 12291
rect 8864 12288 8892 12387
rect 10962 12384 10968 12436
rect 11020 12424 11026 12436
rect 12253 12427 12311 12433
rect 12253 12424 12265 12427
rect 11020 12396 12265 12424
rect 11020 12384 11026 12396
rect 12253 12393 12265 12396
rect 12299 12393 12311 12427
rect 14550 12424 14556 12436
rect 12253 12387 12311 12393
rect 12406 12396 14556 12424
rect 8938 12316 8944 12368
rect 8996 12356 9002 12368
rect 9674 12356 9680 12368
rect 8996 12328 9680 12356
rect 8996 12316 9002 12328
rect 9674 12316 9680 12328
rect 9732 12356 9738 12368
rect 10980 12356 11008 12384
rect 12406 12356 12434 12396
rect 14550 12384 14556 12396
rect 14608 12384 14614 12436
rect 14918 12384 14924 12436
rect 14976 12424 14982 12436
rect 15102 12424 15108 12436
rect 14976 12396 15108 12424
rect 14976 12384 14982 12396
rect 15102 12384 15108 12396
rect 15160 12424 15166 12436
rect 15160 12396 17908 12424
rect 15160 12384 15166 12396
rect 14182 12356 14188 12368
rect 9732 12328 11008 12356
rect 11072 12328 12434 12356
rect 13464 12328 14188 12356
rect 9732 12316 9738 12328
rect 9197 12291 9255 12297
rect 9197 12288 9209 12291
rect 8864 12260 9209 12288
rect 8665 12251 8723 12257
rect 9197 12257 9209 12260
rect 9243 12257 9255 12291
rect 9197 12251 9255 12257
rect 2498 12180 2504 12232
rect 2556 12180 2562 12232
rect 6730 12180 6736 12232
rect 6788 12220 6794 12232
rect 8294 12220 8300 12232
rect 6788 12192 8300 12220
rect 6788 12180 6794 12192
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 7374 12112 7380 12164
rect 7432 12152 7438 12164
rect 8202 12152 8208 12164
rect 7432 12124 8208 12152
rect 7432 12112 7438 12124
rect 8202 12112 8208 12124
rect 8260 12112 8266 12164
rect 3881 12087 3939 12093
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 4706 12084 4712 12096
rect 3927 12056 4712 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 4706 12044 4712 12056
rect 4764 12084 4770 12096
rect 5166 12084 5172 12096
rect 4764 12056 5172 12084
rect 4764 12044 4770 12056
rect 5166 12044 5172 12056
rect 5224 12044 5230 12096
rect 7650 12044 7656 12096
rect 7708 12044 7714 12096
rect 8680 12084 8708 12251
rect 10870 12248 10876 12300
rect 10928 12288 10934 12300
rect 10965 12291 11023 12297
rect 10965 12288 10977 12291
rect 10928 12260 10977 12288
rect 10928 12248 10934 12260
rect 10965 12257 10977 12260
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 8938 12180 8944 12232
rect 8996 12180 9002 12232
rect 9950 12112 9956 12164
rect 10008 12152 10014 12164
rect 10321 12155 10379 12161
rect 10321 12152 10333 12155
rect 10008 12124 10333 12152
rect 10008 12112 10014 12124
rect 10321 12121 10333 12124
rect 10367 12152 10379 12155
rect 11072 12152 11100 12328
rect 11330 12248 11336 12300
rect 11388 12288 11394 12300
rect 13464 12297 13492 12328
rect 14182 12316 14188 12328
rect 14240 12356 14246 12368
rect 14642 12356 14648 12368
rect 14240 12328 14648 12356
rect 14240 12316 14246 12328
rect 14642 12316 14648 12328
rect 14700 12316 14706 12368
rect 15010 12356 15016 12368
rect 14752 12328 15016 12356
rect 13449 12291 13507 12297
rect 13449 12288 13461 12291
rect 11388 12260 13461 12288
rect 11388 12248 11394 12260
rect 13449 12257 13461 12260
rect 13495 12257 13507 12291
rect 13449 12251 13507 12257
rect 13817 12291 13875 12297
rect 13817 12257 13829 12291
rect 13863 12257 13875 12291
rect 13817 12251 13875 12257
rect 14001 12291 14059 12297
rect 14001 12257 14013 12291
rect 14047 12288 14059 12291
rect 14274 12288 14280 12300
rect 14047 12260 14280 12288
rect 14047 12257 14059 12260
rect 14001 12251 14059 12257
rect 12526 12180 12532 12232
rect 12584 12220 12590 12232
rect 13262 12220 13268 12232
rect 12584 12192 13268 12220
rect 12584 12180 12590 12192
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 10367 12124 11100 12152
rect 10367 12121 10379 12124
rect 10321 12115 10379 12121
rect 11974 12112 11980 12164
rect 12032 12152 12038 12164
rect 12434 12152 12440 12164
rect 12032 12124 12440 12152
rect 12032 12112 12038 12124
rect 12434 12112 12440 12124
rect 12492 12152 12498 12164
rect 13832 12152 13860 12251
rect 14274 12248 14280 12260
rect 14332 12288 14338 12300
rect 14752 12288 14780 12328
rect 15010 12316 15016 12328
rect 15068 12356 15074 12368
rect 15068 12328 15424 12356
rect 15068 12316 15074 12328
rect 14332 12260 14780 12288
rect 14332 12248 14338 12260
rect 14826 12248 14832 12300
rect 14884 12248 14890 12300
rect 14918 12248 14924 12300
rect 14976 12248 14982 12300
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 15396 12297 15424 12328
rect 16776 12297 16804 12396
rect 17880 12368 17908 12396
rect 18138 12384 18144 12436
rect 18196 12424 18202 12436
rect 18322 12424 18328 12436
rect 18196 12396 18328 12424
rect 18196 12384 18202 12396
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 18414 12384 18420 12436
rect 18472 12384 18478 12436
rect 19153 12427 19211 12433
rect 19153 12393 19165 12427
rect 19199 12424 19211 12427
rect 19426 12424 19432 12436
rect 19199 12396 19432 12424
rect 19199 12393 19211 12396
rect 19153 12387 19211 12393
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 20346 12384 20352 12436
rect 20404 12424 20410 12436
rect 22738 12424 22744 12436
rect 20404 12396 22744 12424
rect 20404 12384 20410 12396
rect 22738 12384 22744 12396
rect 22796 12384 22802 12436
rect 23014 12384 23020 12436
rect 23072 12424 23078 12436
rect 23411 12427 23469 12433
rect 23411 12424 23423 12427
rect 23072 12396 23423 12424
rect 23072 12384 23078 12396
rect 23411 12393 23423 12396
rect 23457 12424 23469 12427
rect 24946 12424 24952 12436
rect 23457 12396 24952 12424
rect 23457 12393 23469 12396
rect 23411 12387 23469 12393
rect 24946 12384 24952 12396
rect 25004 12384 25010 12436
rect 25314 12384 25320 12436
rect 25372 12424 25378 12436
rect 25593 12427 25651 12433
rect 25593 12424 25605 12427
rect 25372 12396 25605 12424
rect 25372 12384 25378 12396
rect 25593 12393 25605 12396
rect 25639 12393 25651 12427
rect 25593 12387 25651 12393
rect 16850 12316 16856 12368
rect 16908 12356 16914 12368
rect 16908 12328 17264 12356
rect 16908 12316 16914 12328
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 15252 12260 15301 12288
rect 15252 12248 15258 12260
rect 15289 12257 15301 12260
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 15381 12291 15439 12297
rect 15381 12257 15393 12291
rect 15427 12257 15439 12291
rect 15381 12251 15439 12257
rect 16761 12291 16819 12297
rect 16761 12257 16773 12291
rect 16807 12257 16819 12291
rect 16761 12251 16819 12257
rect 17034 12248 17040 12300
rect 17092 12288 17098 12300
rect 17236 12297 17264 12328
rect 17586 12316 17592 12368
rect 17644 12356 17650 12368
rect 17770 12356 17776 12368
rect 17644 12328 17776 12356
rect 17644 12316 17650 12328
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 17862 12316 17868 12368
rect 17920 12356 17926 12368
rect 21542 12356 21548 12368
rect 17920 12328 21548 12356
rect 17920 12316 17926 12328
rect 17129 12291 17187 12297
rect 17129 12288 17141 12291
rect 17092 12260 17141 12288
rect 17092 12248 17098 12260
rect 17129 12257 17141 12260
rect 17175 12257 17187 12291
rect 17129 12251 17187 12257
rect 17221 12291 17279 12297
rect 17221 12257 17233 12291
rect 17267 12288 17279 12291
rect 17497 12291 17555 12297
rect 17497 12288 17509 12291
rect 17267 12260 17509 12288
rect 17267 12257 17279 12260
rect 17221 12251 17279 12257
rect 17497 12257 17509 12260
rect 17543 12257 17555 12291
rect 17497 12251 17555 12257
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12189 16911 12223
rect 17512 12220 17540 12251
rect 17678 12248 17684 12300
rect 17736 12248 17742 12300
rect 18064 12297 18092 12328
rect 18049 12291 18107 12297
rect 18049 12257 18061 12291
rect 18095 12257 18107 12291
rect 18049 12251 18107 12257
rect 18233 12291 18291 12297
rect 18233 12257 18245 12291
rect 18279 12288 18291 12291
rect 18506 12288 18512 12300
rect 18279 12260 18512 12288
rect 18279 12257 18291 12260
rect 18233 12251 18291 12257
rect 18506 12248 18512 12260
rect 18564 12248 18570 12300
rect 18966 12248 18972 12300
rect 19024 12248 19030 12300
rect 19429 12291 19487 12297
rect 19429 12257 19441 12291
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 19444 12220 19472 12251
rect 19610 12248 19616 12300
rect 19668 12248 19674 12300
rect 19996 12297 20024 12328
rect 21542 12316 21548 12328
rect 21600 12316 21606 12368
rect 23201 12359 23259 12365
rect 23201 12325 23213 12359
rect 23247 12356 23259 12359
rect 23658 12356 23664 12368
rect 23247 12328 23664 12356
rect 23247 12325 23259 12328
rect 23201 12319 23259 12325
rect 23658 12316 23664 12328
rect 23716 12316 23722 12368
rect 25038 12316 25044 12368
rect 25096 12356 25102 12368
rect 25096 12328 25544 12356
rect 25096 12316 25102 12328
rect 19981 12291 20039 12297
rect 19981 12257 19993 12291
rect 20027 12257 20039 12291
rect 19981 12251 20039 12257
rect 20165 12291 20223 12297
rect 20165 12257 20177 12291
rect 20211 12288 20223 12291
rect 20346 12288 20352 12300
rect 20211 12260 20352 12288
rect 20211 12257 20223 12260
rect 20165 12251 20223 12257
rect 20346 12248 20352 12260
rect 20404 12248 20410 12300
rect 20438 12248 20444 12300
rect 20496 12288 20502 12300
rect 21453 12291 21511 12297
rect 21453 12288 21465 12291
rect 20496 12260 21465 12288
rect 20496 12248 20502 12260
rect 21453 12257 21465 12260
rect 21499 12257 21511 12291
rect 21560 12288 21588 12316
rect 21821 12291 21879 12297
rect 21821 12288 21833 12291
rect 21560 12260 21833 12288
rect 21453 12251 21511 12257
rect 21821 12257 21833 12260
rect 21867 12257 21879 12291
rect 21821 12251 21879 12257
rect 22465 12291 22523 12297
rect 22465 12257 22477 12291
rect 22511 12288 22523 12291
rect 23750 12288 23756 12300
rect 22511 12260 23756 12288
rect 22511 12257 22523 12260
rect 22465 12251 22523 12257
rect 23750 12248 23756 12260
rect 23808 12248 23814 12300
rect 24486 12248 24492 12300
rect 24544 12288 24550 12300
rect 24866 12291 24924 12297
rect 24866 12288 24878 12291
rect 24544 12260 24878 12288
rect 24544 12248 24550 12260
rect 24866 12257 24878 12260
rect 24912 12257 24924 12291
rect 24866 12251 24924 12257
rect 25130 12248 25136 12300
rect 25188 12248 25194 12300
rect 25516 12297 25544 12328
rect 25225 12291 25283 12297
rect 25225 12257 25237 12291
rect 25271 12257 25283 12291
rect 25225 12251 25283 12257
rect 25501 12291 25559 12297
rect 25501 12257 25513 12291
rect 25547 12257 25559 12291
rect 25501 12251 25559 12257
rect 20990 12220 20996 12232
rect 17512 12192 20996 12220
rect 16853 12183 16911 12189
rect 12492 12124 13860 12152
rect 14461 12155 14519 12161
rect 12492 12112 12498 12124
rect 14461 12121 14473 12155
rect 14507 12152 14519 12155
rect 15010 12152 15016 12164
rect 14507 12124 15016 12152
rect 14507 12121 14519 12124
rect 14461 12115 14519 12121
rect 15010 12112 15016 12124
rect 15068 12112 15074 12164
rect 16316 12124 16528 12152
rect 10134 12084 10140 12096
rect 8680 12056 10140 12084
rect 10134 12044 10140 12056
rect 10192 12044 10198 12096
rect 13078 12044 13084 12096
rect 13136 12044 13142 12096
rect 13262 12044 13268 12096
rect 13320 12084 13326 12096
rect 16316 12084 16344 12124
rect 13320 12056 16344 12084
rect 13320 12044 13326 12056
rect 16390 12044 16396 12096
rect 16448 12044 16454 12096
rect 16500 12084 16528 12124
rect 16574 12112 16580 12164
rect 16632 12152 16638 12164
rect 16868 12152 16896 12183
rect 20990 12180 20996 12192
rect 21048 12220 21054 12232
rect 21545 12223 21603 12229
rect 21545 12220 21557 12223
rect 21048 12192 21557 12220
rect 21048 12180 21054 12192
rect 21545 12189 21557 12192
rect 21591 12189 21603 12223
rect 21545 12183 21603 12189
rect 21634 12180 21640 12232
rect 21692 12220 21698 12232
rect 21729 12223 21787 12229
rect 21729 12220 21741 12223
rect 21692 12192 21741 12220
rect 21692 12180 21698 12192
rect 21729 12189 21741 12192
rect 21775 12189 21787 12223
rect 21729 12183 21787 12189
rect 23290 12180 23296 12232
rect 23348 12220 23354 12232
rect 23474 12220 23480 12232
rect 23348 12192 23480 12220
rect 23348 12180 23354 12192
rect 23474 12180 23480 12192
rect 23532 12180 23538 12232
rect 25240 12220 25268 12251
rect 26878 12220 26884 12232
rect 25148 12192 26884 12220
rect 17586 12152 17592 12164
rect 16632 12124 17592 12152
rect 16632 12112 16638 12124
rect 17586 12112 17592 12124
rect 17644 12112 17650 12164
rect 17678 12112 17684 12164
rect 17736 12152 17742 12164
rect 17736 12124 24256 12152
rect 17736 12112 17742 12124
rect 20070 12084 20076 12096
rect 16500 12056 20076 12084
rect 20070 12044 20076 12056
rect 20128 12044 20134 12096
rect 20254 12044 20260 12096
rect 20312 12084 20318 12096
rect 20349 12087 20407 12093
rect 20349 12084 20361 12087
rect 20312 12056 20361 12084
rect 20312 12044 20318 12056
rect 20349 12053 20361 12056
rect 20395 12053 20407 12087
rect 20349 12047 20407 12053
rect 23106 12044 23112 12096
rect 23164 12084 23170 12096
rect 23385 12087 23443 12093
rect 23385 12084 23397 12087
rect 23164 12056 23397 12084
rect 23164 12044 23170 12056
rect 23385 12053 23397 12056
rect 23431 12053 23443 12087
rect 23385 12047 23443 12053
rect 23566 12044 23572 12096
rect 23624 12044 23630 12096
rect 23658 12044 23664 12096
rect 23716 12084 23722 12096
rect 23753 12087 23811 12093
rect 23753 12084 23765 12087
rect 23716 12056 23765 12084
rect 23716 12044 23722 12056
rect 23753 12053 23765 12056
rect 23799 12053 23811 12087
rect 24228 12084 24256 12124
rect 25148 12084 25176 12192
rect 26878 12180 26884 12192
rect 26936 12180 26942 12232
rect 24228 12056 25176 12084
rect 23753 12047 23811 12053
rect 25222 12044 25228 12096
rect 25280 12084 25286 12096
rect 25317 12087 25375 12093
rect 25317 12084 25329 12087
rect 25280 12056 25329 12084
rect 25280 12044 25286 12056
rect 25317 12053 25329 12056
rect 25363 12084 25375 12087
rect 25406 12084 25412 12096
rect 25363 12056 25412 12084
rect 25363 12053 25375 12056
rect 25317 12047 25375 12053
rect 25406 12044 25412 12056
rect 25464 12044 25470 12096
rect 552 11994 27416 12016
rect 552 11942 3756 11994
rect 3808 11942 3820 11994
rect 3872 11942 3884 11994
rect 3936 11942 3948 11994
rect 4000 11942 4012 11994
rect 4064 11942 10472 11994
rect 10524 11942 10536 11994
rect 10588 11942 10600 11994
rect 10652 11942 10664 11994
rect 10716 11942 10728 11994
rect 10780 11942 17188 11994
rect 17240 11942 17252 11994
rect 17304 11942 17316 11994
rect 17368 11942 17380 11994
rect 17432 11942 17444 11994
rect 17496 11942 23904 11994
rect 23956 11942 23968 11994
rect 24020 11942 24032 11994
rect 24084 11942 24096 11994
rect 24148 11942 24160 11994
rect 24212 11942 27416 11994
rect 552 11920 27416 11942
rect 2961 11883 3019 11889
rect 2961 11849 2973 11883
rect 3007 11880 3019 11883
rect 4246 11880 4252 11892
rect 3007 11852 4252 11880
rect 3007 11849 3019 11852
rect 2961 11843 3019 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 8018 11880 8024 11892
rect 6328 11852 8024 11880
rect 6328 11840 6334 11852
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 10318 11880 10324 11892
rect 8352 11852 10324 11880
rect 8352 11840 8358 11852
rect 10318 11840 10324 11852
rect 10376 11880 10382 11892
rect 11422 11880 11428 11892
rect 10376 11852 11428 11880
rect 10376 11840 10382 11852
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 11974 11840 11980 11892
rect 12032 11840 12038 11892
rect 12406 11852 20024 11880
rect 6288 11812 6316 11840
rect 5000 11784 6316 11812
rect 5000 11688 5028 11784
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 7926 11812 7932 11824
rect 6420 11784 7932 11812
rect 6420 11772 6426 11784
rect 7926 11772 7932 11784
rect 7984 11812 7990 11824
rect 12406 11812 12434 11852
rect 19150 11812 19156 11824
rect 7984 11784 12434 11812
rect 16960 11784 19156 11812
rect 7984 11772 7990 11784
rect 5077 11747 5135 11753
rect 5077 11713 5089 11747
rect 5123 11744 5135 11747
rect 11882 11744 11888 11756
rect 5123 11716 11888 11744
rect 5123 11713 5135 11716
rect 5077 11707 5135 11713
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 13280 11716 14320 11744
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11676 2835 11679
rect 3234 11676 3240 11688
rect 2823 11648 3240 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 3234 11636 3240 11648
rect 3292 11636 3298 11688
rect 4982 11636 4988 11688
rect 5040 11636 5046 11688
rect 5350 11636 5356 11688
rect 5408 11636 5414 11688
rect 5534 11636 5540 11688
rect 5592 11636 5598 11688
rect 6089 11679 6147 11685
rect 6089 11645 6101 11679
rect 6135 11645 6147 11679
rect 6089 11639 6147 11645
rect 5552 11608 5580 11636
rect 6104 11608 6132 11639
rect 6270 11636 6276 11688
rect 6328 11636 6334 11688
rect 6638 11636 6644 11688
rect 6696 11636 6702 11688
rect 6730 11636 6736 11688
rect 6788 11636 6794 11688
rect 7374 11636 7380 11688
rect 7432 11636 7438 11688
rect 7466 11636 7472 11688
rect 7524 11636 7530 11688
rect 7558 11636 7564 11688
rect 7616 11636 7622 11688
rect 7653 11679 7711 11685
rect 7653 11645 7665 11679
rect 7699 11645 7711 11679
rect 7653 11639 7711 11645
rect 6362 11608 6368 11620
rect 5552 11580 6040 11608
rect 6104 11580 6368 11608
rect 4614 11500 4620 11552
rect 4672 11500 4678 11552
rect 5718 11500 5724 11552
rect 5776 11500 5782 11552
rect 6012 11540 6040 11580
rect 6362 11568 6368 11580
rect 6420 11568 6426 11620
rect 6748 11608 6776 11636
rect 6472 11580 6776 11608
rect 7668 11608 7696 11639
rect 7742 11636 7748 11688
rect 7800 11676 7806 11688
rect 7837 11679 7895 11685
rect 7837 11676 7849 11679
rect 7800 11648 7849 11676
rect 7800 11636 7806 11648
rect 7837 11645 7849 11648
rect 7883 11645 7895 11679
rect 7837 11639 7895 11645
rect 8110 11636 8116 11688
rect 8168 11676 8174 11688
rect 8389 11679 8447 11685
rect 8389 11676 8401 11679
rect 8168 11648 8401 11676
rect 8168 11636 8174 11648
rect 8389 11645 8401 11648
rect 8435 11645 8447 11679
rect 8389 11639 8447 11645
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11676 9643 11679
rect 9674 11676 9680 11688
rect 9631 11648 9680 11676
rect 9631 11645 9643 11648
rect 9585 11639 9643 11645
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 9769 11679 9827 11685
rect 9769 11645 9781 11679
rect 9815 11645 9827 11679
rect 9769 11639 9827 11645
rect 8202 11608 8208 11620
rect 7668 11580 8208 11608
rect 6472 11540 6500 11580
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 9784 11608 9812 11639
rect 9858 11636 9864 11688
rect 9916 11676 9922 11688
rect 10137 11679 10195 11685
rect 10137 11676 10149 11679
rect 9916 11648 10149 11676
rect 9916 11636 9922 11648
rect 10137 11645 10149 11648
rect 10183 11645 10195 11679
rect 10137 11639 10195 11645
rect 10318 11636 10324 11688
rect 10376 11636 10382 11688
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11149 11679 11207 11685
rect 11149 11676 11161 11679
rect 11112 11648 11161 11676
rect 11112 11636 11118 11648
rect 11149 11645 11161 11648
rect 11195 11645 11207 11679
rect 11149 11639 11207 11645
rect 11330 11636 11336 11688
rect 11388 11636 11394 11688
rect 11606 11636 11612 11688
rect 11664 11676 11670 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11664 11648 11713 11676
rect 11664 11636 11670 11648
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 11793 11679 11851 11685
rect 11793 11645 11805 11679
rect 11839 11676 11851 11679
rect 13280 11676 13308 11716
rect 14292 11688 14320 11716
rect 11839 11648 13308 11676
rect 11839 11645 11851 11648
rect 11793 11639 11851 11645
rect 11348 11608 11376 11636
rect 8312 11580 11376 11608
rect 6012 11512 6500 11540
rect 7006 11500 7012 11552
rect 7064 11540 7070 11552
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 7064 11512 7205 11540
rect 7064 11500 7070 11512
rect 7193 11509 7205 11512
rect 7239 11509 7251 11543
rect 7193 11503 7251 11509
rect 8018 11500 8024 11552
rect 8076 11540 8082 11552
rect 8312 11540 8340 11580
rect 11422 11568 11428 11620
rect 11480 11608 11486 11620
rect 11808 11608 11836 11639
rect 13354 11636 13360 11688
rect 13412 11636 13418 11688
rect 14274 11636 14280 11688
rect 14332 11676 14338 11688
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 14332 11648 14473 11676
rect 14332 11636 14338 11648
rect 14461 11645 14473 11648
rect 14507 11645 14519 11679
rect 14461 11639 14519 11645
rect 14550 11636 14556 11688
rect 14608 11636 14614 11688
rect 14642 11636 14648 11688
rect 14700 11676 14706 11688
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 14700 11648 14933 11676
rect 14700 11636 14706 11648
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 15013 11679 15071 11685
rect 15013 11645 15025 11679
rect 15059 11676 15071 11679
rect 16960 11676 16988 11784
rect 19150 11772 19156 11784
rect 19208 11772 19214 11824
rect 19996 11812 20024 11852
rect 20070 11840 20076 11892
rect 20128 11880 20134 11892
rect 20128 11852 21220 11880
rect 20128 11840 20134 11852
rect 20346 11812 20352 11824
rect 19996 11784 20352 11812
rect 20346 11772 20352 11784
rect 20404 11772 20410 11824
rect 21192 11812 21220 11852
rect 21266 11840 21272 11892
rect 21324 11880 21330 11892
rect 22925 11883 22983 11889
rect 22925 11880 22937 11883
rect 21324 11852 22937 11880
rect 21324 11840 21330 11852
rect 22925 11849 22937 11852
rect 22971 11880 22983 11883
rect 23474 11880 23480 11892
rect 22971 11852 23480 11880
rect 22971 11849 22983 11852
rect 22925 11843 22983 11849
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 23750 11840 23756 11892
rect 23808 11880 23814 11892
rect 27062 11880 27068 11892
rect 23808 11852 27068 11880
rect 23808 11840 23814 11852
rect 27062 11840 27068 11852
rect 27120 11840 27126 11892
rect 21634 11812 21640 11824
rect 21192 11784 21640 11812
rect 21634 11772 21640 11784
rect 21692 11772 21698 11824
rect 17678 11744 17684 11756
rect 17052 11716 17684 11744
rect 17052 11685 17080 11716
rect 17678 11704 17684 11716
rect 17736 11704 17742 11756
rect 18782 11744 18788 11756
rect 18064 11716 18788 11744
rect 18064 11685 18092 11716
rect 18782 11704 18788 11716
rect 18840 11704 18846 11756
rect 23014 11744 23020 11756
rect 22572 11716 23020 11744
rect 15059 11648 16988 11676
rect 17037 11679 17095 11685
rect 15059 11645 15071 11648
rect 15013 11639 15071 11645
rect 17037 11645 17049 11679
rect 17083 11645 17095 11679
rect 17037 11639 17095 11645
rect 17221 11679 17279 11685
rect 17221 11645 17233 11679
rect 17267 11676 17279 11679
rect 17497 11679 17555 11685
rect 17497 11676 17509 11679
rect 17267 11648 17509 11676
rect 17267 11645 17279 11648
rect 17221 11639 17279 11645
rect 17497 11645 17509 11648
rect 17543 11645 17555 11679
rect 17497 11639 17555 11645
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 11480 11580 11836 11608
rect 13112 11611 13170 11617
rect 11480 11568 11486 11580
rect 13112 11577 13124 11611
rect 13158 11608 13170 11611
rect 13446 11608 13452 11620
rect 13158 11580 13452 11608
rect 13158 11577 13170 11580
rect 13112 11571 13170 11577
rect 13446 11568 13452 11580
rect 13504 11568 13510 11620
rect 14826 11568 14832 11620
rect 14884 11608 14890 11620
rect 15028 11608 15056 11639
rect 16393 11611 16451 11617
rect 16393 11608 16405 11611
rect 14884 11580 15056 11608
rect 15120 11580 16405 11608
rect 14884 11568 14890 11580
rect 8076 11512 8340 11540
rect 8076 11500 8082 11512
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8444 11512 9045 11540
rect 8444 11500 8450 11512
rect 9033 11509 9045 11512
rect 9079 11540 9091 11543
rect 9122 11540 9128 11552
rect 9079 11512 9128 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 9401 11543 9459 11549
rect 9401 11509 9413 11543
rect 9447 11540 9459 11543
rect 9490 11540 9496 11552
rect 9447 11512 9496 11540
rect 9447 11509 9459 11512
rect 9401 11503 9459 11509
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 10965 11543 11023 11549
rect 10965 11509 10977 11543
rect 11011 11540 11023 11543
rect 11146 11540 11152 11552
rect 11011 11512 11152 11540
rect 11011 11509 11023 11512
rect 10965 11503 11023 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 14182 11500 14188 11552
rect 14240 11540 14246 11552
rect 15120 11540 15148 11580
rect 16393 11577 16405 11580
rect 16439 11608 16451 11611
rect 16853 11611 16911 11617
rect 16853 11608 16865 11611
rect 16439 11580 16865 11608
rect 16439 11577 16451 11580
rect 16393 11571 16451 11577
rect 16853 11577 16865 11580
rect 16899 11577 16911 11611
rect 17512 11608 17540 11639
rect 18138 11636 18144 11688
rect 18196 11676 18202 11688
rect 22572 11676 22600 11716
rect 23014 11704 23020 11716
rect 23072 11704 23078 11756
rect 24210 11744 24216 11756
rect 23216 11716 24216 11744
rect 18196 11648 22600 11676
rect 18196 11636 18202 11648
rect 22646 11636 22652 11688
rect 22704 11636 22710 11688
rect 23216 11685 23244 11716
rect 24210 11704 24216 11716
rect 24268 11744 24274 11756
rect 24394 11744 24400 11756
rect 24268 11716 24400 11744
rect 24268 11704 24274 11716
rect 24394 11704 24400 11716
rect 24452 11704 24458 11756
rect 23201 11679 23259 11685
rect 23201 11645 23213 11679
rect 23247 11645 23259 11679
rect 23201 11639 23259 11645
rect 23290 11636 23296 11688
rect 23348 11676 23354 11688
rect 23385 11679 23443 11685
rect 23385 11676 23397 11679
rect 23348 11648 23397 11676
rect 23348 11636 23354 11648
rect 23385 11645 23397 11648
rect 23431 11645 23443 11679
rect 23385 11639 23443 11645
rect 24857 11679 24915 11685
rect 24857 11645 24869 11679
rect 24903 11645 24915 11679
rect 24857 11639 24915 11645
rect 24949 11679 25007 11685
rect 24949 11645 24961 11679
rect 24995 11676 25007 11679
rect 25038 11676 25044 11688
rect 24995 11648 25044 11676
rect 24995 11645 25007 11648
rect 24949 11639 25007 11645
rect 18156 11608 18184 11636
rect 17512 11580 18184 11608
rect 16853 11571 16911 11577
rect 18690 11568 18696 11620
rect 18748 11568 18754 11620
rect 18782 11568 18788 11620
rect 18840 11608 18846 11620
rect 18840 11580 22094 11608
rect 18840 11568 18846 11580
rect 14240 11512 15148 11540
rect 14240 11500 14246 11512
rect 15470 11500 15476 11552
rect 15528 11500 15534 11552
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 16942 11540 16948 11552
rect 16724 11512 16948 11540
rect 16724 11500 16730 11512
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17313 11543 17371 11549
rect 17313 11509 17325 11543
rect 17359 11540 17371 11543
rect 17678 11540 17684 11552
rect 17359 11512 17684 11540
rect 17359 11509 17371 11512
rect 17313 11503 17371 11509
rect 17678 11500 17684 11512
rect 17736 11500 17742 11552
rect 18230 11500 18236 11552
rect 18288 11500 18294 11552
rect 19978 11500 19984 11552
rect 20036 11500 20042 11552
rect 22066 11540 22094 11580
rect 22186 11568 22192 11620
rect 22244 11608 22250 11620
rect 22382 11611 22440 11617
rect 22382 11608 22394 11611
rect 22244 11580 22394 11608
rect 22244 11568 22250 11580
rect 22382 11577 22394 11580
rect 22428 11577 22440 11611
rect 23106 11608 23112 11620
rect 22382 11571 22440 11577
rect 22664 11580 23112 11608
rect 22664 11540 22692 11580
rect 23106 11568 23112 11580
rect 23164 11568 23170 11620
rect 24872 11608 24900 11639
rect 25038 11636 25044 11648
rect 25096 11636 25102 11688
rect 25216 11611 25274 11617
rect 24872 11580 24992 11608
rect 22066 11512 22692 11540
rect 22738 11500 22744 11552
rect 22796 11500 22802 11552
rect 22909 11543 22967 11549
rect 22909 11509 22921 11543
rect 22955 11540 22967 11543
rect 23201 11543 23259 11549
rect 23201 11540 23213 11543
rect 22955 11512 23213 11540
rect 22955 11509 22967 11512
rect 22909 11503 22967 11509
rect 23201 11509 23213 11512
rect 23247 11509 23259 11543
rect 23201 11503 23259 11509
rect 24213 11543 24271 11549
rect 24213 11509 24225 11543
rect 24259 11540 24271 11543
rect 24302 11540 24308 11552
rect 24259 11512 24308 11540
rect 24259 11509 24271 11512
rect 24213 11503 24271 11509
rect 24302 11500 24308 11512
rect 24360 11500 24366 11552
rect 24964 11540 24992 11580
rect 25216 11577 25228 11611
rect 25262 11608 25274 11611
rect 25314 11608 25320 11620
rect 25262 11580 25320 11608
rect 25262 11577 25274 11580
rect 25216 11571 25274 11577
rect 25314 11568 25320 11580
rect 25372 11568 25378 11620
rect 26142 11540 26148 11552
rect 24964 11512 26148 11540
rect 26142 11500 26148 11512
rect 26200 11540 26206 11552
rect 26329 11543 26387 11549
rect 26329 11540 26341 11543
rect 26200 11512 26341 11540
rect 26200 11500 26206 11512
rect 26329 11509 26341 11512
rect 26375 11509 26387 11543
rect 26329 11503 26387 11509
rect 552 11450 27576 11472
rect 552 11398 7114 11450
rect 7166 11398 7178 11450
rect 7230 11398 7242 11450
rect 7294 11398 7306 11450
rect 7358 11398 7370 11450
rect 7422 11398 13830 11450
rect 13882 11398 13894 11450
rect 13946 11398 13958 11450
rect 14010 11398 14022 11450
rect 14074 11398 14086 11450
rect 14138 11398 20546 11450
rect 20598 11398 20610 11450
rect 20662 11398 20674 11450
rect 20726 11398 20738 11450
rect 20790 11398 20802 11450
rect 20854 11398 27262 11450
rect 27314 11398 27326 11450
rect 27378 11398 27390 11450
rect 27442 11398 27454 11450
rect 27506 11398 27518 11450
rect 27570 11398 27576 11450
rect 552 11376 27576 11398
rect 1394 11296 1400 11348
rect 1452 11336 1458 11348
rect 6181 11339 6239 11345
rect 1452 11308 4844 11336
rect 1452 11296 1458 11308
rect 3142 11160 3148 11212
rect 3200 11160 3206 11212
rect 3329 11203 3387 11209
rect 3329 11169 3341 11203
rect 3375 11200 3387 11203
rect 4246 11200 4252 11212
rect 3375 11172 4252 11200
rect 3375 11169 3387 11172
rect 3329 11163 3387 11169
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 4338 11092 4344 11144
rect 4396 11132 4402 11144
rect 4433 11135 4491 11141
rect 4433 11132 4445 11135
rect 4396 11104 4445 11132
rect 4396 11092 4402 11104
rect 4433 11101 4445 11104
rect 4479 11101 4491 11135
rect 4816 11132 4844 11308
rect 6181 11305 6193 11339
rect 6227 11336 6239 11339
rect 7558 11336 7564 11348
rect 6227 11308 7564 11336
rect 6227 11305 6239 11308
rect 6181 11299 6239 11305
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 8110 11296 8116 11348
rect 8168 11296 8174 11348
rect 8202 11296 8208 11348
rect 8260 11296 8266 11348
rect 9309 11339 9367 11345
rect 9309 11336 9321 11339
rect 8864 11308 9321 11336
rect 7006 11277 7012 11280
rect 4908 11240 6960 11268
rect 4908 11209 4936 11240
rect 4893 11203 4951 11209
rect 4893 11169 4905 11203
rect 4939 11169 4951 11203
rect 4893 11163 4951 11169
rect 4982 11160 4988 11212
rect 5040 11200 5046 11212
rect 5077 11203 5135 11209
rect 5077 11200 5089 11203
rect 5040 11172 5089 11200
rect 5040 11160 5046 11172
rect 5077 11169 5089 11172
rect 5123 11169 5135 11203
rect 5077 11163 5135 11169
rect 5166 11160 5172 11212
rect 5224 11200 5230 11212
rect 5445 11203 5503 11209
rect 5445 11200 5457 11203
rect 5224 11172 5457 11200
rect 5224 11160 5230 11172
rect 5445 11169 5457 11172
rect 5491 11169 5503 11203
rect 5445 11163 5503 11169
rect 5994 11160 6000 11212
rect 6052 11160 6058 11212
rect 6733 11203 6791 11209
rect 6733 11169 6745 11203
rect 6779 11200 6791 11203
rect 6822 11200 6828 11212
rect 6779 11172 6828 11200
rect 6779 11169 6791 11172
rect 6733 11163 6791 11169
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 6932 11200 6960 11240
rect 7000 11231 7012 11277
rect 7064 11268 7070 11280
rect 7064 11240 7100 11268
rect 7006 11228 7012 11231
rect 7064 11228 7070 11240
rect 8386 11228 8392 11280
rect 8444 11228 8450 11280
rect 8864 11277 8892 11308
rect 9309 11305 9321 11308
rect 9355 11336 9367 11339
rect 9398 11336 9404 11348
rect 9355 11308 9404 11336
rect 9355 11305 9367 11308
rect 9309 11299 9367 11305
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 13538 11336 13544 11348
rect 12400 11308 13544 11336
rect 12400 11296 12406 11308
rect 13538 11296 13544 11308
rect 13596 11336 13602 11348
rect 13725 11339 13783 11345
rect 13725 11336 13737 11339
rect 13596 11308 13737 11336
rect 13596 11296 13602 11308
rect 13725 11305 13737 11308
rect 13771 11305 13783 11339
rect 13725 11299 13783 11305
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 21450 11336 21456 11348
rect 13872 11308 21456 11336
rect 13872 11296 13878 11308
rect 21450 11296 21456 11308
rect 21508 11296 21514 11348
rect 23290 11296 23296 11348
rect 23348 11336 23354 11348
rect 23677 11339 23735 11345
rect 23677 11336 23689 11339
rect 23348 11308 23689 11336
rect 23348 11296 23354 11308
rect 23677 11305 23689 11308
rect 23723 11305 23735 11339
rect 23677 11299 23735 11305
rect 24486 11296 24492 11348
rect 24544 11296 24550 11348
rect 25314 11296 25320 11348
rect 25372 11296 25378 11348
rect 8849 11271 8907 11277
rect 8849 11237 8861 11271
rect 8895 11237 8907 11271
rect 8849 11231 8907 11237
rect 9122 11228 9128 11280
rect 9180 11268 9186 11280
rect 11517 11271 11575 11277
rect 11517 11268 11529 11271
rect 9180 11240 11529 11268
rect 9180 11228 9186 11240
rect 11517 11237 11529 11240
rect 11563 11237 11575 11271
rect 11517 11231 11575 11237
rect 11882 11228 11888 11280
rect 11940 11268 11946 11280
rect 16574 11268 16580 11280
rect 11940 11240 16580 11268
rect 11940 11228 11946 11240
rect 16574 11228 16580 11240
rect 16632 11228 16638 11280
rect 19242 11228 19248 11280
rect 19300 11228 19306 11280
rect 21542 11228 21548 11280
rect 21600 11228 21606 11280
rect 23474 11228 23480 11280
rect 23532 11228 23538 11280
rect 24210 11228 24216 11280
rect 24268 11268 24274 11280
rect 24765 11271 24823 11277
rect 24765 11268 24777 11271
rect 24268 11240 24777 11268
rect 24268 11228 24274 11240
rect 24765 11237 24777 11240
rect 24811 11237 24823 11271
rect 24765 11231 24823 11237
rect 24854 11228 24860 11280
rect 24912 11268 24918 11280
rect 24912 11240 25912 11268
rect 24912 11228 24918 11240
rect 7466 11200 7472 11212
rect 6932 11172 7472 11200
rect 7466 11160 7472 11172
rect 7524 11160 7530 11212
rect 8573 11203 8631 11209
rect 8573 11169 8585 11203
rect 8619 11169 8631 11203
rect 8573 11163 8631 11169
rect 9033 11203 9091 11209
rect 9033 11169 9045 11203
rect 9079 11200 9091 11203
rect 10042 11200 10048 11212
rect 9079 11172 10048 11200
rect 9079 11169 9091 11172
rect 9033 11163 9091 11169
rect 5353 11135 5411 11141
rect 5353 11132 5365 11135
rect 4816 11104 5365 11132
rect 4433 11095 4491 11101
rect 5353 11101 5365 11104
rect 5399 11132 5411 11135
rect 5534 11132 5540 11144
rect 5399 11104 5540 11132
rect 5399 11101 5411 11104
rect 5353 11095 5411 11101
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11101 5871 11135
rect 8588 11132 8616 11163
rect 9048 11132 9076 11163
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 11054 11160 11060 11212
rect 11112 11200 11118 11212
rect 11149 11203 11207 11209
rect 11149 11200 11161 11203
rect 11112 11172 11161 11200
rect 11112 11160 11118 11172
rect 11149 11169 11161 11172
rect 11195 11169 11207 11203
rect 11149 11163 11207 11169
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 11296 11172 11341 11200
rect 11296 11160 11302 11172
rect 11422 11160 11428 11212
rect 11480 11160 11486 11212
rect 11698 11209 11704 11212
rect 11655 11203 11704 11209
rect 11655 11169 11667 11203
rect 11701 11169 11704 11203
rect 11655 11163 11704 11169
rect 11698 11160 11704 11163
rect 11756 11160 11762 11212
rect 12618 11209 12624 11212
rect 12612 11163 12624 11209
rect 12618 11160 12624 11163
rect 12676 11160 12682 11212
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11200 16267 11203
rect 16298 11200 16304 11212
rect 16255 11172 16304 11200
rect 16255 11169 16267 11172
rect 16209 11163 16267 11169
rect 16298 11160 16304 11172
rect 16356 11160 16362 11212
rect 16482 11209 16488 11212
rect 16476 11163 16488 11209
rect 16482 11160 16488 11163
rect 16540 11160 16546 11212
rect 17586 11160 17592 11212
rect 17644 11200 17650 11212
rect 18325 11203 18383 11209
rect 18325 11200 18337 11203
rect 17644 11172 18337 11200
rect 17644 11160 17650 11172
rect 18325 11169 18337 11172
rect 18371 11169 18383 11203
rect 18325 11163 18383 11169
rect 18506 11160 18512 11212
rect 18564 11160 18570 11212
rect 18874 11160 18880 11212
rect 18932 11160 18938 11212
rect 19518 11160 19524 11212
rect 19576 11160 19582 11212
rect 19610 11160 19616 11212
rect 19668 11160 19674 11212
rect 19702 11160 19708 11212
rect 19760 11160 19766 11212
rect 19886 11160 19892 11212
rect 19944 11160 19950 11212
rect 22646 11160 22652 11212
rect 22704 11200 22710 11212
rect 23293 11203 23351 11209
rect 23293 11200 23305 11203
rect 22704 11172 23305 11200
rect 22704 11160 22710 11172
rect 23293 11169 23305 11172
rect 23339 11200 23351 11203
rect 25038 11200 25044 11212
rect 23339 11172 25044 11200
rect 23339 11169 23351 11172
rect 23293 11163 23351 11169
rect 25038 11160 25044 11172
rect 25096 11160 25102 11212
rect 25130 11160 25136 11212
rect 25188 11200 25194 11212
rect 25501 11203 25559 11209
rect 25501 11200 25513 11203
rect 25188 11172 25513 11200
rect 25188 11160 25194 11172
rect 25501 11169 25513 11172
rect 25547 11200 25559 11203
rect 25682 11200 25688 11212
rect 25547 11172 25688 11200
rect 25547 11169 25559 11172
rect 25501 11163 25559 11169
rect 25682 11160 25688 11172
rect 25740 11160 25746 11212
rect 8588 11104 9076 11132
rect 5813 11095 5871 11101
rect 5074 11024 5080 11076
rect 5132 11064 5138 11076
rect 5828 11064 5856 11095
rect 9858 11092 9864 11144
rect 9916 11092 9922 11144
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 11020 11104 12357 11132
rect 11020 11092 11026 11104
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 5132 11036 5856 11064
rect 5132 11024 5138 11036
rect 9398 11024 9404 11076
rect 9456 11064 9462 11076
rect 9674 11064 9680 11076
rect 9456 11036 9680 11064
rect 9456 11024 9462 11036
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 3326 10956 3332 11008
rect 3384 10956 3390 11008
rect 8386 10956 8392 11008
rect 8444 10996 8450 11008
rect 8665 10999 8723 11005
rect 8665 10996 8677 10999
rect 8444 10968 8677 10996
rect 8444 10956 8450 10968
rect 8665 10965 8677 10968
rect 8711 10965 8723 10999
rect 8665 10959 8723 10965
rect 11793 10999 11851 11005
rect 11793 10965 11805 10999
rect 11839 10996 11851 10999
rect 12158 10996 12164 11008
rect 11839 10968 12164 10996
rect 11839 10965 11851 10968
rect 11793 10959 11851 10965
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 12360 10996 12388 11095
rect 18598 11092 18604 11144
rect 18656 11092 18662 11144
rect 18693 11135 18751 11141
rect 18693 11101 18705 11135
rect 18739 11132 18751 11135
rect 20530 11132 20536 11144
rect 18739 11104 20536 11132
rect 18739 11101 18751 11104
rect 18693 11095 18751 11101
rect 20530 11092 20536 11104
rect 20588 11092 20594 11144
rect 23566 11092 23572 11144
rect 23624 11132 23630 11144
rect 24029 11135 24087 11141
rect 24029 11132 24041 11135
rect 23624 11104 24041 11132
rect 23624 11092 23630 11104
rect 24029 11101 24041 11104
rect 24075 11101 24087 11135
rect 24029 11095 24087 11101
rect 24118 11092 24124 11144
rect 24176 11092 24182 11144
rect 24210 11092 24216 11144
rect 24268 11092 24274 11144
rect 24302 11092 24308 11144
rect 24360 11092 24366 11144
rect 25590 11132 25596 11144
rect 25056 11104 25596 11132
rect 17589 11067 17647 11073
rect 17589 11033 17601 11067
rect 17635 11064 17647 11067
rect 17954 11064 17960 11076
rect 17635 11036 17960 11064
rect 17635 11033 17647 11036
rect 17589 11027 17647 11033
rect 17954 11024 17960 11036
rect 18012 11024 18018 11076
rect 19061 11067 19119 11073
rect 19061 11033 19073 11067
rect 19107 11064 19119 11067
rect 20070 11064 20076 11076
rect 19107 11036 20076 11064
rect 19107 11033 19119 11036
rect 19061 11027 19119 11033
rect 20070 11024 20076 11036
rect 20128 11024 20134 11076
rect 23845 11067 23903 11073
rect 23845 11033 23857 11067
rect 23891 11064 23903 11067
rect 25056 11064 25084 11104
rect 25590 11092 25596 11104
rect 25648 11132 25654 11144
rect 25884 11141 25912 11240
rect 26142 11160 26148 11212
rect 26200 11160 26206 11212
rect 25777 11135 25835 11141
rect 25777 11132 25789 11135
rect 25648 11104 25789 11132
rect 25648 11092 25654 11104
rect 25777 11101 25789 11104
rect 25823 11101 25835 11135
rect 25777 11095 25835 11101
rect 25869 11135 25927 11141
rect 25869 11101 25881 11135
rect 25915 11101 25927 11135
rect 25869 11095 25927 11101
rect 23891 11036 25084 11064
rect 25133 11067 25191 11073
rect 23891 11033 23903 11036
rect 23845 11027 23903 11033
rect 25133 11033 25145 11067
rect 25179 11064 25191 11067
rect 26160 11064 26188 11160
rect 25179 11036 26188 11064
rect 25179 11033 25191 11036
rect 25133 11027 25191 11033
rect 13354 10996 13360 11008
rect 12360 10968 13360 10996
rect 13354 10956 13360 10968
rect 13412 10996 13418 11008
rect 14274 10996 14280 11008
rect 13412 10968 14280 10996
rect 13412 10956 13418 10968
rect 14274 10956 14280 10968
rect 14332 10956 14338 11008
rect 16942 10956 16948 11008
rect 17000 10996 17006 11008
rect 22554 10996 22560 11008
rect 17000 10968 22560 10996
rect 17000 10956 17006 10968
rect 22554 10956 22560 10968
rect 22612 10956 22618 11008
rect 23566 10956 23572 11008
rect 23624 10996 23630 11008
rect 23661 10999 23719 11005
rect 23661 10996 23673 10999
rect 23624 10968 23673 10996
rect 23624 10956 23630 10968
rect 23661 10965 23673 10968
rect 23707 10996 23719 10999
rect 24210 10996 24216 11008
rect 23707 10968 24216 10996
rect 23707 10965 23719 10968
rect 23661 10959 23719 10965
rect 24210 10956 24216 10968
rect 24268 10956 24274 11008
rect 25225 10999 25283 11005
rect 25225 10965 25237 10999
rect 25271 10996 25283 10999
rect 25685 10999 25743 11005
rect 25685 10996 25697 10999
rect 25271 10968 25697 10996
rect 25271 10965 25283 10968
rect 25225 10959 25283 10965
rect 25685 10965 25697 10968
rect 25731 10996 25743 10999
rect 25774 10996 25780 11008
rect 25731 10968 25780 10996
rect 25731 10965 25743 10968
rect 25685 10959 25743 10965
rect 25774 10956 25780 10968
rect 25832 10956 25838 11008
rect 25866 10956 25872 11008
rect 25924 10996 25930 11008
rect 25961 10999 26019 11005
rect 25961 10996 25973 10999
rect 25924 10968 25973 10996
rect 25924 10956 25930 10968
rect 25961 10965 25973 10968
rect 26007 10965 26019 10999
rect 25961 10959 26019 10965
rect 26050 10956 26056 11008
rect 26108 10956 26114 11008
rect 552 10906 27416 10928
rect 552 10854 3756 10906
rect 3808 10854 3820 10906
rect 3872 10854 3884 10906
rect 3936 10854 3948 10906
rect 4000 10854 4012 10906
rect 4064 10854 10472 10906
rect 10524 10854 10536 10906
rect 10588 10854 10600 10906
rect 10652 10854 10664 10906
rect 10716 10854 10728 10906
rect 10780 10854 17188 10906
rect 17240 10854 17252 10906
rect 17304 10854 17316 10906
rect 17368 10854 17380 10906
rect 17432 10854 17444 10906
rect 17496 10854 23904 10906
rect 23956 10854 23968 10906
rect 24020 10854 24032 10906
rect 24084 10854 24096 10906
rect 24148 10854 24160 10906
rect 24212 10854 27416 10906
rect 552 10832 27416 10854
rect 7742 10792 7748 10804
rect 7576 10764 7748 10792
rect 4617 10727 4675 10733
rect 4617 10693 4629 10727
rect 4663 10724 4675 10727
rect 4890 10724 4896 10736
rect 4663 10696 4896 10724
rect 4663 10693 4675 10696
rect 4617 10687 4675 10693
rect 4890 10684 4896 10696
rect 4948 10724 4954 10736
rect 4948 10696 5304 10724
rect 4948 10684 4954 10696
rect 5276 10665 5304 10696
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10656 5319 10659
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 5307 10628 5457 10656
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 5445 10625 5457 10628
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 2498 10588 2504 10600
rect 1719 10560 2504 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 2498 10548 2504 10560
rect 2556 10588 2562 10600
rect 3237 10591 3295 10597
rect 3237 10588 3249 10591
rect 2556 10560 3249 10588
rect 2556 10548 2562 10560
rect 3237 10557 3249 10560
rect 3283 10557 3295 10591
rect 3237 10551 3295 10557
rect 3326 10548 3332 10600
rect 3384 10588 3390 10600
rect 3493 10591 3551 10597
rect 3493 10588 3505 10591
rect 3384 10560 3505 10588
rect 3384 10548 3390 10560
rect 3493 10557 3505 10560
rect 3539 10557 3551 10591
rect 3493 10551 3551 10557
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10588 5687 10591
rect 5994 10588 6000 10600
rect 5675 10560 6000 10588
rect 5675 10557 5687 10560
rect 5629 10551 5687 10557
rect 5994 10548 6000 10560
rect 6052 10588 6058 10600
rect 6362 10588 6368 10600
rect 6052 10560 6368 10588
rect 6052 10548 6058 10560
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 7576 10597 7604 10764
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 9769 10795 9827 10801
rect 9769 10761 9781 10795
rect 9815 10792 9827 10795
rect 9858 10792 9864 10804
rect 9815 10764 9864 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11296 10764 12572 10792
rect 11296 10752 11302 10764
rect 7926 10684 7932 10736
rect 7984 10684 7990 10736
rect 8386 10684 8392 10736
rect 8444 10684 8450 10736
rect 12342 10724 12348 10736
rect 11404 10696 12348 10724
rect 8404 10656 8432 10684
rect 7760 10628 8432 10656
rect 7760 10597 7788 10628
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 11404 10656 11432 10696
rect 12342 10684 12348 10696
rect 12400 10684 12406 10736
rect 12544 10724 12572 10764
rect 12618 10752 12624 10804
rect 12676 10752 12682 10804
rect 15562 10792 15568 10804
rect 13096 10764 15568 10792
rect 13096 10724 13124 10764
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 16301 10795 16359 10801
rect 16301 10761 16313 10795
rect 16347 10792 16359 10795
rect 16482 10792 16488 10804
rect 16347 10764 16488 10792
rect 16347 10761 16359 10764
rect 16301 10755 16359 10761
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 18693 10795 18751 10801
rect 18693 10761 18705 10795
rect 18739 10792 18751 10795
rect 18874 10792 18880 10804
rect 18739 10764 18880 10792
rect 18739 10761 18751 10764
rect 18693 10755 18751 10761
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 19702 10752 19708 10804
rect 19760 10792 19766 10804
rect 20165 10795 20223 10801
rect 20165 10792 20177 10795
rect 19760 10764 20177 10792
rect 19760 10752 19766 10764
rect 20165 10761 20177 10764
rect 20211 10761 20223 10795
rect 20165 10755 20223 10761
rect 21266 10752 21272 10804
rect 21324 10752 21330 10804
rect 22094 10752 22100 10804
rect 22152 10752 22158 10804
rect 22186 10752 22192 10804
rect 22244 10752 22250 10804
rect 23750 10752 23756 10804
rect 23808 10792 23814 10804
rect 23937 10795 23995 10801
rect 23937 10792 23949 10795
rect 23808 10764 23949 10792
rect 23808 10752 23814 10764
rect 23937 10761 23949 10764
rect 23983 10761 23995 10795
rect 23937 10755 23995 10761
rect 12544 10696 13124 10724
rect 10192 10628 11432 10656
rect 10192 10616 10198 10628
rect 7561 10591 7619 10597
rect 7561 10557 7573 10591
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 1940 10523 1998 10529
rect 1940 10489 1952 10523
rect 1986 10520 1998 10523
rect 2406 10520 2412 10532
rect 1986 10492 2412 10520
rect 1986 10489 1998 10492
rect 1940 10483 1998 10489
rect 2406 10480 2412 10492
rect 2464 10480 2470 10532
rect 7576 10520 7604 10551
rect 7834 10548 7840 10600
rect 7892 10548 7898 10600
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10588 8079 10591
rect 8110 10588 8116 10600
rect 8067 10560 8116 10588
rect 8067 10557 8079 10560
rect 8021 10551 8079 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 8389 10591 8447 10597
rect 8389 10588 8401 10591
rect 8352 10560 8401 10588
rect 8352 10548 8358 10560
rect 8389 10557 8401 10560
rect 8435 10588 8447 10591
rect 8938 10588 8944 10600
rect 8435 10560 8944 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11404 10597 11432 10628
rect 11241 10591 11299 10597
rect 11241 10588 11253 10591
rect 11112 10560 11253 10588
rect 11112 10548 11118 10560
rect 11241 10557 11253 10560
rect 11287 10557 11299 10591
rect 11241 10551 11299 10557
rect 11389 10591 11447 10597
rect 11389 10557 11401 10591
rect 11435 10557 11447 10591
rect 11389 10551 11447 10557
rect 11698 10548 11704 10600
rect 11756 10597 11762 10600
rect 11756 10588 11764 10597
rect 11756 10560 11801 10588
rect 11756 10551 11764 10560
rect 11756 10548 11762 10551
rect 11974 10548 11980 10600
rect 12032 10548 12038 10600
rect 12158 10548 12164 10600
rect 12216 10548 12222 10600
rect 12250 10548 12256 10600
rect 12308 10548 12314 10600
rect 12360 10597 12388 10684
rect 12345 10591 12403 10597
rect 12345 10557 12357 10591
rect 12391 10557 12403 10591
rect 12345 10551 12403 10557
rect 12710 10548 12716 10600
rect 12768 10548 12774 10600
rect 13096 10597 13124 10696
rect 16574 10684 16580 10736
rect 16632 10684 16638 10736
rect 16666 10684 16672 10736
rect 16724 10684 16730 10736
rect 20070 10684 20076 10736
rect 20128 10684 20134 10736
rect 22480 10696 22876 10724
rect 16684 10656 16712 10684
rect 16500 10628 16712 10656
rect 12897 10591 12955 10597
rect 12897 10588 12909 10591
rect 12820 10560 12909 10588
rect 7926 10520 7932 10532
rect 7576 10492 7932 10520
rect 7926 10480 7932 10492
rect 7984 10480 7990 10532
rect 8205 10523 8263 10529
rect 8205 10489 8217 10523
rect 8251 10520 8263 10523
rect 8634 10523 8692 10529
rect 8634 10520 8646 10523
rect 8251 10492 8646 10520
rect 8251 10489 8263 10492
rect 8205 10483 8263 10489
rect 8634 10489 8646 10492
rect 8680 10489 8692 10523
rect 8634 10483 8692 10489
rect 11514 10480 11520 10532
rect 11572 10480 11578 10532
rect 11609 10523 11667 10529
rect 11609 10489 11621 10523
rect 11655 10489 11667 10523
rect 12820 10520 12848 10560
rect 12897 10557 12909 10560
rect 12943 10557 12955 10591
rect 12897 10551 12955 10557
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10557 13047 10591
rect 12989 10551 13047 10557
rect 13081 10591 13139 10597
rect 13081 10557 13093 10591
rect 13127 10557 13139 10591
rect 13081 10551 13139 10557
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10588 14243 10591
rect 14274 10588 14280 10600
rect 14231 10560 14280 10588
rect 14231 10557 14243 10560
rect 14185 10551 14243 10557
rect 13004 10520 13032 10551
rect 14274 10548 14280 10560
rect 14332 10548 14338 10600
rect 15654 10548 15660 10600
rect 15712 10588 15718 10600
rect 16500 10597 16528 10628
rect 17954 10616 17960 10668
rect 18012 10616 18018 10668
rect 20088 10656 20116 10684
rect 19996 10628 20116 10656
rect 20180 10628 21404 10656
rect 16485 10591 16543 10597
rect 16485 10588 16497 10591
rect 15712 10560 16497 10588
rect 15712 10548 15718 10560
rect 16485 10557 16497 10560
rect 16531 10557 16543 10591
rect 16485 10551 16543 10557
rect 16666 10548 16672 10600
rect 16724 10548 16730 10600
rect 16758 10548 16764 10600
rect 16816 10548 16822 10600
rect 16942 10548 16948 10600
rect 17000 10548 17006 10600
rect 19817 10591 19875 10597
rect 19817 10557 19829 10591
rect 19863 10588 19875 10591
rect 19996 10588 20024 10628
rect 19863 10560 20024 10588
rect 19863 10557 19875 10560
rect 19817 10551 19875 10557
rect 20070 10548 20076 10600
rect 20128 10548 20134 10600
rect 11609 10483 11667 10489
rect 12268 10492 12848 10520
rect 12912 10492 13032 10520
rect 13357 10523 13415 10529
rect 3053 10455 3111 10461
rect 3053 10421 3065 10455
rect 3099 10452 3111 10455
rect 4154 10452 4160 10464
rect 3099 10424 4160 10452
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 4706 10412 4712 10464
rect 4764 10412 4770 10464
rect 5813 10455 5871 10461
rect 5813 10421 5825 10455
rect 5859 10452 5871 10455
rect 9122 10452 9128 10464
rect 5859 10424 9128 10452
rect 5859 10421 5871 10424
rect 5813 10415 5871 10421
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 11624 10452 11652 10483
rect 9732 10424 11652 10452
rect 11885 10455 11943 10461
rect 9732 10412 9738 10424
rect 11885 10421 11897 10455
rect 11931 10452 11943 10455
rect 12268 10452 12296 10492
rect 12912 10464 12940 10492
rect 13357 10489 13369 10523
rect 13403 10520 13415 10523
rect 14430 10523 14488 10529
rect 14430 10520 14442 10523
rect 13403 10492 14442 10520
rect 13403 10489 13415 10492
rect 13357 10483 13415 10489
rect 14430 10489 14442 10492
rect 14476 10489 14488 10523
rect 14430 10483 14488 10489
rect 18138 10480 18144 10532
rect 18196 10520 18202 10532
rect 18322 10520 18328 10532
rect 18196 10492 18328 10520
rect 18196 10480 18202 10492
rect 18322 10480 18328 10492
rect 18380 10520 18386 10532
rect 20180 10520 20208 10628
rect 20346 10588 20352 10600
rect 18380 10492 20208 10520
rect 20272 10560 20352 10588
rect 18380 10480 18386 10492
rect 11931 10424 12296 10452
rect 11931 10421 11943 10424
rect 11885 10415 11943 10421
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12894 10452 12900 10464
rect 12492 10424 12900 10452
rect 12492 10412 12498 10424
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 17405 10455 17463 10461
rect 17405 10452 17417 10455
rect 17276 10424 17417 10452
rect 17276 10412 17282 10424
rect 17405 10421 17417 10424
rect 17451 10421 17463 10455
rect 17405 10415 17463 10421
rect 18046 10412 18052 10464
rect 18104 10452 18110 10464
rect 20272 10452 20300 10560
rect 20346 10548 20352 10560
rect 20404 10548 20410 10600
rect 20530 10548 20536 10600
rect 20588 10548 20594 10600
rect 21082 10548 21088 10600
rect 21140 10548 21146 10600
rect 21269 10591 21327 10597
rect 21269 10557 21281 10591
rect 21315 10557 21327 10591
rect 21376 10588 21404 10628
rect 21450 10616 21456 10668
rect 21508 10616 21514 10668
rect 22480 10665 22508 10696
rect 22465 10659 22523 10665
rect 22465 10625 22477 10659
rect 22511 10625 22523 10659
rect 22465 10619 22523 10625
rect 22554 10616 22560 10668
rect 22612 10616 22618 10668
rect 22848 10656 22876 10696
rect 22922 10684 22928 10736
rect 22980 10684 22986 10736
rect 23492 10696 23980 10724
rect 22848 10628 23336 10656
rect 21729 10591 21787 10597
rect 21729 10588 21741 10591
rect 21376 10560 21741 10588
rect 21269 10551 21327 10557
rect 21729 10557 21741 10560
rect 21775 10557 21787 10591
rect 21729 10551 21787 10557
rect 21284 10520 21312 10551
rect 22370 10548 22376 10600
rect 22428 10548 22434 10600
rect 22649 10591 22707 10597
rect 22649 10557 22661 10591
rect 22695 10590 22707 10591
rect 22738 10590 22744 10600
rect 22695 10562 22744 10590
rect 22695 10557 22707 10562
rect 22649 10551 22707 10557
rect 22738 10548 22744 10562
rect 22796 10548 22802 10600
rect 21450 10520 21456 10532
rect 21284 10492 21456 10520
rect 21450 10480 21456 10492
rect 21508 10480 21514 10532
rect 23308 10529 23336 10628
rect 23492 10597 23520 10696
rect 23952 10656 23980 10696
rect 24118 10684 24124 10736
rect 24176 10684 24182 10736
rect 25774 10684 25780 10736
rect 25832 10684 25838 10736
rect 23952 10628 24808 10656
rect 23477 10591 23535 10597
rect 23477 10557 23489 10591
rect 23523 10557 23535 10591
rect 23477 10551 23535 10557
rect 23671 10591 23729 10597
rect 23671 10557 23683 10591
rect 23717 10557 23729 10591
rect 23671 10551 23729 10557
rect 23845 10591 23903 10597
rect 23845 10557 23857 10591
rect 23891 10588 23903 10591
rect 23952 10588 23980 10628
rect 24780 10600 24808 10628
rect 23891 10560 23980 10588
rect 23891 10557 23903 10560
rect 23845 10551 23903 10557
rect 23293 10523 23351 10529
rect 22664 10492 22952 10520
rect 18104 10424 20300 10452
rect 18104 10412 18110 10424
rect 20898 10412 20904 10464
rect 20956 10412 20962 10464
rect 21266 10412 21272 10464
rect 21324 10452 21330 10464
rect 21637 10455 21695 10461
rect 21637 10452 21649 10455
rect 21324 10424 21649 10452
rect 21324 10412 21330 10424
rect 21637 10421 21649 10424
rect 21683 10421 21695 10455
rect 21637 10415 21695 10421
rect 21818 10412 21824 10464
rect 21876 10452 21882 10464
rect 22664 10452 22692 10492
rect 21876 10424 22692 10452
rect 21876 10412 21882 10424
rect 22830 10412 22836 10464
rect 22888 10412 22894 10464
rect 22924 10452 22952 10492
rect 23293 10489 23305 10523
rect 23339 10520 23351 10523
rect 23566 10520 23572 10532
rect 23339 10492 23572 10520
rect 23339 10489 23351 10492
rect 23293 10483 23351 10489
rect 23566 10480 23572 10492
rect 23624 10480 23630 10532
rect 23692 10520 23720 10551
rect 24026 10548 24032 10600
rect 24084 10548 24090 10600
rect 24670 10588 24676 10600
rect 24136 10560 24676 10588
rect 24136 10520 24164 10560
rect 24670 10548 24676 10560
rect 24728 10548 24734 10600
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 25590 10548 25596 10600
rect 25648 10548 25654 10600
rect 25866 10548 25872 10600
rect 25924 10548 25930 10600
rect 23692 10492 24164 10520
rect 24305 10523 24363 10529
rect 24305 10489 24317 10523
rect 24351 10520 24363 10523
rect 24489 10523 24547 10529
rect 24489 10520 24501 10523
rect 24351 10492 24501 10520
rect 24351 10489 24363 10492
rect 24305 10483 24363 10489
rect 24489 10489 24501 10492
rect 24535 10489 24547 10523
rect 24489 10483 24547 10489
rect 23477 10455 23535 10461
rect 23477 10452 23489 10455
rect 22924 10424 23489 10452
rect 23477 10421 23489 10424
rect 23523 10421 23535 10455
rect 23477 10415 23535 10421
rect 25409 10455 25467 10461
rect 25409 10421 25421 10455
rect 25455 10452 25467 10455
rect 25774 10452 25780 10464
rect 25455 10424 25780 10452
rect 25455 10421 25467 10424
rect 25409 10415 25467 10421
rect 25774 10412 25780 10424
rect 25832 10412 25838 10464
rect 552 10362 27576 10384
rect 552 10310 7114 10362
rect 7166 10310 7178 10362
rect 7230 10310 7242 10362
rect 7294 10310 7306 10362
rect 7358 10310 7370 10362
rect 7422 10310 13830 10362
rect 13882 10310 13894 10362
rect 13946 10310 13958 10362
rect 14010 10310 14022 10362
rect 14074 10310 14086 10362
rect 14138 10310 20546 10362
rect 20598 10310 20610 10362
rect 20662 10310 20674 10362
rect 20726 10310 20738 10362
rect 20790 10310 20802 10362
rect 20854 10310 27262 10362
rect 27314 10310 27326 10362
rect 27378 10310 27390 10362
rect 27442 10310 27454 10362
rect 27506 10310 27518 10362
rect 27570 10310 27576 10362
rect 552 10288 27576 10310
rect 2406 10208 2412 10260
rect 2464 10248 2470 10260
rect 2501 10251 2559 10257
rect 2501 10248 2513 10251
rect 2464 10220 2513 10248
rect 2464 10208 2470 10220
rect 2501 10217 2513 10220
rect 2547 10217 2559 10251
rect 2501 10211 2559 10217
rect 4154 10208 4160 10260
rect 4212 10208 4218 10260
rect 4246 10208 4252 10260
rect 4304 10208 4310 10260
rect 6181 10251 6239 10257
rect 6181 10217 6193 10251
rect 6227 10248 6239 10251
rect 7834 10248 7840 10260
rect 6227 10220 7840 10248
rect 6227 10217 6239 10220
rect 6181 10211 6239 10217
rect 7834 10208 7840 10220
rect 7892 10208 7898 10260
rect 9122 10208 9128 10260
rect 9180 10248 9186 10260
rect 16666 10248 16672 10260
rect 9180 10220 16672 10248
rect 9180 10208 9186 10220
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 16758 10208 16764 10260
rect 16816 10248 16822 10260
rect 17037 10251 17095 10257
rect 17037 10248 17049 10251
rect 16816 10220 17049 10248
rect 16816 10208 16822 10220
rect 17037 10217 17049 10220
rect 17083 10217 17095 10251
rect 17037 10211 17095 10217
rect 17954 10208 17960 10260
rect 18012 10208 18018 10260
rect 18506 10208 18512 10260
rect 18564 10208 18570 10260
rect 18690 10208 18696 10260
rect 18748 10248 18754 10260
rect 18748 10220 19656 10248
rect 18748 10208 18754 10220
rect 3602 10180 3608 10192
rect 2240 10152 3608 10180
rect 2038 10072 2044 10124
rect 2096 10072 2102 10124
rect 2240 10121 2268 10152
rect 3602 10140 3608 10152
rect 3660 10140 3666 10192
rect 4172 10180 4200 10208
rect 9585 10183 9643 10189
rect 3712 10152 5120 10180
rect 2225 10115 2283 10121
rect 2225 10081 2237 10115
rect 2271 10081 2283 10115
rect 2225 10075 2283 10081
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 2866 10112 2872 10124
rect 2731 10084 2872 10112
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 3712 10121 3740 10152
rect 5092 10124 5120 10152
rect 9585 10149 9597 10183
rect 9631 10180 9643 10183
rect 9861 10183 9919 10189
rect 9861 10180 9873 10183
rect 9631 10152 9873 10180
rect 9631 10149 9643 10152
rect 9585 10143 9643 10149
rect 9861 10149 9873 10152
rect 9907 10180 9919 10183
rect 11425 10183 11483 10189
rect 11425 10180 11437 10183
rect 9907 10152 11437 10180
rect 9907 10149 9919 10152
rect 9861 10143 9919 10149
rect 11425 10149 11437 10152
rect 11471 10149 11483 10183
rect 12434 10180 12440 10192
rect 11425 10143 11483 10149
rect 12084 10152 12440 10180
rect 3697 10115 3755 10121
rect 3697 10081 3709 10115
rect 3743 10081 3755 10115
rect 3697 10075 3755 10081
rect 3973 10115 4031 10121
rect 3973 10081 3985 10115
rect 4019 10081 4031 10115
rect 3973 10075 4031 10081
rect 4157 10115 4215 10121
rect 4157 10081 4169 10115
rect 4203 10112 4215 10115
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 4203 10084 4537 10112
rect 4203 10081 4215 10084
rect 4157 10075 4215 10081
rect 4525 10081 4537 10084
rect 4571 10112 4583 10115
rect 4706 10112 4712 10124
rect 4571 10084 4712 10112
rect 4571 10081 4583 10084
rect 4525 10075 4583 10081
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10044 3019 10047
rect 3053 10047 3111 10053
rect 3053 10044 3065 10047
rect 3007 10016 3065 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 3053 10013 3065 10016
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 2869 9979 2927 9985
rect 2869 9945 2881 9979
rect 2915 9976 2927 9979
rect 3142 9976 3148 9988
rect 2915 9948 3148 9976
rect 2915 9945 2927 9948
rect 2869 9939 2927 9945
rect 3142 9936 3148 9948
rect 3200 9976 3206 9988
rect 3789 9979 3847 9985
rect 3789 9976 3801 9979
rect 3200 9948 3801 9976
rect 3200 9936 3206 9948
rect 3789 9945 3801 9948
rect 3835 9945 3847 9979
rect 3988 9976 4016 10075
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 4890 10072 4896 10124
rect 4948 10072 4954 10124
rect 5074 10072 5080 10124
rect 5132 10072 5138 10124
rect 5166 10072 5172 10124
rect 5224 10112 5230 10124
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 5224 10084 5457 10112
rect 5224 10072 5230 10084
rect 5445 10081 5457 10084
rect 5491 10081 5503 10115
rect 5445 10075 5503 10081
rect 5902 10072 5908 10124
rect 5960 10072 5966 10124
rect 5997 10115 6055 10121
rect 5997 10081 6009 10115
rect 6043 10112 6055 10115
rect 6362 10112 6368 10124
rect 6043 10084 6368 10112
rect 6043 10081 6055 10084
rect 5997 10075 6055 10081
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7377 10115 7435 10121
rect 7377 10112 7389 10115
rect 6972 10084 7389 10112
rect 6972 10072 6978 10084
rect 7377 10081 7389 10084
rect 7423 10081 7435 10115
rect 7377 10075 7435 10081
rect 7644 10115 7702 10121
rect 7644 10081 7656 10115
rect 7690 10112 7702 10115
rect 8202 10112 8208 10124
rect 7690 10084 8208 10112
rect 7690 10081 7702 10084
rect 7644 10075 7702 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 10042 10072 10048 10124
rect 10100 10072 10106 10124
rect 11054 10072 11060 10124
rect 11112 10072 11118 10124
rect 11238 10121 11244 10124
rect 11205 10115 11244 10121
rect 11205 10081 11217 10115
rect 11205 10075 11244 10081
rect 11238 10072 11244 10075
rect 11296 10072 11302 10124
rect 11330 10072 11336 10124
rect 11388 10072 11394 10124
rect 11522 10115 11580 10121
rect 11522 10081 11534 10115
rect 11568 10112 11580 10115
rect 11698 10112 11704 10124
rect 11568 10084 11704 10112
rect 11568 10081 11580 10084
rect 11522 10075 11580 10081
rect 4246 10004 4252 10056
rect 4304 10004 4310 10056
rect 4430 10004 4436 10056
rect 4488 10004 4494 10056
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 11072 10044 11100 10072
rect 11422 10044 11428 10056
rect 11072 10016 11428 10044
rect 8941 10007 8999 10013
rect 4448 9976 4476 10004
rect 5261 9979 5319 9985
rect 5261 9976 5273 9979
rect 3988 9948 5273 9976
rect 3789 9939 3847 9945
rect 4264 9920 4292 9948
rect 5261 9945 5273 9948
rect 5307 9945 5319 9979
rect 5261 9939 5319 9945
rect 8757 9979 8815 9985
rect 8757 9945 8769 9979
rect 8803 9976 8815 9979
rect 8956 9976 8984 10007
rect 11422 10004 11428 10016
rect 11480 10004 11486 10056
rect 8803 9948 8984 9976
rect 8803 9945 8815 9948
rect 8757 9939 8815 9945
rect 2222 9868 2228 9920
rect 2280 9868 2286 9920
rect 4246 9868 4252 9920
rect 4304 9868 4310 9920
rect 4709 9911 4767 9917
rect 4709 9877 4721 9911
rect 4755 9908 4767 9911
rect 5074 9908 5080 9920
rect 4755 9880 5080 9908
rect 4755 9877 4767 9880
rect 4709 9871 4767 9877
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 9677 9911 9735 9917
rect 9677 9908 9689 9911
rect 8444 9880 9689 9908
rect 8444 9868 8450 9880
rect 9677 9877 9689 9880
rect 9723 9877 9735 9911
rect 11624 9908 11652 10084
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10112 11851 10115
rect 11882 10112 11888 10124
rect 11839 10084 11888 10112
rect 11839 10081 11851 10084
rect 11793 10075 11851 10081
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 12084 10121 12112 10152
rect 12434 10140 12440 10152
rect 12492 10140 12498 10192
rect 14274 10180 14280 10192
rect 12544 10152 14280 10180
rect 12544 10121 12572 10152
rect 14274 10140 14280 10152
rect 14332 10140 14338 10192
rect 17218 10140 17224 10192
rect 17276 10140 17282 10192
rect 17405 10183 17463 10189
rect 17405 10149 17417 10183
rect 17451 10180 17463 10183
rect 17678 10180 17684 10192
rect 17451 10152 17684 10180
rect 17451 10149 17463 10152
rect 17405 10143 17463 10149
rect 17678 10140 17684 10152
rect 17736 10140 17742 10192
rect 17972 10180 18000 10208
rect 19242 10189 19248 10192
rect 18233 10183 18291 10189
rect 18233 10180 18245 10183
rect 17972 10152 18245 10180
rect 18233 10149 18245 10152
rect 18279 10149 18291 10183
rect 19236 10180 19248 10189
rect 19203 10152 19248 10180
rect 18233 10143 18291 10149
rect 19236 10143 19248 10152
rect 19242 10140 19248 10143
rect 19300 10140 19306 10192
rect 19628 10180 19656 10220
rect 19702 10208 19708 10260
rect 19760 10248 19766 10260
rect 22738 10248 22744 10260
rect 19760 10220 22744 10248
rect 19760 10208 19766 10220
rect 22738 10208 22744 10220
rect 22796 10208 22802 10260
rect 23290 10208 23296 10260
rect 23348 10208 23354 10260
rect 24670 10208 24676 10260
rect 24728 10248 24734 10260
rect 25225 10251 25283 10257
rect 25225 10248 25237 10251
rect 24728 10220 25237 10248
rect 24728 10208 24734 10220
rect 25225 10217 25237 10220
rect 25271 10248 25283 10251
rect 26050 10248 26056 10260
rect 25271 10220 26056 10248
rect 25271 10217 25283 10220
rect 25225 10211 25283 10217
rect 26050 10208 26056 10220
rect 26108 10208 26114 10260
rect 20898 10180 20904 10192
rect 19628 10152 20904 10180
rect 20898 10140 20904 10152
rect 20956 10140 20962 10192
rect 22646 10180 22652 10192
rect 21284 10152 22652 10180
rect 11977 10115 12035 10121
rect 11977 10081 11989 10115
rect 12023 10081 12035 10115
rect 11977 10075 12035 10081
rect 12069 10115 12127 10121
rect 12069 10081 12081 10115
rect 12115 10081 12127 10115
rect 12069 10075 12127 10081
rect 12161 10115 12219 10121
rect 12161 10081 12173 10115
rect 12207 10112 12219 10115
rect 12529 10115 12587 10121
rect 12207 10084 12388 10112
rect 12207 10081 12219 10084
rect 12161 10075 12219 10081
rect 11992 10044 12020 10075
rect 11716 10016 12020 10044
rect 11716 9985 11744 10016
rect 11701 9979 11759 9985
rect 11701 9945 11713 9979
rect 11747 9945 11759 9979
rect 11701 9939 11759 9945
rect 11790 9936 11796 9988
rect 11848 9976 11854 9988
rect 12360 9976 12388 10084
rect 12529 10081 12541 10115
rect 12575 10081 12587 10115
rect 12785 10115 12843 10121
rect 12785 10112 12797 10115
rect 12529 10075 12587 10081
rect 12636 10084 12797 10112
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10044 12495 10047
rect 12636 10044 12664 10084
rect 12785 10081 12797 10084
rect 12831 10081 12843 10115
rect 12785 10075 12843 10081
rect 14366 10072 14372 10124
rect 14424 10112 14430 10124
rect 17957 10115 18015 10121
rect 17957 10112 17969 10115
rect 14424 10084 17969 10112
rect 14424 10072 14430 10084
rect 17957 10081 17969 10084
rect 18003 10112 18015 10115
rect 18046 10112 18052 10124
rect 18003 10084 18052 10112
rect 18003 10081 18015 10084
rect 17957 10075 18015 10081
rect 18046 10072 18052 10084
rect 18104 10072 18110 10124
rect 18141 10115 18199 10121
rect 18141 10081 18153 10115
rect 18187 10081 18199 10115
rect 18141 10075 18199 10081
rect 18371 10115 18429 10121
rect 18371 10081 18383 10115
rect 18417 10112 18429 10115
rect 19702 10112 19708 10124
rect 18417 10084 19708 10112
rect 18417 10081 18429 10084
rect 18371 10075 18429 10081
rect 12483 10016 12664 10044
rect 18156 10044 18184 10075
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 21284 10121 21312 10152
rect 22646 10140 22652 10152
rect 22704 10140 22710 10192
rect 23308 10180 23336 10208
rect 23032 10152 23336 10180
rect 23032 10124 23060 10152
rect 23474 10140 23480 10192
rect 23532 10140 23538 10192
rect 23661 10183 23719 10189
rect 23661 10149 23673 10183
rect 23707 10180 23719 10183
rect 24302 10180 24308 10192
rect 23707 10152 24308 10180
rect 23707 10149 23719 10152
rect 23661 10143 23719 10149
rect 24302 10140 24308 10152
rect 24360 10180 24366 10192
rect 24397 10183 24455 10189
rect 24397 10180 24409 10183
rect 24360 10152 24409 10180
rect 24360 10140 24366 10152
rect 24397 10149 24409 10152
rect 24443 10180 24455 10183
rect 25498 10180 25504 10192
rect 24443 10152 25504 10180
rect 24443 10149 24455 10152
rect 24397 10143 24455 10149
rect 21542 10121 21548 10124
rect 21269 10115 21327 10121
rect 21269 10081 21281 10115
rect 21315 10081 21327 10115
rect 21269 10075 21327 10081
rect 21536 10075 21548 10121
rect 21542 10072 21548 10075
rect 21600 10072 21606 10124
rect 23014 10072 23020 10124
rect 23072 10072 23078 10124
rect 24872 10121 24900 10152
rect 25498 10140 25504 10152
rect 25556 10140 25562 10192
rect 23293 10115 23351 10121
rect 23293 10081 23305 10115
rect 23339 10081 23351 10115
rect 23293 10075 23351 10081
rect 24581 10115 24639 10121
rect 24581 10081 24593 10115
rect 24627 10081 24639 10115
rect 24581 10075 24639 10081
rect 24857 10115 24915 10121
rect 24857 10081 24869 10115
rect 24903 10081 24915 10115
rect 24857 10075 24915 10081
rect 25041 10115 25099 10121
rect 25041 10081 25053 10115
rect 25087 10081 25099 10115
rect 25041 10075 25099 10081
rect 25133 10115 25191 10121
rect 25133 10081 25145 10115
rect 25179 10112 25191 10115
rect 25222 10112 25228 10124
rect 25179 10084 25228 10112
rect 25179 10081 25191 10084
rect 25133 10075 25191 10081
rect 18690 10044 18696 10056
rect 18156 10016 18696 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 18969 10047 19027 10053
rect 18969 10013 18981 10047
rect 19015 10013 19027 10047
rect 18969 10007 19027 10013
rect 11848 9948 12388 9976
rect 11848 9936 11854 9948
rect 12250 9908 12256 9920
rect 11624 9880 12256 9908
rect 9677 9871 9735 9877
rect 12250 9868 12256 9880
rect 12308 9868 12314 9920
rect 12360 9908 12388 9948
rect 13909 9979 13967 9985
rect 13909 9945 13921 9979
rect 13955 9976 13967 9979
rect 14458 9976 14464 9988
rect 13955 9948 14464 9976
rect 13955 9945 13967 9948
rect 13909 9939 13967 9945
rect 13924 9908 13952 9939
rect 14458 9936 14464 9948
rect 14516 9936 14522 9988
rect 12360 9880 13952 9908
rect 18984 9908 19012 10007
rect 22554 10004 22560 10056
rect 22612 10044 22618 10056
rect 22922 10044 22928 10056
rect 22612 10016 22928 10044
rect 22612 10004 22618 10016
rect 22922 10004 22928 10016
rect 22980 10044 22986 10056
rect 23201 10047 23259 10053
rect 23201 10044 23213 10047
rect 22980 10016 23213 10044
rect 22980 10004 22986 10016
rect 23201 10013 23213 10016
rect 23247 10044 23259 10047
rect 23308 10044 23336 10075
rect 23247 10016 23336 10044
rect 24596 10044 24624 10075
rect 25056 10044 25084 10075
rect 25222 10072 25228 10084
rect 25280 10072 25286 10124
rect 25314 10072 25320 10124
rect 25372 10072 25378 10124
rect 24596 10016 25084 10044
rect 23247 10013 23259 10016
rect 23201 10007 23259 10013
rect 20346 9936 20352 9988
rect 20404 9936 20410 9988
rect 23658 9976 23664 9988
rect 22199 9948 23664 9976
rect 19334 9908 19340 9920
rect 18984 9880 19340 9908
rect 19334 9868 19340 9880
rect 19392 9908 19398 9920
rect 20070 9908 20076 9920
rect 19392 9880 20076 9908
rect 19392 9868 19398 9880
rect 20070 9868 20076 9880
rect 20128 9868 20134 9920
rect 21082 9868 21088 9920
rect 21140 9908 21146 9920
rect 22199 9908 22227 9948
rect 23658 9936 23664 9948
rect 23716 9976 23722 9988
rect 24596 9976 24624 10016
rect 23716 9948 24624 9976
rect 23716 9936 23722 9948
rect 21140 9880 22227 9908
rect 21140 9868 21146 9880
rect 22554 9868 22560 9920
rect 22612 9908 22618 9920
rect 22649 9911 22707 9917
rect 22649 9908 22661 9911
rect 22612 9880 22661 9908
rect 22612 9868 22618 9880
rect 22649 9877 22661 9880
rect 22695 9877 22707 9911
rect 22649 9871 22707 9877
rect 22738 9868 22744 9920
rect 22796 9908 22802 9920
rect 22833 9911 22891 9917
rect 22833 9908 22845 9911
rect 22796 9880 22845 9908
rect 22796 9868 22802 9880
rect 22833 9877 22845 9880
rect 22879 9908 22891 9911
rect 22922 9908 22928 9920
rect 22879 9880 22928 9908
rect 22879 9877 22891 9880
rect 22833 9871 22891 9877
rect 22922 9868 22928 9880
rect 22980 9868 22986 9920
rect 24026 9868 24032 9920
rect 24084 9908 24090 9920
rect 24762 9908 24768 9920
rect 24084 9880 24768 9908
rect 24084 9868 24090 9880
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 24854 9868 24860 9920
rect 24912 9868 24918 9920
rect 552 9818 27416 9840
rect 552 9766 3756 9818
rect 3808 9766 3820 9818
rect 3872 9766 3884 9818
rect 3936 9766 3948 9818
rect 4000 9766 4012 9818
rect 4064 9766 10472 9818
rect 10524 9766 10536 9818
rect 10588 9766 10600 9818
rect 10652 9766 10664 9818
rect 10716 9766 10728 9818
rect 10780 9766 17188 9818
rect 17240 9766 17252 9818
rect 17304 9766 17316 9818
rect 17368 9766 17380 9818
rect 17432 9766 17444 9818
rect 17496 9766 23904 9818
rect 23956 9766 23968 9818
rect 24020 9766 24032 9818
rect 24084 9766 24096 9818
rect 24148 9766 24160 9818
rect 24212 9766 27416 9818
rect 552 9744 27416 9766
rect 1857 9707 1915 9713
rect 1857 9673 1869 9707
rect 1903 9704 1915 9707
rect 2038 9704 2044 9716
rect 1903 9676 2044 9704
rect 1903 9673 1915 9676
rect 1857 9667 1915 9673
rect 2038 9664 2044 9676
rect 2096 9664 2102 9716
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 3053 9707 3111 9713
rect 3053 9704 3065 9707
rect 2924 9676 3065 9704
rect 2924 9664 2930 9676
rect 3053 9673 3065 9676
rect 3099 9673 3111 9707
rect 3053 9667 3111 9673
rect 4154 9664 4160 9716
rect 4212 9704 4218 9716
rect 4798 9704 4804 9716
rect 4212 9676 4804 9704
rect 4212 9664 4218 9676
rect 4798 9664 4804 9676
rect 4856 9664 4862 9716
rect 8202 9664 8208 9716
rect 8260 9664 8266 9716
rect 16574 9704 16580 9716
rect 16316 9676 16580 9704
rect 2130 9596 2136 9648
rect 2188 9636 2194 9648
rect 3237 9639 3295 9645
rect 3237 9636 3249 9639
rect 2188 9608 3249 9636
rect 2188 9596 2194 9608
rect 3237 9605 3249 9608
rect 3283 9605 3295 9639
rect 3237 9599 3295 9605
rect 3602 9596 3608 9648
rect 3660 9636 3666 9648
rect 3973 9639 4031 9645
rect 3973 9636 3985 9639
rect 3660 9608 3985 9636
rect 3660 9596 3666 9608
rect 3973 9605 3985 9608
rect 4019 9605 4031 9639
rect 5074 9636 5080 9648
rect 3973 9599 4031 9605
rect 4172 9608 5080 9636
rect 1946 9528 1952 9580
rect 2004 9528 2010 9580
rect 2222 9528 2228 9580
rect 2280 9568 2286 9580
rect 4172 9577 4200 9608
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 7193 9639 7251 9645
rect 7193 9605 7205 9639
rect 7239 9636 7251 9639
rect 7742 9636 7748 9648
rect 7239 9608 7748 9636
rect 7239 9605 7251 9608
rect 7193 9599 7251 9605
rect 7742 9596 7748 9608
rect 7800 9596 7806 9648
rect 8110 9636 8116 9648
rect 7852 9608 8116 9636
rect 2501 9571 2559 9577
rect 2501 9568 2513 9571
rect 2280 9540 2513 9568
rect 2280 9528 2286 9540
rect 2501 9537 2513 9540
rect 2547 9537 2559 9571
rect 4157 9571 4215 9577
rect 4157 9568 4169 9571
rect 2501 9531 2559 9537
rect 2792 9540 4169 9568
rect 2792 9509 2820 9540
rect 4157 9537 4169 9540
rect 4203 9537 4215 9571
rect 5261 9571 5319 9577
rect 5261 9568 5273 9571
rect 4157 9531 4215 9537
rect 4816 9540 5273 9568
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9500 1639 9503
rect 2777 9503 2835 9509
rect 2777 9500 2789 9503
rect 1627 9472 2789 9500
rect 1627 9469 1639 9472
rect 1581 9463 1639 9469
rect 2777 9469 2789 9472
rect 2823 9469 2835 9503
rect 2777 9463 2835 9469
rect 2866 9460 2872 9512
rect 2924 9500 2930 9512
rect 2924 9472 3740 9500
rect 2924 9460 2930 9472
rect 1857 9435 1915 9441
rect 1857 9401 1869 9435
rect 1903 9432 1915 9435
rect 2130 9432 2136 9444
rect 1903 9404 2136 9432
rect 1903 9401 1915 9404
rect 1857 9395 1915 9401
rect 2130 9392 2136 9404
rect 2188 9392 2194 9444
rect 3050 9392 3056 9444
rect 3108 9392 3114 9444
rect 1673 9367 1731 9373
rect 1673 9333 1685 9367
rect 1719 9364 1731 9367
rect 2590 9364 2596 9376
rect 1719 9336 2596 9364
rect 1719 9333 1731 9336
rect 1673 9327 1731 9333
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 3712 9364 3740 9472
rect 3786 9460 3792 9512
rect 3844 9460 3850 9512
rect 4246 9460 4252 9512
rect 4304 9460 4310 9512
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9469 4399 9503
rect 4341 9463 4399 9469
rect 3804 9432 3832 9460
rect 4356 9432 4384 9463
rect 4430 9460 4436 9512
rect 4488 9460 4494 9512
rect 4816 9432 4844 9540
rect 5261 9537 5273 9540
rect 5307 9568 5319 9571
rect 5902 9568 5908 9580
rect 5307 9540 5908 9568
rect 5307 9537 5319 9540
rect 5261 9531 5319 9537
rect 5902 9528 5908 9540
rect 5960 9528 5966 9580
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9568 6607 9571
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 6595 9540 7113 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7852 9568 7880 9608
rect 8110 9596 8116 9608
rect 8168 9636 8174 9648
rect 8570 9636 8576 9648
rect 8168 9608 8576 9636
rect 8168 9596 8174 9608
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 8665 9639 8723 9645
rect 8665 9605 8677 9639
rect 8711 9636 8723 9639
rect 9766 9636 9772 9648
rect 8711 9608 9772 9636
rect 8711 9605 8723 9608
rect 8665 9599 8723 9605
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 13538 9636 13544 9648
rect 12768 9608 13544 9636
rect 12768 9596 12774 9608
rect 13538 9596 13544 9608
rect 13596 9596 13602 9648
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 15841 9639 15899 9645
rect 15841 9636 15853 9639
rect 15252 9608 15853 9636
rect 15252 9596 15258 9608
rect 15841 9605 15853 9608
rect 15887 9636 15899 9639
rect 16316 9636 16344 9676
rect 16574 9664 16580 9676
rect 16632 9664 16638 9716
rect 16850 9664 16856 9716
rect 16908 9704 16914 9716
rect 16908 9676 17264 9704
rect 16908 9664 16914 9676
rect 15887 9608 16344 9636
rect 17236 9636 17264 9676
rect 21542 9664 21548 9716
rect 21600 9704 21606 9716
rect 21729 9707 21787 9713
rect 21729 9704 21741 9707
rect 21600 9676 21741 9704
rect 21600 9664 21606 9676
rect 21729 9673 21741 9676
rect 21775 9673 21787 9707
rect 21729 9667 21787 9673
rect 22186 9664 22192 9716
rect 22244 9704 22250 9716
rect 22554 9704 22560 9716
rect 22244 9676 22560 9704
rect 22244 9664 22250 9676
rect 22554 9664 22560 9676
rect 22612 9664 22618 9716
rect 22925 9707 22983 9713
rect 22925 9673 22937 9707
rect 22971 9704 22983 9707
rect 23014 9704 23020 9716
rect 22971 9676 23020 9704
rect 22971 9673 22983 9676
rect 22925 9667 22983 9673
rect 23014 9664 23020 9676
rect 23072 9664 23078 9716
rect 25593 9707 25651 9713
rect 25593 9673 25605 9707
rect 25639 9704 25651 9707
rect 25774 9704 25780 9716
rect 25639 9676 25780 9704
rect 25639 9673 25651 9676
rect 25593 9667 25651 9673
rect 19242 9636 19248 9648
rect 17236 9608 19248 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 19242 9596 19248 9608
rect 19300 9596 19306 9648
rect 19337 9639 19395 9645
rect 19337 9605 19349 9639
rect 19383 9636 19395 9639
rect 19610 9636 19616 9648
rect 19383 9608 19616 9636
rect 19383 9605 19395 9608
rect 19337 9599 19395 9605
rect 19610 9596 19616 9608
rect 19668 9596 19674 9648
rect 21361 9639 21419 9645
rect 21361 9636 21373 9639
rect 19720 9608 21373 9636
rect 7101 9531 7159 9537
rect 7300 9540 7880 9568
rect 5074 9460 5080 9512
rect 5132 9460 5138 9512
rect 5166 9460 5172 9512
rect 5224 9460 5230 9512
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9500 5411 9503
rect 5626 9500 5632 9512
rect 5399 9472 5632 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 5626 9460 5632 9472
rect 5684 9500 5690 9512
rect 6089 9503 6147 9509
rect 6089 9500 6101 9503
rect 5684 9472 6101 9500
rect 5684 9460 5690 9472
rect 6089 9469 6101 9472
rect 6135 9500 6147 9503
rect 6181 9503 6239 9509
rect 6181 9500 6193 9503
rect 6135 9472 6193 9500
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 6181 9469 6193 9472
rect 6227 9469 6239 9503
rect 6181 9463 6239 9469
rect 6362 9460 6368 9512
rect 6420 9460 6426 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 6914 9500 6920 9512
rect 6871 9472 6920 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7300 9509 7328 9540
rect 8018 9528 8024 9580
rect 8076 9568 8082 9580
rect 13446 9568 13452 9580
rect 8076 9540 9076 9568
rect 8076 9528 8082 9540
rect 7009 9503 7067 9509
rect 7009 9469 7021 9503
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9500 7527 9503
rect 7561 9503 7619 9509
rect 7561 9500 7573 9503
rect 7515 9472 7573 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 7561 9469 7573 9472
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 3804 9404 4844 9432
rect 5092 9432 5120 9460
rect 5721 9435 5779 9441
rect 5721 9432 5733 9435
rect 5092 9404 5733 9432
rect 5721 9401 5733 9404
rect 5767 9401 5779 9435
rect 5721 9395 5779 9401
rect 5902 9392 5908 9444
rect 5960 9392 5966 9444
rect 7024 9432 7052 9463
rect 8386 9460 8392 9512
rect 8444 9460 8450 9512
rect 8570 9460 8576 9512
rect 8628 9460 8634 9512
rect 8754 9460 8760 9512
rect 8812 9460 8818 9512
rect 9048 9509 9076 9540
rect 9324 9540 13452 9568
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9500 9091 9503
rect 9214 9500 9220 9512
rect 9079 9472 9220 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 8404 9432 8432 9460
rect 7024 9404 8432 9432
rect 8864 9432 8892 9463
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 9324 9509 9352 9540
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 13998 9528 14004 9580
rect 14056 9528 14062 9580
rect 14108 9540 15884 9568
rect 9309 9503 9367 9509
rect 9309 9469 9321 9503
rect 9355 9469 9367 9503
rect 9309 9463 9367 9469
rect 9582 9460 9588 9512
rect 9640 9500 9646 9512
rect 9769 9503 9827 9509
rect 9769 9500 9781 9503
rect 9640 9472 9781 9500
rect 9640 9460 9646 9472
rect 9769 9469 9781 9472
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 11422 9460 11428 9512
rect 11480 9500 11486 9512
rect 11698 9509 11704 9512
rect 11517 9503 11575 9509
rect 11517 9500 11529 9503
rect 11480 9472 11529 9500
rect 11480 9460 11486 9472
rect 11517 9469 11529 9472
rect 11563 9469 11575 9503
rect 11517 9463 11575 9469
rect 11665 9503 11704 9509
rect 11665 9469 11677 9503
rect 11665 9463 11704 9469
rect 11698 9460 11704 9463
rect 11756 9460 11762 9512
rect 12023 9503 12081 9509
rect 12023 9469 12035 9503
rect 12069 9500 12081 9503
rect 12250 9500 12256 9512
rect 12069 9472 12256 9500
rect 12069 9469 12081 9472
rect 12023 9463 12081 9469
rect 12250 9460 12256 9472
rect 12308 9460 12314 9512
rect 12342 9460 12348 9512
rect 12400 9460 12406 9512
rect 13354 9460 13360 9512
rect 13412 9500 13418 9512
rect 14108 9500 14136 9540
rect 13412 9472 14136 9500
rect 13412 9460 13418 9472
rect 9493 9435 9551 9441
rect 8864 9404 9260 9432
rect 4246 9364 4252 9376
rect 3712 9336 4252 9364
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 4893 9367 4951 9373
rect 4893 9333 4905 9367
rect 4939 9364 4951 9367
rect 4982 9364 4988 9376
rect 4939 9336 4988 9364
rect 4939 9333 4951 9336
rect 4893 9327 4951 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5074 9324 5080 9376
rect 5132 9364 5138 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 5132 9336 5549 9364
rect 5132 9324 5138 9336
rect 5537 9333 5549 9336
rect 5583 9333 5595 9367
rect 5537 9327 5595 9333
rect 5810 9324 5816 9376
rect 5868 9324 5874 9376
rect 8389 9367 8447 9373
rect 8389 9333 8401 9367
rect 8435 9364 8447 9367
rect 8478 9364 8484 9376
rect 8435 9336 8484 9364
rect 8435 9333 8447 9336
rect 8389 9327 8447 9333
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 9122 9324 9128 9376
rect 9180 9324 9186 9376
rect 9232 9364 9260 9404
rect 9493 9401 9505 9435
rect 9539 9432 9551 9435
rect 10042 9432 10048 9444
rect 9539 9404 10048 9432
rect 9539 9401 9551 9404
rect 9493 9395 9551 9401
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 11330 9392 11336 9444
rect 11388 9432 11394 9444
rect 11790 9432 11796 9444
rect 11388 9404 11796 9432
rect 11388 9392 11394 9404
rect 11790 9392 11796 9404
rect 11848 9392 11854 9444
rect 11885 9435 11943 9441
rect 11885 9401 11897 9435
rect 11931 9401 11943 9435
rect 15654 9432 15660 9444
rect 11885 9395 11943 9401
rect 11992 9404 15660 9432
rect 9674 9364 9680 9376
rect 9232 9336 9680 9364
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 9858 9324 9864 9376
rect 9916 9364 9922 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 9916 9336 10425 9364
rect 9916 9324 9922 9336
rect 10413 9333 10425 9336
rect 10459 9364 10471 9367
rect 11900 9364 11928 9395
rect 11992 9376 12020 9404
rect 15654 9392 15660 9404
rect 15712 9392 15718 9444
rect 15746 9392 15752 9444
rect 15804 9392 15810 9444
rect 15856 9432 15884 9540
rect 18322 9528 18328 9580
rect 18380 9568 18386 9580
rect 19720 9568 19748 9608
rect 21361 9605 21373 9608
rect 21407 9605 21419 9639
rect 21361 9599 21419 9605
rect 21453 9639 21511 9645
rect 21453 9605 21465 9639
rect 21499 9636 21511 9639
rect 22830 9636 22836 9648
rect 21499 9608 22836 9636
rect 21499 9605 21511 9608
rect 21453 9599 21511 9605
rect 22830 9596 22836 9608
rect 22888 9596 22894 9648
rect 23032 9636 23060 9664
rect 23032 9608 24247 9636
rect 18380 9540 19748 9568
rect 22480 9540 23152 9568
rect 18380 9528 18386 9540
rect 22480 9512 22508 9540
rect 16482 9460 16488 9512
rect 16540 9500 16546 9512
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 16540 9472 17233 9500
rect 16540 9460 16546 9472
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 17957 9503 18015 9509
rect 17957 9469 17969 9503
rect 18003 9500 18015 9503
rect 18782 9500 18788 9512
rect 18003 9472 18788 9500
rect 18003 9469 18015 9472
rect 17957 9463 18015 9469
rect 18782 9460 18788 9472
rect 18840 9500 18846 9512
rect 18969 9503 19027 9509
rect 18969 9500 18981 9503
rect 18840 9472 18981 9500
rect 18840 9460 18846 9472
rect 18969 9469 18981 9472
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 19516 9503 19574 9509
rect 19516 9469 19528 9503
rect 19562 9500 19574 9503
rect 19562 9472 19840 9500
rect 19562 9469 19574 9472
rect 19516 9463 19574 9469
rect 16758 9432 16764 9444
rect 15856 9404 16764 9432
rect 16758 9392 16764 9404
rect 16816 9392 16822 9444
rect 16850 9392 16856 9444
rect 16908 9432 16914 9444
rect 16954 9435 17012 9441
rect 16954 9432 16966 9435
rect 16908 9404 16966 9432
rect 16908 9392 16914 9404
rect 16954 9401 16966 9404
rect 17000 9401 17012 9435
rect 19613 9435 19671 9441
rect 16954 9395 17012 9401
rect 17052 9404 19564 9432
rect 10459 9336 11928 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 11974 9324 11980 9376
rect 12032 9324 12038 9376
rect 12158 9324 12164 9376
rect 12216 9324 12222 9376
rect 12802 9324 12808 9376
rect 12860 9364 12866 9376
rect 12897 9367 12955 9373
rect 12897 9364 12909 9367
rect 12860 9336 12909 9364
rect 12860 9324 12866 9336
rect 12897 9333 12909 9336
rect 12943 9333 12955 9367
rect 12897 9327 12955 9333
rect 16114 9324 16120 9376
rect 16172 9364 16178 9376
rect 17052 9364 17080 9404
rect 19536 9376 19564 9404
rect 19613 9401 19625 9435
rect 19659 9401 19671 9435
rect 19613 9395 19671 9401
rect 16172 9336 17080 9364
rect 17773 9367 17831 9373
rect 16172 9324 16178 9336
rect 17773 9333 17785 9367
rect 17819 9364 17831 9367
rect 17862 9364 17868 9376
rect 17819 9336 17868 9364
rect 17819 9333 17831 9336
rect 17773 9327 17831 9333
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 18785 9367 18843 9373
rect 18785 9333 18797 9367
rect 18831 9364 18843 9367
rect 19242 9364 19248 9376
rect 18831 9336 19248 9364
rect 18831 9333 18843 9336
rect 18785 9327 18843 9333
rect 19242 9324 19248 9336
rect 19300 9324 19306 9376
rect 19518 9324 19524 9376
rect 19576 9324 19582 9376
rect 19628 9364 19656 9395
rect 19702 9392 19708 9444
rect 19760 9392 19766 9444
rect 19812 9432 19840 9472
rect 19886 9460 19892 9512
rect 19944 9460 19950 9512
rect 19981 9503 20039 9509
rect 19981 9469 19993 9503
rect 20027 9500 20039 9503
rect 20898 9500 20904 9512
rect 20027 9472 20904 9500
rect 20027 9469 20039 9472
rect 19981 9463 20039 9469
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 21174 9460 21180 9512
rect 21232 9500 21238 9512
rect 21269 9503 21327 9509
rect 21269 9500 21281 9503
rect 21232 9472 21281 9500
rect 21232 9460 21238 9472
rect 21269 9469 21281 9472
rect 21315 9469 21327 9503
rect 21269 9463 21327 9469
rect 21450 9460 21456 9512
rect 21508 9500 21514 9512
rect 21545 9503 21603 9509
rect 21545 9500 21557 9503
rect 21508 9472 21557 9500
rect 21508 9460 21514 9472
rect 21545 9469 21557 9472
rect 21591 9500 21603 9503
rect 22005 9503 22063 9509
rect 22005 9500 22017 9503
rect 21591 9472 22017 9500
rect 21591 9469 21603 9472
rect 21545 9463 21603 9469
rect 22005 9469 22017 9472
rect 22051 9469 22063 9503
rect 22005 9463 22063 9469
rect 22186 9460 22192 9512
rect 22244 9460 22250 9512
rect 22373 9503 22431 9509
rect 22373 9469 22385 9503
rect 22419 9469 22431 9503
rect 22373 9463 22431 9469
rect 20162 9432 20168 9444
rect 19812 9404 20168 9432
rect 20162 9392 20168 9404
rect 20220 9392 20226 9444
rect 22388 9432 22416 9463
rect 22462 9460 22468 9512
rect 22520 9460 22526 9512
rect 23124 9509 23152 9540
rect 24026 9509 24032 9512
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9469 22983 9503
rect 22925 9463 22983 9469
rect 23109 9503 23167 9509
rect 23109 9469 23121 9503
rect 23155 9500 23167 9503
rect 23845 9503 23903 9509
rect 23845 9500 23857 9503
rect 23155 9472 23857 9500
rect 23155 9469 23167 9472
rect 23109 9463 23167 9469
rect 23845 9469 23857 9472
rect 23891 9469 23903 9503
rect 23845 9463 23903 9469
rect 24003 9503 24032 9509
rect 24003 9469 24015 9503
rect 24003 9463 24032 9469
rect 22940 9432 22968 9463
rect 24026 9460 24032 9463
rect 24084 9460 24090 9512
rect 24121 9503 24179 9509
rect 24121 9469 24133 9503
rect 24167 9500 24179 9503
rect 24219 9500 24247 9608
rect 24394 9528 24400 9580
rect 24452 9568 24458 9580
rect 24581 9571 24639 9577
rect 24581 9568 24593 9571
rect 24452 9540 24593 9568
rect 24452 9528 24458 9540
rect 24581 9537 24593 9540
rect 24627 9537 24639 9571
rect 24946 9568 24952 9580
rect 24581 9531 24639 9537
rect 24780 9540 24952 9568
rect 24167 9472 24247 9500
rect 24305 9503 24363 9509
rect 24167 9469 24179 9472
rect 24121 9463 24179 9469
rect 24305 9469 24317 9503
rect 24351 9469 24363 9503
rect 24305 9463 24363 9469
rect 22388 9404 24072 9432
rect 24044 9376 24072 9404
rect 24210 9392 24216 9444
rect 24268 9392 24274 9444
rect 24320 9432 24348 9463
rect 24486 9460 24492 9512
rect 24544 9460 24550 9512
rect 24780 9509 24808 9540
rect 24946 9528 24952 9540
rect 25004 9568 25010 9580
rect 25608 9568 25636 9667
rect 25774 9664 25780 9676
rect 25832 9664 25838 9716
rect 26786 9568 26792 9580
rect 25004 9540 25636 9568
rect 25700 9540 26792 9568
rect 25004 9528 25010 9540
rect 24765 9503 24823 9509
rect 24765 9469 24777 9503
rect 24811 9469 24823 9503
rect 24765 9463 24823 9469
rect 24854 9460 24860 9512
rect 24912 9500 24918 9512
rect 25041 9503 25099 9509
rect 25041 9500 25053 9503
rect 24912 9472 25053 9500
rect 24912 9460 24918 9472
rect 25041 9469 25053 9472
rect 25087 9469 25099 9503
rect 25041 9463 25099 9469
rect 25314 9460 25320 9512
rect 25372 9460 25378 9512
rect 25700 9509 25728 9540
rect 26786 9528 26792 9540
rect 26844 9528 26850 9580
rect 25685 9503 25743 9509
rect 25685 9469 25697 9503
rect 25731 9469 25743 9503
rect 25685 9463 25743 9469
rect 25774 9460 25780 9512
rect 25832 9460 25838 9512
rect 25869 9435 25927 9441
rect 25869 9432 25881 9435
rect 24320 9404 25881 9432
rect 25424 9376 25452 9404
rect 25869 9401 25881 9404
rect 25915 9401 25927 9435
rect 25869 9395 25927 9401
rect 21082 9364 21088 9376
rect 19628 9336 21088 9364
rect 21082 9324 21088 9336
rect 21140 9324 21146 9376
rect 24026 9324 24032 9376
rect 24084 9364 24090 9376
rect 24949 9367 25007 9373
rect 24949 9364 24961 9367
rect 24084 9336 24961 9364
rect 24084 9324 24090 9336
rect 24949 9333 24961 9336
rect 24995 9333 25007 9367
rect 24949 9327 25007 9333
rect 25133 9367 25191 9373
rect 25133 9333 25145 9367
rect 25179 9364 25191 9367
rect 25314 9364 25320 9376
rect 25179 9336 25320 9364
rect 25179 9333 25191 9336
rect 25133 9327 25191 9333
rect 25314 9324 25320 9336
rect 25372 9324 25378 9376
rect 25406 9324 25412 9376
rect 25464 9324 25470 9376
rect 552 9274 27576 9296
rect 552 9222 7114 9274
rect 7166 9222 7178 9274
rect 7230 9222 7242 9274
rect 7294 9222 7306 9274
rect 7358 9222 7370 9274
rect 7422 9222 13830 9274
rect 13882 9222 13894 9274
rect 13946 9222 13958 9274
rect 14010 9222 14022 9274
rect 14074 9222 14086 9274
rect 14138 9222 20546 9274
rect 20598 9222 20610 9274
rect 20662 9222 20674 9274
rect 20726 9222 20738 9274
rect 20790 9222 20802 9274
rect 20854 9222 27262 9274
rect 27314 9222 27326 9274
rect 27378 9222 27390 9274
rect 27442 9222 27454 9274
rect 27506 9222 27518 9274
rect 27570 9222 27576 9274
rect 552 9200 27576 9222
rect 2869 9163 2927 9169
rect 2869 9129 2881 9163
rect 2915 9160 2927 9163
rect 3786 9160 3792 9172
rect 2915 9132 3792 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 5626 9120 5632 9172
rect 5684 9120 5690 9172
rect 6549 9163 6607 9169
rect 6549 9129 6561 9163
rect 6595 9160 6607 9163
rect 8754 9160 8760 9172
rect 6595 9132 8760 9160
rect 6595 9129 6607 9132
rect 6549 9123 6607 9129
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 9582 9120 9588 9172
rect 9640 9120 9646 9172
rect 9674 9120 9680 9172
rect 9732 9120 9738 9172
rect 11974 9160 11980 9172
rect 9784 9132 11980 9160
rect 1756 9095 1814 9101
rect 1756 9061 1768 9095
rect 1802 9092 1814 9095
rect 1946 9092 1952 9104
rect 1802 9064 1952 9092
rect 1802 9061 1814 9064
rect 1756 9055 1814 9061
rect 1946 9052 1952 9064
rect 2004 9052 2010 9104
rect 3050 9052 3056 9104
rect 3108 9092 3114 9104
rect 4430 9092 4436 9104
rect 3108 9064 4436 9092
rect 3108 9052 3114 9064
rect 4430 9052 4436 9064
rect 4488 9052 4494 9104
rect 5166 9052 5172 9104
rect 5224 9092 5230 9104
rect 5810 9092 5816 9104
rect 5224 9064 5816 9092
rect 5224 9052 5230 9064
rect 5810 9052 5816 9064
rect 5868 9052 5874 9104
rect 9122 9092 9128 9104
rect 7668 9064 9128 9092
rect 4516 9027 4574 9033
rect 4516 8993 4528 9027
rect 4562 9024 4574 9027
rect 5258 9024 5264 9036
rect 4562 8996 5264 9024
rect 4562 8993 4574 8996
rect 4516 8987 4574 8993
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 6362 8984 6368 9036
rect 6420 8984 6426 9036
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 7668 9033 7696 9064
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 9214 9052 9220 9104
rect 9272 9092 9278 9104
rect 9784 9092 9812 9132
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12342 9120 12348 9172
rect 12400 9120 12406 9172
rect 12621 9163 12679 9169
rect 12621 9129 12633 9163
rect 12667 9160 12679 9163
rect 12986 9160 12992 9172
rect 12667 9132 12992 9160
rect 12667 9129 12679 9132
rect 12621 9123 12679 9129
rect 12986 9120 12992 9132
rect 13044 9120 13050 9172
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 13504 9132 16528 9160
rect 13504 9120 13510 9132
rect 9272 9064 9812 9092
rect 9272 9052 9278 9064
rect 9858 9052 9864 9104
rect 9916 9052 9922 9104
rect 10042 9052 10048 9104
rect 10100 9052 10106 9104
rect 10152 9064 11376 9092
rect 7469 9027 7527 9033
rect 7469 9024 7481 9027
rect 6972 8996 7481 9024
rect 6972 8984 6978 8996
rect 7469 8993 7481 8996
rect 7515 8993 7527 9027
rect 7469 8987 7527 8993
rect 7653 9027 7711 9033
rect 7653 8993 7665 9027
rect 7699 8993 7711 9027
rect 7653 8987 7711 8993
rect 1486 8916 1492 8968
rect 1544 8916 1550 8968
rect 4246 8916 4252 8968
rect 4304 8916 4310 8968
rect 6086 8916 6092 8968
rect 6144 8956 6150 8968
rect 6181 8959 6239 8965
rect 6181 8956 6193 8959
rect 6144 8928 6193 8956
rect 6144 8916 6150 8928
rect 6181 8925 6193 8928
rect 6227 8925 6239 8959
rect 7484 8956 7512 8987
rect 7834 8984 7840 9036
rect 7892 8984 7898 9036
rect 7929 9027 7987 9033
rect 7929 8993 7941 9027
rect 7975 9024 7987 9027
rect 8110 9024 8116 9036
rect 7975 8996 8116 9024
rect 7975 8993 7987 8996
rect 7929 8987 7987 8993
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 8205 9027 8263 9033
rect 8205 8993 8217 9027
rect 8251 9024 8263 9027
rect 8294 9024 8300 9036
rect 8251 8996 8300 9024
rect 8251 8993 8263 8996
rect 8205 8987 8263 8993
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 8478 9033 8484 9036
rect 8472 9024 8484 9033
rect 8439 8996 8484 9024
rect 8472 8987 8484 8996
rect 8478 8984 8484 8987
rect 8536 8984 8542 9036
rect 10152 9024 10180 9064
rect 11238 9033 11244 9036
rect 9232 8996 10180 9024
rect 8018 8956 8024 8968
rect 7484 8928 8024 8956
rect 6181 8919 6239 8925
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 7745 8891 7803 8897
rect 7745 8888 7757 8891
rect 7064 8860 7757 8888
rect 7064 8848 7070 8860
rect 7745 8857 7757 8860
rect 7791 8857 7803 8891
rect 7745 8851 7803 8857
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 6270 8820 6276 8832
rect 4488 8792 6276 8820
rect 4488 8780 4494 8792
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 8110 8780 8116 8832
rect 8168 8780 8174 8832
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 9232 8820 9260 8996
rect 11232 8987 11244 9033
rect 11238 8984 11244 8987
rect 11296 8984 11302 9036
rect 11348 9024 11376 9064
rect 11514 9052 11520 9104
rect 11572 9092 11578 9104
rect 11882 9092 11888 9104
rect 11572 9064 11888 9092
rect 11572 9052 11578 9064
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 12158 9052 12164 9104
rect 12216 9092 12222 9104
rect 13998 9092 14004 9104
rect 12216 9064 13768 9092
rect 12216 9052 12222 9064
rect 12437 9027 12495 9033
rect 12437 9024 12449 9027
rect 11348 8996 12449 9024
rect 12437 8993 12449 8996
rect 12483 9024 12495 9027
rect 13170 9024 13176 9036
rect 12483 8996 13176 9024
rect 12483 8993 12495 8996
rect 12437 8987 12495 8993
rect 13170 8984 13176 8996
rect 13228 8984 13234 9036
rect 13538 8984 13544 9036
rect 13596 8984 13602 9036
rect 13740 9033 13768 9064
rect 13832 9064 14004 9092
rect 13832 9033 13860 9064
rect 13998 9052 14004 9064
rect 14056 9052 14062 9104
rect 14185 9095 14243 9101
rect 14185 9061 14197 9095
rect 14231 9092 14243 9095
rect 14522 9095 14580 9101
rect 14522 9092 14534 9095
rect 14231 9064 14534 9092
rect 14231 9061 14243 9064
rect 14185 9055 14243 9061
rect 14522 9061 14534 9064
rect 14568 9061 14580 9095
rect 14522 9055 14580 9061
rect 14734 9052 14740 9104
rect 14792 9052 14798 9104
rect 16500 9101 16528 9132
rect 16850 9120 16856 9172
rect 16908 9120 16914 9172
rect 19058 9160 19064 9172
rect 17236 9132 19064 9160
rect 16485 9095 16543 9101
rect 16485 9061 16497 9095
rect 16531 9061 16543 9095
rect 16485 9055 16543 9061
rect 16758 9052 16764 9104
rect 16816 9092 16822 9104
rect 17236 9092 17264 9132
rect 19058 9120 19064 9132
rect 19116 9120 19122 9172
rect 24486 9160 24492 9172
rect 19812 9132 24492 9160
rect 18414 9092 18420 9104
rect 16816 9064 17264 9092
rect 16816 9052 16822 9064
rect 13725 9027 13783 9033
rect 13725 8993 13737 9027
rect 13771 8993 13783 9027
rect 13725 8987 13783 8993
rect 13817 9027 13875 9033
rect 13817 8993 13829 9027
rect 13863 8993 13875 9027
rect 13817 8987 13875 8993
rect 13909 9027 13967 9033
rect 13909 8993 13921 9027
rect 13955 8993 13967 9027
rect 13909 8987 13967 8993
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 9732 8928 10977 8956
rect 9732 8916 9738 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 12216 8928 12817 8956
rect 12216 8916 12222 8928
rect 12805 8925 12817 8928
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 12894 8916 12900 8968
rect 12952 8956 12958 8968
rect 13262 8956 13268 8968
rect 12952 8928 13268 8956
rect 12952 8916 12958 8928
rect 13262 8916 13268 8928
rect 13320 8956 13326 8968
rect 13832 8956 13860 8987
rect 13320 8928 13860 8956
rect 13924 8956 13952 8987
rect 14274 8984 14280 9036
rect 14332 8984 14338 9036
rect 14752 9024 14780 9052
rect 14384 8996 15332 9024
rect 14384 8956 14412 8996
rect 13924 8928 14412 8956
rect 13320 8916 13326 8928
rect 9306 8848 9312 8900
rect 9364 8888 9370 8900
rect 10134 8888 10140 8900
rect 9364 8860 10140 8888
rect 9364 8848 9370 8860
rect 10134 8848 10140 8860
rect 10192 8888 10198 8900
rect 10502 8888 10508 8900
rect 10192 8860 10508 8888
rect 10192 8848 10198 8860
rect 10502 8848 10508 8860
rect 10560 8848 10566 8900
rect 11974 8848 11980 8900
rect 12032 8888 12038 8900
rect 15304 8888 15332 8996
rect 16114 8984 16120 9036
rect 16172 8984 16178 9036
rect 16210 9027 16268 9033
rect 16210 8993 16222 9027
rect 16256 8993 16268 9027
rect 16210 8987 16268 8993
rect 16224 8956 16252 8987
rect 16298 8984 16304 9036
rect 16356 9024 16362 9036
rect 16393 9027 16451 9033
rect 16393 9024 16405 9027
rect 16356 8996 16405 9024
rect 16356 8984 16362 8996
rect 16393 8993 16405 8996
rect 16439 8993 16451 9027
rect 16393 8987 16451 8993
rect 16623 9027 16681 9033
rect 16623 8993 16635 9027
rect 16669 9024 16681 9027
rect 16850 9024 16856 9036
rect 16669 8996 16856 9024
rect 16669 8993 16681 8996
rect 16623 8987 16681 8993
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 17126 8984 17132 9036
rect 17184 8984 17190 9036
rect 17236 9033 17264 9064
rect 17512 9064 18420 9092
rect 17512 9033 17540 9064
rect 18414 9052 18420 9064
rect 18472 9052 18478 9104
rect 17221 9027 17279 9033
rect 17221 8993 17233 9027
rect 17267 8993 17279 9027
rect 17221 8987 17279 8993
rect 17313 9027 17371 9033
rect 17313 8993 17325 9027
rect 17359 8993 17371 9027
rect 17313 8987 17371 8993
rect 17497 9027 17555 9033
rect 17497 8993 17509 9027
rect 17543 8993 17555 9027
rect 17497 8987 17555 8993
rect 17589 9027 17647 9033
rect 17589 8993 17601 9027
rect 17635 9024 17647 9027
rect 17678 9024 17684 9036
rect 17635 8996 17684 9024
rect 17635 8993 17647 8996
rect 17589 8987 17647 8993
rect 17328 8956 17356 8987
rect 17678 8984 17684 8996
rect 17736 8984 17742 9036
rect 17862 8984 17868 9036
rect 17920 9024 17926 9036
rect 17957 9027 18015 9033
rect 17957 9024 17969 9027
rect 17920 8996 17969 9024
rect 17920 8984 17926 8996
rect 17957 8993 17969 8996
rect 18003 8993 18015 9027
rect 17957 8987 18015 8993
rect 18322 8984 18328 9036
rect 18380 8984 18386 9036
rect 18509 9027 18567 9033
rect 18509 8993 18521 9027
rect 18555 9024 18567 9027
rect 19150 9024 19156 9036
rect 18555 8996 19156 9024
rect 18555 8993 18567 8996
rect 18509 8987 18567 8993
rect 19150 8984 19156 8996
rect 19208 8984 19214 9036
rect 19242 8984 19248 9036
rect 19300 9024 19306 9036
rect 19812 9033 19840 9132
rect 24486 9120 24492 9132
rect 24544 9120 24550 9172
rect 24578 9120 24584 9172
rect 24636 9160 24642 9172
rect 24636 9132 25268 9160
rect 24636 9120 24642 9132
rect 21542 9092 21548 9104
rect 20364 9064 21548 9092
rect 20364 9033 20392 9064
rect 21542 9052 21548 9064
rect 21600 9092 21606 9104
rect 21818 9092 21824 9104
rect 21600 9064 21824 9092
rect 21600 9052 21606 9064
rect 21818 9052 21824 9064
rect 21876 9052 21882 9104
rect 24946 9092 24952 9104
rect 24780 9064 24952 9092
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 19300 8996 19625 9024
rect 19300 8984 19306 8996
rect 19613 8993 19625 8996
rect 19659 8993 19671 9027
rect 19613 8987 19671 8993
rect 19797 9027 19855 9033
rect 19797 8993 19809 9027
rect 19843 8993 19855 9027
rect 19797 8987 19855 8993
rect 20349 9027 20407 9033
rect 20349 8993 20361 9027
rect 20395 8993 20407 9027
rect 20349 8987 20407 8993
rect 20441 9027 20499 9033
rect 20441 8993 20453 9027
rect 20487 8993 20499 9027
rect 20441 8987 20499 8993
rect 18046 8956 18052 8968
rect 15672 8928 16252 8956
rect 16776 8928 17356 8956
rect 17788 8928 18052 8956
rect 15672 8897 15700 8928
rect 16776 8897 16804 8928
rect 17788 8897 17816 8928
rect 18046 8916 18052 8928
rect 18104 8956 18110 8968
rect 18340 8956 18368 8984
rect 18104 8928 18368 8956
rect 19981 8959 20039 8965
rect 18104 8916 18110 8928
rect 19981 8925 19993 8959
rect 20027 8956 20039 8959
rect 20456 8956 20484 8987
rect 22462 8984 22468 9036
rect 22520 9024 22526 9036
rect 24780 9033 24808 9064
rect 24946 9052 24952 9064
rect 25004 9052 25010 9104
rect 23661 9027 23719 9033
rect 23661 9024 23673 9027
rect 22520 8996 23673 9024
rect 22520 8984 22526 8996
rect 23661 8993 23673 8996
rect 23707 8993 23719 9027
rect 23661 8987 23719 8993
rect 24673 9027 24731 9033
rect 24673 8993 24685 9027
rect 24719 8993 24731 9027
rect 24673 8987 24731 8993
rect 24765 9027 24823 9033
rect 24765 8993 24777 9027
rect 24811 8993 24823 9027
rect 24765 8987 24823 8993
rect 20027 8928 20484 8956
rect 24121 8959 24179 8965
rect 20027 8925 20039 8928
rect 19981 8919 20039 8925
rect 24121 8925 24133 8959
rect 24167 8956 24179 8959
rect 24302 8956 24308 8968
rect 24167 8928 24308 8956
rect 24167 8925 24179 8928
rect 24121 8919 24179 8925
rect 24302 8916 24308 8928
rect 24360 8916 24366 8968
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8925 24639 8959
rect 24688 8956 24716 8987
rect 24854 8984 24860 9036
rect 24912 9024 24918 9036
rect 25041 9027 25099 9033
rect 25041 9024 25053 9027
rect 24912 8996 25053 9024
rect 24912 8984 24918 8996
rect 25041 8993 25053 8996
rect 25087 8993 25099 9027
rect 25041 8987 25099 8993
rect 25130 8984 25136 9036
rect 25188 8984 25194 9036
rect 25240 8956 25268 9132
rect 26421 9095 26479 9101
rect 26421 9092 26433 9095
rect 25516 9064 26433 9092
rect 25314 8984 25320 9036
rect 25372 8984 25378 9036
rect 25406 8984 25412 9036
rect 25464 8984 25470 9036
rect 25516 9033 25544 9064
rect 26421 9061 26433 9064
rect 26467 9061 26479 9095
rect 26421 9055 26479 9061
rect 25501 9027 25559 9033
rect 25501 8993 25513 9027
rect 25547 8993 25559 9027
rect 25501 8987 25559 8993
rect 25590 8984 25596 9036
rect 25648 9024 25654 9036
rect 25774 9024 25780 9036
rect 25648 8996 25780 9024
rect 25648 8984 25654 8996
rect 25774 8984 25780 8996
rect 25832 9024 25838 9036
rect 25869 9027 25927 9033
rect 25869 9024 25881 9027
rect 25832 8996 25881 9024
rect 25832 8984 25838 8996
rect 25869 8993 25881 8996
rect 25915 8993 25927 9027
rect 25869 8987 25927 8993
rect 25958 8984 25964 9036
rect 26016 9024 26022 9036
rect 26053 9027 26111 9033
rect 26053 9024 26065 9027
rect 26016 8996 26065 9024
rect 26016 8984 26022 8996
rect 26053 8993 26065 8996
rect 26099 8993 26111 9027
rect 26053 8987 26111 8993
rect 26145 9027 26203 9033
rect 26145 8993 26157 9027
rect 26191 8993 26203 9027
rect 26145 8987 26203 8993
rect 26160 8956 26188 8987
rect 24688 8928 24900 8956
rect 25240 8928 26188 8956
rect 24581 8919 24639 8925
rect 15657 8891 15715 8897
rect 15657 8888 15669 8891
rect 12032 8860 14320 8888
rect 15304 8860 15669 8888
rect 12032 8848 12038 8860
rect 8260 8792 9260 8820
rect 8260 8780 8266 8792
rect 11606 8780 11612 8832
rect 11664 8820 11670 8832
rect 12526 8820 12532 8832
rect 11664 8792 12532 8820
rect 11664 8780 11670 8792
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 14292 8820 14320 8860
rect 15657 8857 15669 8860
rect 15703 8857 15715 8891
rect 15657 8851 15715 8857
rect 16761 8891 16819 8897
rect 16761 8857 16773 8891
rect 16807 8857 16819 8891
rect 16761 8851 16819 8857
rect 17773 8891 17831 8897
rect 17773 8857 17785 8891
rect 17819 8857 17831 8891
rect 17773 8851 17831 8857
rect 17954 8848 17960 8900
rect 18012 8888 18018 8900
rect 18417 8891 18475 8897
rect 18417 8888 18429 8891
rect 18012 8860 18429 8888
rect 18012 8848 18018 8860
rect 18417 8857 18429 8860
rect 18463 8857 18475 8891
rect 18417 8851 18475 8857
rect 19518 8848 19524 8900
rect 19576 8888 19582 8900
rect 20165 8891 20223 8897
rect 20165 8888 20177 8891
rect 19576 8860 20177 8888
rect 19576 8848 19582 8860
rect 20165 8857 20177 8860
rect 20211 8857 20223 8891
rect 24486 8888 24492 8900
rect 20165 8851 20223 8857
rect 23952 8860 24492 8888
rect 16942 8820 16948 8832
rect 14292 8792 16948 8820
rect 16942 8780 16948 8792
rect 17000 8820 17006 8832
rect 18141 8823 18199 8829
rect 18141 8820 18153 8823
rect 17000 8792 18153 8820
rect 17000 8780 17006 8792
rect 18141 8789 18153 8792
rect 18187 8789 18199 8823
rect 18141 8783 18199 8789
rect 20622 8780 20628 8832
rect 20680 8780 20686 8832
rect 23952 8829 23980 8860
rect 24486 8848 24492 8860
rect 24544 8888 24550 8900
rect 24596 8888 24624 8919
rect 24872 8897 24900 8928
rect 26786 8916 26792 8968
rect 26844 8956 26850 8968
rect 26973 8959 27031 8965
rect 26973 8956 26985 8959
rect 26844 8928 26985 8956
rect 26844 8916 26850 8928
rect 26973 8925 26985 8928
rect 27019 8925 27031 8959
rect 26973 8919 27031 8925
rect 24544 8860 24624 8888
rect 24857 8891 24915 8897
rect 24544 8848 24550 8860
rect 24857 8857 24869 8891
rect 24903 8888 24915 8891
rect 25958 8888 25964 8900
rect 24903 8860 25964 8888
rect 24903 8857 24915 8860
rect 24857 8851 24915 8857
rect 25958 8848 25964 8860
rect 26016 8848 26022 8900
rect 23937 8823 23995 8829
rect 23937 8789 23949 8823
rect 23983 8789 23995 8823
rect 23937 8783 23995 8789
rect 24026 8780 24032 8832
rect 24084 8820 24090 8832
rect 24305 8823 24363 8829
rect 24305 8820 24317 8823
rect 24084 8792 24317 8820
rect 24084 8780 24090 8792
rect 24305 8789 24317 8792
rect 24351 8789 24363 8823
rect 24305 8783 24363 8789
rect 24670 8780 24676 8832
rect 24728 8780 24734 8832
rect 24762 8780 24768 8832
rect 24820 8780 24826 8832
rect 25774 8780 25780 8832
rect 25832 8780 25838 8832
rect 25866 8780 25872 8832
rect 25924 8780 25930 8832
rect 552 8730 27416 8752
rect 552 8678 3756 8730
rect 3808 8678 3820 8730
rect 3872 8678 3884 8730
rect 3936 8678 3948 8730
rect 4000 8678 4012 8730
rect 4064 8678 10472 8730
rect 10524 8678 10536 8730
rect 10588 8678 10600 8730
rect 10652 8678 10664 8730
rect 10716 8678 10728 8730
rect 10780 8678 17188 8730
rect 17240 8678 17252 8730
rect 17304 8678 17316 8730
rect 17368 8678 17380 8730
rect 17432 8678 17444 8730
rect 17496 8678 23904 8730
rect 23956 8678 23968 8730
rect 24020 8678 24032 8730
rect 24084 8678 24096 8730
rect 24148 8678 24160 8730
rect 24212 8678 27416 8730
rect 552 8656 27416 8678
rect 4798 8616 4804 8628
rect 3252 8588 4804 8616
rect 3252 8480 3280 8588
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 4985 8619 5043 8625
rect 4985 8585 4997 8619
rect 5031 8616 5043 8619
rect 5031 8588 5304 8616
rect 5031 8585 5043 8588
rect 4985 8579 5043 8585
rect 3329 8551 3387 8557
rect 3329 8517 3341 8551
rect 3375 8548 3387 8551
rect 4154 8548 4160 8560
rect 3375 8520 4160 8548
rect 3375 8517 3387 8520
rect 3329 8511 3387 8517
rect 4154 8508 4160 8520
rect 4212 8548 4218 8560
rect 4617 8551 4675 8557
rect 4617 8548 4629 8551
rect 4212 8520 4629 8548
rect 4212 8508 4218 8520
rect 4617 8517 4629 8520
rect 4663 8548 4675 8551
rect 5074 8548 5080 8560
rect 4663 8520 5080 8548
rect 4663 8517 4675 8520
rect 4617 8511 4675 8517
rect 5074 8508 5080 8520
rect 5132 8508 5138 8560
rect 5169 8551 5227 8557
rect 5169 8517 5181 8551
rect 5215 8517 5227 8551
rect 5276 8548 5304 8588
rect 7006 8576 7012 8628
rect 7064 8576 7070 8628
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 7883 8588 9812 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 6638 8548 6644 8560
rect 5276 8520 6644 8548
rect 5169 8511 5227 8517
rect 3513 8483 3571 8489
rect 3513 8480 3525 8483
rect 3252 8452 3525 8480
rect 3513 8449 3525 8452
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 4062 8440 4068 8492
rect 4120 8480 4126 8492
rect 4249 8483 4307 8489
rect 4249 8480 4261 8483
rect 4120 8452 4261 8480
rect 4120 8440 4126 8452
rect 4249 8449 4261 8452
rect 4295 8480 4307 8483
rect 4295 8452 5120 8480
rect 4295 8449 4307 8452
rect 4249 8443 4307 8449
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 4341 8415 4399 8421
rect 4341 8381 4353 8415
rect 4387 8381 4399 8415
rect 4341 8375 4399 8381
rect 3252 8344 3280 8375
rect 3605 8347 3663 8353
rect 3605 8344 3617 8347
rect 3252 8316 3617 8344
rect 3605 8313 3617 8316
rect 3651 8313 3663 8347
rect 4356 8344 4384 8375
rect 4522 8372 4528 8424
rect 4580 8372 4586 8424
rect 4706 8344 4712 8356
rect 4356 8316 4712 8344
rect 3605 8307 3663 8313
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 4982 8304 4988 8356
rect 5040 8304 5046 8356
rect 5092 8344 5120 8452
rect 5184 8412 5212 8511
rect 6638 8508 6644 8520
rect 6696 8508 6702 8560
rect 9784 8548 9812 8588
rect 11238 8576 11244 8628
rect 11296 8576 11302 8628
rect 13541 8619 13599 8625
rect 13541 8616 13553 8619
rect 11716 8588 13553 8616
rect 11609 8551 11667 8557
rect 11609 8548 11621 8551
rect 9784 8520 11621 8548
rect 11609 8517 11621 8520
rect 11655 8517 11667 8551
rect 11609 8511 11667 8517
rect 6362 8440 6368 8492
rect 6420 8480 6426 8492
rect 6420 8452 7696 8480
rect 6420 8440 6426 8452
rect 5445 8415 5503 8421
rect 5445 8412 5457 8415
rect 5184 8384 5457 8412
rect 5445 8381 5457 8384
rect 5491 8381 5503 8415
rect 5445 8375 5503 8381
rect 5902 8372 5908 8424
rect 5960 8372 5966 8424
rect 6840 8421 6868 8452
rect 6457 8415 6515 8421
rect 6457 8381 6469 8415
rect 6503 8412 6515 8415
rect 6641 8415 6699 8421
rect 6641 8412 6653 8415
rect 6503 8384 6653 8412
rect 6503 8381 6515 8384
rect 6457 8375 6515 8381
rect 6641 8381 6653 8384
rect 6687 8381 6699 8415
rect 6641 8375 6699 8381
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 7466 8372 7472 8424
rect 7524 8372 7530 8424
rect 7668 8421 7696 8452
rect 9582 8440 9588 8492
rect 9640 8480 9646 8492
rect 9640 8452 11468 8480
rect 9640 8440 9646 8452
rect 11440 8424 11468 8452
rect 7653 8415 7711 8421
rect 7653 8381 7665 8415
rect 7699 8412 7711 8415
rect 8202 8412 8208 8424
rect 7699 8384 8208 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 8389 8415 8447 8421
rect 8389 8381 8401 8415
rect 8435 8412 8447 8415
rect 9674 8412 9680 8424
rect 8435 8384 9680 8412
rect 8435 8381 8447 8384
rect 8389 8375 8447 8381
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 11422 8372 11428 8424
rect 11480 8372 11486 8424
rect 11517 8415 11575 8421
rect 11517 8381 11529 8415
rect 11563 8412 11575 8415
rect 11606 8412 11612 8424
rect 11563 8384 11612 8412
rect 11563 8381 11575 8384
rect 11517 8375 11575 8381
rect 11606 8372 11612 8384
rect 11664 8372 11670 8424
rect 11716 8421 11744 8588
rect 13541 8585 13553 8588
rect 13587 8585 13599 8619
rect 13541 8579 13599 8585
rect 13630 8576 13636 8628
rect 13688 8616 13694 8628
rect 14185 8619 14243 8625
rect 14185 8616 14197 8619
rect 13688 8588 14197 8616
rect 13688 8576 13694 8588
rect 14185 8585 14197 8588
rect 14231 8616 14243 8619
rect 17313 8619 17371 8625
rect 14231 8588 15608 8616
rect 14231 8585 14243 8588
rect 14185 8579 14243 8585
rect 12710 8508 12716 8560
rect 12768 8508 12774 8560
rect 15580 8548 15608 8588
rect 17313 8585 17325 8619
rect 17359 8616 17371 8619
rect 17586 8616 17592 8628
rect 17359 8588 17592 8616
rect 17359 8585 17371 8588
rect 17313 8579 17371 8585
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 19334 8616 19340 8628
rect 18708 8588 19340 8616
rect 18138 8548 18144 8560
rect 13372 8520 14412 8548
rect 15580 8520 18144 8548
rect 12158 8480 12164 8492
rect 11808 8452 12164 8480
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8381 11759 8415
rect 11701 8375 11759 8381
rect 6086 8344 6092 8356
rect 5092 8316 6092 8344
rect 6086 8304 6092 8316
rect 6144 8304 6150 8356
rect 8110 8304 8116 8356
rect 8168 8344 8174 8356
rect 8634 8347 8692 8353
rect 8634 8344 8646 8347
rect 8168 8316 8646 8344
rect 8168 8304 8174 8316
rect 8634 8313 8646 8316
rect 8680 8313 8692 8347
rect 11808 8344 11836 8452
rect 12158 8440 12164 8452
rect 12216 8440 12222 8492
rect 12250 8440 12256 8492
rect 12308 8440 12314 8492
rect 11882 8372 11888 8424
rect 11940 8372 11946 8424
rect 11977 8415 12035 8421
rect 11977 8381 11989 8415
rect 12023 8381 12035 8415
rect 11977 8375 12035 8381
rect 8634 8307 8692 8313
rect 9784 8316 11836 8344
rect 11992 8344 12020 8375
rect 12066 8372 12072 8424
rect 12124 8372 12130 8424
rect 12268 8412 12296 8440
rect 12728 8421 12756 8508
rect 13372 8489 13400 8520
rect 13357 8483 13415 8489
rect 13357 8449 13369 8483
rect 13403 8449 13415 8483
rect 13357 8443 13415 8449
rect 12442 8415 12500 8421
rect 12442 8412 12454 8415
rect 12176 8384 12454 8412
rect 12176 8356 12204 8384
rect 12442 8381 12454 8384
rect 12488 8381 12500 8415
rect 12728 8415 12795 8421
rect 12728 8384 12749 8415
rect 12442 8375 12500 8381
rect 12737 8381 12749 8384
rect 12783 8381 12795 8415
rect 12737 8375 12795 8381
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8381 12955 8415
rect 12989 8415 13047 8421
rect 12989 8412 13001 8415
rect 12897 8375 12955 8381
rect 12984 8381 13001 8412
rect 13035 8381 13047 8415
rect 13127 8415 13185 8421
rect 13127 8412 13139 8415
rect 12984 8375 13047 8381
rect 13116 8381 13139 8412
rect 13173 8406 13185 8415
rect 13446 8406 13452 8424
rect 13173 8390 13308 8406
rect 13372 8390 13452 8406
rect 13173 8381 13452 8390
rect 13116 8378 13452 8381
rect 13127 8375 13185 8378
rect 11992 8316 12066 8344
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 3513 8279 3571 8285
rect 3513 8276 3525 8279
rect 3476 8248 3525 8276
rect 3476 8236 3482 8248
rect 3513 8245 3525 8248
rect 3559 8245 3571 8279
rect 3513 8239 3571 8245
rect 4430 8236 4436 8288
rect 4488 8236 4494 8288
rect 5258 8236 5264 8288
rect 5316 8236 5322 8288
rect 9784 8285 9812 8316
rect 9769 8279 9827 8285
rect 9769 8245 9781 8279
rect 9815 8245 9827 8279
rect 9769 8239 9827 8245
rect 11330 8236 11336 8288
rect 11388 8276 11394 8288
rect 12038 8276 12066 8316
rect 12158 8304 12164 8356
rect 12216 8304 12222 8356
rect 12250 8304 12256 8356
rect 12308 8304 12314 8356
rect 12342 8304 12348 8356
rect 12400 8304 12406 8356
rect 12526 8276 12532 8288
rect 11388 8248 12532 8276
rect 11388 8236 11394 8248
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 12621 8279 12679 8285
rect 12621 8245 12633 8279
rect 12667 8276 12679 8279
rect 12912 8276 12940 8375
rect 12667 8248 12940 8276
rect 12984 8276 13012 8375
rect 13280 8362 13400 8378
rect 13446 8372 13452 8378
rect 13504 8372 13510 8424
rect 14384 8412 14412 8520
rect 18138 8508 18144 8520
rect 18196 8508 18202 8560
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8480 15623 8483
rect 16482 8480 16488 8492
rect 15611 8452 16488 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 16482 8440 16488 8452
rect 16540 8480 16546 8492
rect 18708 8489 18736 8588
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 19886 8576 19892 8628
rect 19944 8616 19950 8628
rect 20073 8619 20131 8625
rect 20073 8616 20085 8619
rect 19944 8588 20085 8616
rect 19944 8576 19950 8588
rect 20073 8585 20085 8588
rect 20119 8585 20131 8619
rect 20073 8579 20131 8585
rect 21174 8576 21180 8628
rect 21232 8576 21238 8628
rect 21637 8619 21695 8625
rect 21637 8585 21649 8619
rect 21683 8616 21695 8619
rect 22462 8616 22468 8628
rect 21683 8588 22468 8616
rect 21683 8585 21695 8588
rect 21637 8579 21695 8585
rect 22462 8576 22468 8588
rect 22520 8576 22526 8628
rect 23860 8588 24808 8616
rect 21192 8548 21220 8576
rect 23860 8548 23888 8588
rect 21192 8520 23888 8548
rect 24780 8548 24808 8588
rect 25130 8548 25136 8560
rect 24780 8520 25136 8548
rect 25130 8508 25136 8520
rect 25188 8508 25194 8560
rect 18693 8483 18751 8489
rect 18693 8480 18705 8483
rect 16540 8452 18705 8480
rect 16540 8440 16546 8452
rect 18693 8449 18705 8452
rect 18739 8449 18751 8483
rect 22646 8480 22652 8492
rect 18693 8443 18751 8449
rect 22066 8452 22652 8480
rect 15298 8415 15356 8421
rect 15298 8412 15310 8415
rect 14384 8384 15310 8412
rect 15298 8381 15310 8384
rect 15344 8381 15356 8415
rect 15298 8375 15356 8381
rect 17034 8372 17040 8424
rect 17092 8412 17098 8424
rect 17129 8415 17187 8421
rect 17129 8412 17141 8415
rect 17092 8384 17141 8412
rect 17092 8372 17098 8384
rect 17129 8381 17141 8384
rect 17175 8381 17187 8415
rect 17129 8375 17187 8381
rect 17770 8372 17776 8424
rect 17828 8372 17834 8424
rect 17954 8372 17960 8424
rect 18012 8372 18018 8424
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 13725 8347 13783 8353
rect 13725 8313 13737 8347
rect 13771 8344 13783 8347
rect 13814 8344 13820 8356
rect 13771 8316 13820 8344
rect 13771 8313 13783 8316
rect 13725 8307 13783 8313
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 13906 8304 13912 8356
rect 13964 8304 13970 8356
rect 13998 8304 14004 8356
rect 14056 8344 14062 8356
rect 18064 8344 18092 8375
rect 18138 8372 18144 8424
rect 18196 8372 18202 8424
rect 20257 8415 20315 8421
rect 20257 8381 20269 8415
rect 20303 8412 20315 8415
rect 22066 8412 22094 8452
rect 22646 8440 22652 8452
rect 22704 8480 22710 8492
rect 23845 8483 23903 8489
rect 23845 8480 23857 8483
rect 22704 8452 23857 8480
rect 22704 8440 22710 8452
rect 23845 8449 23857 8452
rect 23891 8449 23903 8483
rect 23845 8443 23903 8449
rect 20303 8384 22094 8412
rect 22281 8415 22339 8421
rect 20303 8381 20315 8384
rect 20257 8375 20315 8381
rect 22281 8381 22293 8415
rect 22327 8381 22339 8415
rect 22281 8375 22339 8381
rect 14056 8316 14596 8344
rect 14056 8304 14062 8316
rect 14568 8288 14596 8316
rect 17880 8316 18092 8344
rect 18417 8347 18475 8353
rect 13262 8276 13268 8288
rect 12984 8248 13268 8276
rect 12667 8245 12679 8248
rect 12621 8239 12679 8245
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 13538 8236 13544 8288
rect 13596 8276 13602 8288
rect 14366 8276 14372 8288
rect 13596 8248 14372 8276
rect 13596 8236 13602 8248
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 14550 8236 14556 8288
rect 14608 8276 14614 8288
rect 16758 8276 16764 8288
rect 14608 8248 16764 8276
rect 14608 8236 14614 8248
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 16942 8236 16948 8288
rect 17000 8276 17006 8288
rect 17880 8276 17908 8316
rect 18417 8313 18429 8347
rect 18463 8344 18475 8347
rect 18938 8347 18996 8353
rect 18938 8344 18950 8347
rect 18463 8316 18950 8344
rect 18463 8313 18475 8316
rect 18417 8307 18475 8313
rect 18938 8313 18950 8316
rect 18984 8313 18996 8347
rect 18938 8307 18996 8313
rect 20524 8347 20582 8353
rect 20524 8313 20536 8347
rect 20570 8344 20582 8347
rect 20622 8344 20628 8356
rect 20570 8316 20628 8344
rect 20570 8313 20582 8316
rect 20524 8307 20582 8313
rect 20622 8304 20628 8316
rect 20680 8304 20686 8356
rect 20898 8304 20904 8356
rect 20956 8344 20962 8356
rect 21729 8347 21787 8353
rect 21729 8344 21741 8347
rect 20956 8316 21741 8344
rect 20956 8304 20962 8316
rect 21729 8313 21741 8316
rect 21775 8313 21787 8347
rect 22296 8344 22324 8375
rect 23014 8372 23020 8424
rect 23072 8372 23078 8424
rect 23860 8412 23888 8443
rect 25774 8421 25780 8424
rect 25501 8415 25559 8421
rect 25501 8412 25513 8415
rect 23860 8384 25513 8412
rect 25501 8381 25513 8384
rect 25547 8381 25559 8415
rect 25768 8412 25780 8421
rect 25735 8384 25780 8412
rect 25501 8375 25559 8381
rect 25768 8375 25780 8384
rect 25774 8372 25780 8375
rect 25832 8372 25838 8424
rect 21729 8307 21787 8313
rect 22066 8316 22324 8344
rect 17000 8248 17908 8276
rect 17000 8236 17006 8248
rect 21266 8236 21272 8288
rect 21324 8276 21330 8288
rect 22066 8276 22094 8316
rect 23658 8304 23664 8356
rect 23716 8344 23722 8356
rect 24090 8347 24148 8353
rect 24090 8344 24102 8347
rect 23716 8316 24102 8344
rect 23716 8304 23722 8316
rect 24090 8313 24102 8316
rect 24136 8313 24148 8347
rect 24090 8307 24148 8313
rect 24486 8304 24492 8356
rect 24544 8344 24550 8356
rect 24946 8344 24952 8356
rect 24544 8316 24952 8344
rect 24544 8304 24550 8316
rect 24946 8304 24952 8316
rect 25004 8344 25010 8356
rect 25004 8316 25268 8344
rect 25004 8304 25010 8316
rect 21324 8248 22094 8276
rect 21324 8236 21330 8248
rect 22370 8236 22376 8288
rect 22428 8276 22434 8288
rect 25240 8285 25268 8316
rect 22465 8279 22523 8285
rect 22465 8276 22477 8279
rect 22428 8248 22477 8276
rect 22428 8236 22434 8248
rect 22465 8245 22477 8248
rect 22511 8245 22523 8279
rect 22465 8239 22523 8245
rect 25225 8279 25283 8285
rect 25225 8245 25237 8279
rect 25271 8245 25283 8279
rect 25225 8239 25283 8245
rect 26786 8236 26792 8288
rect 26844 8276 26850 8288
rect 26881 8279 26939 8285
rect 26881 8276 26893 8279
rect 26844 8248 26893 8276
rect 26844 8236 26850 8248
rect 26881 8245 26893 8248
rect 26927 8245 26939 8279
rect 26881 8239 26939 8245
rect 552 8186 27576 8208
rect 552 8134 7114 8186
rect 7166 8134 7178 8186
rect 7230 8134 7242 8186
rect 7294 8134 7306 8186
rect 7358 8134 7370 8186
rect 7422 8134 13830 8186
rect 13882 8134 13894 8186
rect 13946 8134 13958 8186
rect 14010 8134 14022 8186
rect 14074 8134 14086 8186
rect 14138 8134 20546 8186
rect 20598 8134 20610 8186
rect 20662 8134 20674 8186
rect 20726 8134 20738 8186
rect 20790 8134 20802 8186
rect 20854 8134 27262 8186
rect 27314 8134 27326 8186
rect 27378 8134 27390 8186
rect 27442 8134 27454 8186
rect 27506 8134 27518 8186
rect 27570 8134 27576 8186
rect 552 8112 27576 8134
rect 4249 8075 4307 8081
rect 4249 8041 4261 8075
rect 4295 8072 4307 8075
rect 4706 8072 4712 8084
rect 4295 8044 4712 8072
rect 4295 8041 4307 8044
rect 4249 8035 4307 8041
rect 4706 8032 4712 8044
rect 4764 8072 4770 8084
rect 5350 8072 5356 8084
rect 4764 8044 5356 8072
rect 4764 8032 4770 8044
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 5902 8032 5908 8084
rect 5960 8072 5966 8084
rect 6181 8075 6239 8081
rect 6181 8072 6193 8075
rect 5960 8044 6193 8072
rect 5960 8032 5966 8044
rect 6181 8041 6193 8044
rect 6227 8041 6239 8075
rect 6181 8035 6239 8041
rect 6457 8075 6515 8081
rect 6457 8041 6469 8075
rect 6503 8072 6515 8075
rect 6914 8072 6920 8084
rect 6503 8044 6920 8072
rect 6503 8041 6515 8044
rect 6457 8035 6515 8041
rect 6914 8032 6920 8044
rect 6972 8072 6978 8084
rect 7466 8072 7472 8084
rect 6972 8044 7472 8072
rect 6972 8032 6978 8044
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 8570 8032 8576 8084
rect 8628 8072 8634 8084
rect 9582 8072 9588 8084
rect 8628 8044 9588 8072
rect 8628 8032 8634 8044
rect 2216 8007 2274 8013
rect 2216 7973 2228 8007
rect 2262 8004 2274 8007
rect 3513 8007 3571 8013
rect 3513 8004 3525 8007
rect 2262 7976 3525 8004
rect 2262 7973 2274 7976
rect 2216 7967 2274 7973
rect 3513 7973 3525 7976
rect 3559 7973 3571 8007
rect 4154 8004 4160 8016
rect 3513 7967 3571 7973
rect 3896 7976 4160 8004
rect 1486 7896 1492 7948
rect 1544 7936 1550 7948
rect 1946 7936 1952 7948
rect 1544 7908 1952 7936
rect 1544 7896 1550 7908
rect 1946 7896 1952 7908
rect 2004 7896 2010 7948
rect 3418 7896 3424 7948
rect 3476 7896 3482 7948
rect 3896 7945 3924 7976
rect 4154 7964 4160 7976
rect 4212 8004 4218 8016
rect 4401 8007 4459 8013
rect 4401 8004 4413 8007
rect 4212 7976 4413 8004
rect 4212 7964 4218 7976
rect 4401 7973 4413 7976
rect 4447 7973 4459 8007
rect 4401 7967 4459 7973
rect 4617 8007 4675 8013
rect 4617 7973 4629 8007
rect 4663 7973 4675 8007
rect 4617 7967 4675 7973
rect 3605 7939 3663 7945
rect 3605 7905 3617 7939
rect 3651 7936 3663 7939
rect 3881 7939 3939 7945
rect 3651 7908 3740 7936
rect 3651 7905 3663 7908
rect 3605 7899 3663 7905
rect 3712 7809 3740 7908
rect 3881 7905 3893 7939
rect 3927 7905 3939 7939
rect 3881 7899 3939 7905
rect 4062 7896 4068 7948
rect 4120 7896 4126 7948
rect 4632 7936 4660 7967
rect 4801 7939 4859 7945
rect 4801 7936 4813 7939
rect 4632 7908 4813 7936
rect 4801 7905 4813 7908
rect 4847 7936 4859 7939
rect 4890 7936 4896 7948
rect 4847 7908 4896 7936
rect 4847 7905 4859 7908
rect 4801 7899 4859 7905
rect 4890 7896 4896 7908
rect 4948 7936 4954 7948
rect 5920 7936 5948 8032
rect 6086 7964 6092 8016
rect 6144 7964 6150 8016
rect 8294 7964 8300 8016
rect 8352 8004 8358 8016
rect 8941 8007 8999 8013
rect 8941 8004 8953 8007
rect 8352 7976 8953 8004
rect 8352 7964 8358 7976
rect 8941 7973 8953 7976
rect 8987 7973 8999 8007
rect 8941 7967 8999 7973
rect 4948 7908 5948 7936
rect 5997 7939 6055 7945
rect 4948 7896 4954 7908
rect 5997 7905 6009 7939
rect 6043 7905 6055 7939
rect 5997 7899 6055 7905
rect 5074 7828 5080 7880
rect 5132 7868 5138 7880
rect 6012 7868 6040 7899
rect 8846 7896 8852 7948
rect 8904 7896 8910 7948
rect 9048 7936 9076 8044
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 12526 8072 12532 8084
rect 9692 8044 12532 8072
rect 9309 8007 9367 8013
rect 9309 7973 9321 8007
rect 9355 8004 9367 8007
rect 9355 7976 9628 8004
rect 9355 7973 9367 7976
rect 9309 7967 9367 7973
rect 9125 7939 9183 7945
rect 9125 7936 9137 7939
rect 9048 7908 9137 7936
rect 9125 7905 9137 7908
rect 9171 7905 9183 7939
rect 9125 7899 9183 7905
rect 9398 7896 9404 7948
rect 9456 7896 9462 7948
rect 9600 7945 9628 7976
rect 9692 7945 9720 8044
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 16298 8072 16304 8084
rect 12676 8044 13860 8072
rect 12676 8032 12682 8044
rect 10870 8004 10876 8016
rect 10796 7976 10876 8004
rect 10796 7945 10824 7976
rect 10870 7964 10876 7976
rect 10928 8004 10934 8016
rect 11701 8007 11759 8013
rect 11701 8004 11713 8007
rect 10928 7976 11713 8004
rect 10928 7964 10934 7976
rect 11701 7973 11713 7976
rect 11747 7973 11759 8007
rect 11701 7967 11759 7973
rect 13832 8004 13860 8044
rect 14108 8044 16304 8072
rect 14108 8004 14136 8044
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 19153 8075 19211 8081
rect 19153 8072 19165 8075
rect 18196 8044 19165 8072
rect 18196 8032 18202 8044
rect 19153 8041 19165 8044
rect 19199 8041 19211 8075
rect 20346 8072 20352 8084
rect 19153 8035 19211 8041
rect 19306 8044 20352 8072
rect 13832 7976 14136 8004
rect 9585 7939 9643 7945
rect 9585 7905 9597 7939
rect 9631 7905 9643 7939
rect 9585 7899 9643 7905
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 9769 7939 9827 7945
rect 9769 7905 9781 7939
rect 9815 7936 9827 7939
rect 10137 7939 10195 7945
rect 10137 7936 10149 7939
rect 9815 7908 10149 7936
rect 9815 7905 9827 7908
rect 9769 7899 9827 7905
rect 10137 7905 10149 7908
rect 10183 7905 10195 7939
rect 10137 7899 10195 7905
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 5132 7840 6040 7868
rect 6365 7871 6423 7877
rect 5132 7828 5138 7840
rect 6365 7837 6377 7871
rect 6411 7868 6423 7871
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6411 7840 7021 7868
rect 6411 7837 6423 7840
rect 6365 7831 6423 7837
rect 7009 7837 7021 7840
rect 7055 7868 7067 7871
rect 7190 7868 7196 7880
rect 7055 7840 7196 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 9692 7868 9720 7899
rect 11330 7896 11336 7948
rect 11388 7896 11394 7948
rect 11514 7945 11520 7948
rect 11481 7939 11520 7945
rect 11481 7905 11493 7939
rect 11481 7899 11520 7905
rect 11514 7896 11520 7899
rect 11572 7896 11578 7948
rect 11609 7939 11667 7945
rect 11609 7905 11621 7939
rect 11655 7905 11667 7939
rect 11609 7899 11667 7905
rect 11839 7939 11897 7945
rect 11839 7905 11851 7939
rect 11885 7936 11897 7939
rect 12158 7936 12164 7948
rect 11885 7908 12164 7936
rect 11885 7905 11897 7908
rect 11839 7899 11897 7905
rect 8812 7840 9720 7868
rect 11624 7868 11652 7899
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 12342 7945 12348 7948
rect 12336 7899 12348 7945
rect 12342 7896 12348 7899
rect 12400 7896 12406 7948
rect 12710 7896 12716 7948
rect 12768 7936 12774 7948
rect 13722 7945 13728 7948
rect 13541 7939 13599 7945
rect 13541 7936 13553 7939
rect 12768 7908 13553 7936
rect 12768 7896 12774 7908
rect 13541 7905 13553 7908
rect 13587 7905 13599 7939
rect 13541 7899 13599 7905
rect 13689 7939 13728 7945
rect 13689 7905 13701 7939
rect 13689 7899 13728 7905
rect 11698 7868 11704 7880
rect 11624 7840 11704 7868
rect 8812 7828 8818 7840
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7837 12127 7871
rect 13556 7868 13584 7899
rect 13722 7896 13728 7899
rect 13780 7896 13786 7948
rect 13832 7945 13860 7976
rect 14366 7964 14372 8016
rect 14424 8004 14430 8016
rect 14424 7976 16804 8004
rect 14424 7964 14430 7976
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7905 13875 7939
rect 13817 7899 13875 7905
rect 13906 7896 13912 7948
rect 13964 7896 13970 7948
rect 13998 7896 14004 7948
rect 14056 7945 14062 7948
rect 14056 7936 14064 7945
rect 14283 7939 14341 7945
rect 14056 7908 14101 7936
rect 14056 7899 14064 7908
rect 14283 7905 14295 7939
rect 14329 7936 14341 7939
rect 14384 7936 14412 7964
rect 14329 7908 14412 7936
rect 14461 7939 14519 7945
rect 14329 7905 14341 7908
rect 14283 7899 14341 7905
rect 14461 7905 14473 7939
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 14056 7896 14062 7899
rect 14476 7868 14504 7899
rect 14550 7896 14556 7948
rect 14608 7896 14614 7948
rect 14645 7939 14703 7945
rect 14645 7905 14657 7939
rect 14691 7936 14703 7939
rect 16117 7939 16175 7945
rect 16117 7936 16129 7939
rect 14691 7908 16129 7936
rect 14691 7905 14703 7908
rect 14645 7899 14703 7905
rect 16117 7905 16129 7908
rect 16163 7905 16175 7939
rect 16117 7899 16175 7905
rect 13556 7840 13676 7868
rect 12069 7831 12127 7837
rect 3697 7803 3755 7809
rect 3697 7769 3709 7803
rect 3743 7800 3755 7803
rect 5166 7800 5172 7812
rect 3743 7772 5172 7800
rect 3743 7769 3755 7772
rect 3697 7763 3755 7769
rect 5166 7760 5172 7772
rect 5224 7760 5230 7812
rect 11606 7760 11612 7812
rect 11664 7800 11670 7812
rect 12084 7800 12112 7831
rect 11664 7772 12112 7800
rect 11664 7760 11670 7772
rect 3329 7735 3387 7741
rect 3329 7701 3341 7735
rect 3375 7732 3387 7735
rect 4062 7732 4068 7744
rect 3375 7704 4068 7732
rect 3375 7701 3387 7704
rect 3329 7695 3387 7701
rect 4062 7692 4068 7704
rect 4120 7732 4126 7744
rect 4433 7735 4491 7741
rect 4433 7732 4445 7735
rect 4120 7704 4445 7732
rect 4120 7692 4126 7704
rect 4433 7701 4445 7704
rect 4479 7701 4491 7735
rect 4433 7695 4491 7701
rect 5258 7692 5264 7744
rect 5316 7732 5322 7744
rect 5353 7735 5411 7741
rect 5353 7732 5365 7735
rect 5316 7704 5365 7732
rect 5316 7692 5322 7704
rect 5353 7701 5365 7704
rect 5399 7701 5411 7735
rect 5353 7695 5411 7701
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7732 5871 7735
rect 5994 7732 6000 7744
rect 5859 7704 6000 7732
rect 5859 7701 5871 7704
rect 5813 7695 5871 7701
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 10042 7692 10048 7744
rect 10100 7692 10106 7744
rect 11977 7735 12035 7741
rect 11977 7701 11989 7735
rect 12023 7732 12035 7735
rect 12710 7732 12716 7744
rect 12023 7704 12716 7732
rect 12023 7701 12035 7704
rect 11977 7695 12035 7701
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 13449 7735 13507 7741
rect 13449 7701 13461 7735
rect 13495 7732 13507 7735
rect 13538 7732 13544 7744
rect 13495 7704 13544 7732
rect 13495 7701 13507 7704
rect 13449 7695 13507 7701
rect 13538 7692 13544 7704
rect 13596 7692 13602 7744
rect 13648 7732 13676 7840
rect 14200 7840 14504 7868
rect 14921 7871 14979 7877
rect 14200 7809 14228 7840
rect 14921 7837 14933 7871
rect 14967 7868 14979 7871
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 14967 7840 15577 7868
rect 14967 7837 14979 7840
rect 14921 7831 14979 7837
rect 15565 7837 15577 7840
rect 15611 7837 15623 7871
rect 15565 7831 15623 7837
rect 15930 7828 15936 7880
rect 15988 7868 15994 7880
rect 16669 7871 16727 7877
rect 16669 7868 16681 7871
rect 15988 7840 16681 7868
rect 15988 7828 15994 7840
rect 16669 7837 16681 7840
rect 16715 7837 16727 7871
rect 16669 7831 16727 7837
rect 14185 7803 14243 7809
rect 14185 7769 14197 7803
rect 14231 7769 14243 7803
rect 16114 7800 16120 7812
rect 14185 7763 14243 7769
rect 14292 7772 16120 7800
rect 14292 7732 14320 7772
rect 16114 7760 16120 7772
rect 16172 7760 16178 7812
rect 16776 7800 16804 7976
rect 17770 7964 17776 8016
rect 17828 8004 17834 8016
rect 19306 8004 19334 8044
rect 20346 8032 20352 8044
rect 20404 8032 20410 8084
rect 20438 8032 20444 8084
rect 20496 8032 20502 8084
rect 21085 8075 21143 8081
rect 21085 8041 21097 8075
rect 21131 8072 21143 8075
rect 23014 8072 23020 8084
rect 21131 8044 23020 8072
rect 21131 8041 21143 8044
rect 21085 8035 21143 8041
rect 23014 8032 23020 8044
rect 23072 8032 23078 8084
rect 23658 8032 23664 8084
rect 23716 8032 23722 8084
rect 25130 8032 25136 8084
rect 25188 8072 25194 8084
rect 25188 8044 25728 8072
rect 25188 8032 25194 8044
rect 20456 8004 20484 8032
rect 22094 8004 22100 8016
rect 17828 7976 19334 8004
rect 19904 7976 22100 8004
rect 17828 7964 17834 7976
rect 17034 7896 17040 7948
rect 17092 7936 17098 7948
rect 17405 7939 17463 7945
rect 17405 7936 17417 7939
rect 17092 7908 17417 7936
rect 17092 7896 17098 7908
rect 17405 7905 17417 7908
rect 17451 7936 17463 7939
rect 17862 7936 17868 7948
rect 17451 7908 17868 7936
rect 17451 7905 17463 7908
rect 17405 7899 17463 7905
rect 17862 7896 17868 7908
rect 17920 7896 17926 7948
rect 19794 7896 19800 7948
rect 19852 7896 19858 7948
rect 19904 7945 19932 7976
rect 19889 7939 19947 7945
rect 19889 7905 19901 7939
rect 19935 7905 19947 7939
rect 19889 7899 19947 7905
rect 20346 7896 20352 7948
rect 20404 7936 20410 7948
rect 20441 7939 20499 7945
rect 20441 7936 20453 7939
rect 20404 7908 20453 7936
rect 20404 7896 20410 7908
rect 20441 7905 20453 7908
rect 20487 7905 20499 7939
rect 20441 7899 20499 7905
rect 20622 7896 20628 7948
rect 20680 7896 20686 7948
rect 20732 7945 20760 7976
rect 22094 7964 22100 7976
rect 22152 7964 22158 8016
rect 24213 8007 24271 8013
rect 24213 7973 24225 8007
rect 24259 8004 24271 8007
rect 24259 7976 25360 8004
rect 24259 7973 24271 7976
rect 24213 7967 24271 7973
rect 20717 7939 20775 7945
rect 20717 7905 20729 7939
rect 20763 7905 20775 7939
rect 20717 7899 20775 7905
rect 20809 7939 20867 7945
rect 20809 7905 20821 7939
rect 20855 7936 20867 7939
rect 20898 7936 20904 7948
rect 20855 7908 20904 7936
rect 20855 7905 20867 7908
rect 20809 7899 20867 7905
rect 20898 7896 20904 7908
rect 20956 7896 20962 7948
rect 22370 7896 22376 7948
rect 22428 7945 22434 7948
rect 22428 7936 22440 7945
rect 22428 7908 22473 7936
rect 22428 7899 22440 7908
rect 22428 7896 22434 7899
rect 22646 7896 22652 7948
rect 22704 7896 22710 7948
rect 23014 7896 23020 7948
rect 23072 7896 23078 7948
rect 23198 7896 23204 7948
rect 23256 7896 23262 7948
rect 23293 7939 23351 7945
rect 23293 7905 23305 7939
rect 23339 7905 23351 7939
rect 23293 7899 23351 7905
rect 23385 7939 23443 7945
rect 23385 7905 23397 7939
rect 23431 7905 23443 7939
rect 23385 7899 23443 7905
rect 24305 7939 24363 7945
rect 24305 7905 24317 7939
rect 24351 7936 24363 7939
rect 24854 7936 24860 7948
rect 24351 7908 24860 7936
rect 24351 7905 24363 7908
rect 24305 7899 24363 7905
rect 16850 7828 16856 7880
rect 16908 7868 16914 7880
rect 16908 7840 21404 7868
rect 16908 7828 16914 7840
rect 17589 7803 17647 7809
rect 17589 7800 17601 7803
rect 16776 7772 17601 7800
rect 17589 7769 17601 7772
rect 17635 7800 17647 7803
rect 18414 7800 18420 7812
rect 17635 7772 18420 7800
rect 17635 7769 17647 7772
rect 17589 7763 17647 7769
rect 18414 7760 18420 7772
rect 18472 7800 18478 7812
rect 19978 7800 19984 7812
rect 18472 7772 19984 7800
rect 18472 7760 18478 7772
rect 19978 7760 19984 7772
rect 20036 7800 20042 7812
rect 21082 7800 21088 7812
rect 20036 7772 21088 7800
rect 20036 7760 20042 7772
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 21266 7760 21272 7812
rect 21324 7760 21330 7812
rect 13648 7704 14320 7732
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 15013 7735 15071 7741
rect 15013 7732 15025 7735
rect 14884 7704 15025 7732
rect 14884 7692 14890 7704
rect 15013 7701 15025 7704
rect 15059 7701 15071 7735
rect 15013 7695 15071 7701
rect 19058 7692 19064 7744
rect 19116 7732 19122 7744
rect 20073 7735 20131 7741
rect 20073 7732 20085 7735
rect 19116 7704 20085 7732
rect 19116 7692 19122 7704
rect 20073 7701 20085 7704
rect 20119 7701 20131 7735
rect 21376 7732 21404 7840
rect 23308 7800 23336 7899
rect 23400 7868 23428 7899
rect 24854 7896 24860 7908
rect 24912 7896 24918 7948
rect 24946 7896 24952 7948
rect 25004 7896 25010 7948
rect 25332 7945 25360 7976
rect 25317 7939 25375 7945
rect 25317 7905 25329 7939
rect 25363 7905 25375 7939
rect 25317 7899 25375 7905
rect 25590 7896 25596 7948
rect 25648 7896 25654 7948
rect 25700 7936 25728 8044
rect 26605 8007 26663 8013
rect 26605 7973 26617 8007
rect 26651 8004 26663 8007
rect 26970 8004 26976 8016
rect 26651 7976 26976 8004
rect 26651 7973 26663 7976
rect 26605 7967 26663 7973
rect 26970 7964 26976 7976
rect 27028 7964 27034 8016
rect 25869 7939 25927 7945
rect 25869 7936 25881 7939
rect 25700 7908 25881 7936
rect 25869 7905 25881 7908
rect 25915 7905 25927 7939
rect 25869 7899 25927 7905
rect 26786 7896 26792 7948
rect 26844 7896 26850 7948
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 23400 7840 24409 7868
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 25222 7828 25228 7880
rect 25280 7868 25286 7880
rect 25409 7871 25467 7877
rect 25409 7868 25421 7871
rect 25280 7840 25421 7868
rect 25280 7828 25286 7840
rect 25409 7837 25421 7840
rect 25455 7837 25467 7871
rect 25409 7831 25467 7837
rect 26050 7828 26056 7880
rect 26108 7868 26114 7880
rect 26145 7871 26203 7877
rect 26145 7868 26157 7871
rect 26108 7840 26157 7868
rect 26108 7828 26114 7840
rect 26145 7837 26157 7840
rect 26191 7837 26203 7871
rect 26145 7831 26203 7837
rect 24762 7800 24768 7812
rect 23308 7772 24768 7800
rect 24762 7760 24768 7772
rect 24820 7760 24826 7812
rect 25958 7800 25964 7812
rect 25608 7772 25964 7800
rect 22462 7732 22468 7744
rect 21376 7704 22468 7732
rect 20073 7695 20131 7701
rect 22462 7692 22468 7704
rect 22520 7692 22526 7744
rect 25038 7692 25044 7744
rect 25096 7732 25102 7744
rect 25608 7741 25636 7772
rect 25958 7760 25964 7772
rect 26016 7800 26022 7812
rect 26421 7803 26479 7809
rect 26421 7800 26433 7803
rect 26016 7772 26433 7800
rect 26016 7760 26022 7772
rect 26421 7769 26433 7772
rect 26467 7769 26479 7803
rect 26421 7763 26479 7769
rect 25133 7735 25191 7741
rect 25133 7732 25145 7735
rect 25096 7704 25145 7732
rect 25096 7692 25102 7704
rect 25133 7701 25145 7704
rect 25179 7701 25191 7735
rect 25133 7695 25191 7701
rect 25593 7735 25651 7741
rect 25593 7701 25605 7735
rect 25639 7701 25651 7735
rect 25593 7695 25651 7701
rect 25682 7692 25688 7744
rect 25740 7692 25746 7744
rect 25866 7692 25872 7744
rect 25924 7732 25930 7744
rect 26053 7735 26111 7741
rect 26053 7732 26065 7735
rect 25924 7704 26065 7732
rect 25924 7692 25930 7704
rect 26053 7701 26065 7704
rect 26099 7701 26111 7735
rect 26053 7695 26111 7701
rect 552 7642 27416 7664
rect 552 7590 3756 7642
rect 3808 7590 3820 7642
rect 3872 7590 3884 7642
rect 3936 7590 3948 7642
rect 4000 7590 4012 7642
rect 4064 7590 10472 7642
rect 10524 7590 10536 7642
rect 10588 7590 10600 7642
rect 10652 7590 10664 7642
rect 10716 7590 10728 7642
rect 10780 7590 17188 7642
rect 17240 7590 17252 7642
rect 17304 7590 17316 7642
rect 17368 7590 17380 7642
rect 17432 7590 17444 7642
rect 17496 7590 23904 7642
rect 23956 7590 23968 7642
rect 24020 7590 24032 7642
rect 24084 7590 24096 7642
rect 24148 7590 24160 7642
rect 24212 7590 27416 7642
rect 552 7568 27416 7590
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 4580 7500 5089 7528
rect 4580 7488 4586 7500
rect 5077 7497 5089 7500
rect 5123 7497 5135 7531
rect 5077 7491 5135 7497
rect 5166 7488 5172 7540
rect 5224 7488 5230 7540
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 5537 7531 5595 7537
rect 5537 7528 5549 7531
rect 5408 7500 5549 7528
rect 5408 7488 5414 7500
rect 5537 7497 5549 7500
rect 5583 7497 5595 7531
rect 6914 7528 6920 7540
rect 5537 7491 5595 7497
rect 5644 7500 6920 7528
rect 4890 7420 4896 7472
rect 4948 7420 4954 7472
rect 1946 7352 1952 7404
rect 2004 7392 2010 7404
rect 2004 7364 2774 7392
rect 2004 7352 2010 7364
rect 2746 7324 2774 7364
rect 4798 7352 4804 7404
rect 4856 7392 4862 7404
rect 4985 7395 5043 7401
rect 4985 7392 4997 7395
rect 4856 7364 4997 7392
rect 4856 7352 4862 7364
rect 4985 7361 4997 7364
rect 5031 7392 5043 7395
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 5031 7364 5365 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 5353 7361 5365 7364
rect 5399 7392 5411 7395
rect 5534 7392 5540 7404
rect 5399 7364 5540 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 3513 7327 3571 7333
rect 3513 7324 3525 7327
rect 2746 7296 3525 7324
rect 3513 7293 3525 7296
rect 3559 7324 3571 7327
rect 4246 7324 4252 7336
rect 3559 7296 4252 7324
rect 3559 7293 3571 7296
rect 3513 7287 3571 7293
rect 4246 7284 4252 7296
rect 4304 7324 4310 7336
rect 4304 7296 5120 7324
rect 4304 7284 4310 7296
rect 3780 7259 3838 7265
rect 3780 7225 3792 7259
rect 3826 7256 3838 7259
rect 4430 7256 4436 7268
rect 3826 7228 4436 7256
rect 3826 7225 3838 7228
rect 3780 7219 3838 7225
rect 4430 7216 4436 7228
rect 4488 7216 4494 7268
rect 5092 7256 5120 7296
rect 5258 7284 5264 7336
rect 5316 7284 5322 7336
rect 5644 7333 5672 7500
rect 6914 7488 6920 7500
rect 6972 7488 6978 7540
rect 7190 7488 7196 7540
rect 7248 7488 7254 7540
rect 12342 7488 12348 7540
rect 12400 7488 12406 7540
rect 15930 7488 15936 7540
rect 15988 7488 15994 7540
rect 20622 7488 20628 7540
rect 20680 7528 20686 7540
rect 20901 7531 20959 7537
rect 20901 7528 20913 7531
rect 20680 7500 20913 7528
rect 20680 7488 20686 7500
rect 20901 7497 20913 7500
rect 20947 7497 20959 7531
rect 20901 7491 20959 7497
rect 21082 7488 21088 7540
rect 21140 7528 21146 7540
rect 23014 7528 23020 7540
rect 21140 7500 23020 7528
rect 21140 7488 21146 7500
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 23198 7488 23204 7540
rect 23256 7528 23262 7540
rect 23845 7531 23903 7537
rect 23845 7528 23857 7531
rect 23256 7500 23857 7528
rect 23256 7488 23262 7500
rect 23845 7497 23857 7500
rect 23891 7497 23903 7531
rect 23845 7491 23903 7497
rect 24397 7531 24455 7537
rect 24397 7497 24409 7531
rect 24443 7528 24455 7531
rect 25590 7528 25596 7540
rect 24443 7500 25596 7528
rect 24443 7497 24455 7500
rect 24397 7491 24455 7497
rect 25590 7488 25596 7500
rect 25648 7488 25654 7540
rect 26050 7488 26056 7540
rect 26108 7488 26114 7540
rect 11333 7463 11391 7469
rect 8588 7432 9444 7460
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7324 5871 7327
rect 6822 7324 6828 7336
rect 5859 7296 6828 7324
rect 5859 7293 5871 7296
rect 5813 7287 5871 7293
rect 5828 7256 5856 7287
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7324 8539 7327
rect 8588 7324 8616 7432
rect 9416 7404 9444 7432
rect 11333 7429 11345 7463
rect 11379 7460 11391 7463
rect 13906 7460 13912 7472
rect 11379 7432 12020 7460
rect 11379 7429 11391 7432
rect 11333 7423 11391 7429
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 9217 7395 9275 7401
rect 9217 7392 9229 7395
rect 9171 7364 9229 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 9217 7361 9229 7364
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 11992 7401 12020 7432
rect 13188 7432 13912 7460
rect 11977 7395 12035 7401
rect 9456 7364 10088 7392
rect 9456 7352 9462 7364
rect 8527 7296 8616 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 8662 7284 8668 7336
rect 8720 7284 8726 7336
rect 8754 7284 8760 7336
rect 8812 7284 8818 7336
rect 8849 7327 8907 7333
rect 8849 7293 8861 7327
rect 8895 7293 8907 7327
rect 8849 7287 8907 7293
rect 5092 7228 5856 7256
rect 5902 7216 5908 7268
rect 5960 7256 5966 7268
rect 6058 7259 6116 7265
rect 6058 7256 6070 7259
rect 5960 7228 6070 7256
rect 5960 7216 5966 7228
rect 6058 7225 6070 7228
rect 6104 7225 6116 7259
rect 6058 7219 6116 7225
rect 5353 7191 5411 7197
rect 5353 7157 5365 7191
rect 5399 7188 5411 7191
rect 5810 7188 5816 7200
rect 5399 7160 5816 7188
rect 5399 7157 5411 7160
rect 5353 7151 5411 7157
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 8864 7188 8892 7287
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 9953 7327 10011 7333
rect 9953 7324 9965 7327
rect 9732 7296 9965 7324
rect 9732 7284 9738 7296
rect 9953 7293 9965 7296
rect 9999 7293 10011 7327
rect 10060 7324 10088 7364
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 13188 7392 13216 7432
rect 13906 7420 13912 7432
rect 13964 7420 13970 7472
rect 12023 7364 13216 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 13538 7352 13544 7404
rect 13596 7352 13602 7404
rect 15948 7392 15976 7488
rect 16669 7463 16727 7469
rect 16669 7429 16681 7463
rect 16715 7460 16727 7463
rect 18690 7460 18696 7472
rect 16715 7432 18696 7460
rect 16715 7429 16727 7432
rect 16669 7423 16727 7429
rect 18690 7420 18696 7432
rect 18748 7420 18754 7472
rect 20073 7463 20131 7469
rect 20073 7429 20085 7463
rect 20119 7460 20131 7463
rect 20119 7432 20760 7460
rect 20119 7429 20131 7432
rect 20073 7423 20131 7429
rect 16850 7392 16856 7404
rect 15948 7364 16160 7392
rect 10060 7296 10364 7324
rect 9953 7287 10011 7293
rect 9861 7259 9919 7265
rect 9861 7225 9873 7259
rect 9907 7256 9919 7259
rect 10198 7259 10256 7265
rect 10198 7256 10210 7259
rect 9907 7228 10210 7256
rect 9907 7225 9919 7228
rect 9861 7219 9919 7225
rect 10198 7225 10210 7228
rect 10244 7225 10256 7259
rect 10336 7256 10364 7296
rect 11698 7284 11704 7336
rect 11756 7324 11762 7336
rect 12250 7324 12256 7336
rect 11756 7296 12256 7324
rect 11756 7284 11762 7296
rect 12250 7284 12256 7296
rect 12308 7324 12314 7336
rect 12618 7324 12624 7336
rect 12308 7296 12624 7324
rect 12308 7284 12314 7296
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 12802 7284 12808 7336
rect 12860 7324 12866 7336
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 12860 7296 12909 7324
rect 12860 7284 12866 7296
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 13081 7327 13139 7333
rect 13081 7293 13093 7327
rect 13127 7324 13139 7327
rect 13170 7324 13176 7336
rect 13127 7296 13176 7324
rect 13127 7293 13139 7296
rect 13081 7287 13139 7293
rect 13170 7284 13176 7296
rect 13228 7284 13234 7336
rect 13556 7296 14504 7324
rect 13556 7256 13584 7296
rect 10336 7228 13584 7256
rect 10198 7219 10256 7225
rect 13630 7216 13636 7268
rect 13688 7256 13694 7268
rect 14185 7259 14243 7265
rect 14185 7256 14197 7259
rect 13688 7228 14197 7256
rect 13688 7216 13694 7228
rect 14185 7225 14197 7228
rect 14231 7225 14243 7259
rect 14185 7219 14243 7225
rect 11425 7191 11483 7197
rect 11425 7188 11437 7191
rect 8864 7160 11437 7188
rect 11425 7157 11437 7160
rect 11471 7157 11483 7191
rect 11425 7151 11483 7157
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 13170 7188 13176 7200
rect 12676 7160 13176 7188
rect 12676 7148 12682 7160
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13265 7191 13323 7197
rect 13265 7157 13277 7191
rect 13311 7188 13323 7191
rect 14366 7188 14372 7200
rect 13311 7160 14372 7188
rect 13311 7157 13323 7160
rect 13265 7151 13323 7157
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 14476 7188 14504 7296
rect 14550 7284 14556 7336
rect 14608 7284 14614 7336
rect 14826 7333 14832 7336
rect 14820 7324 14832 7333
rect 14787 7296 14832 7324
rect 14820 7287 14832 7296
rect 14826 7284 14832 7287
rect 14884 7284 14890 7336
rect 16022 7284 16028 7336
rect 16080 7284 16086 7336
rect 16132 7333 16160 7364
rect 16546 7364 16856 7392
rect 16546 7333 16574 7364
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 20732 7401 20760 7432
rect 20990 7420 20996 7472
rect 21048 7460 21054 7472
rect 21048 7432 21312 7460
rect 21048 7420 21054 7432
rect 20717 7395 20775 7401
rect 18064 7364 18819 7392
rect 16118 7327 16176 7333
rect 16118 7293 16130 7327
rect 16164 7293 16176 7327
rect 16118 7287 16176 7293
rect 16531 7327 16589 7333
rect 16531 7293 16543 7327
rect 16577 7293 16589 7327
rect 16531 7287 16589 7293
rect 16761 7327 16819 7333
rect 16761 7293 16773 7327
rect 16807 7324 16819 7327
rect 17034 7324 17040 7336
rect 16807 7296 17040 7324
rect 16807 7293 16819 7296
rect 16761 7287 16819 7293
rect 17034 7284 17040 7296
rect 17092 7284 17098 7336
rect 17586 7284 17592 7336
rect 17644 7324 17650 7336
rect 17681 7327 17739 7333
rect 17681 7324 17693 7327
rect 17644 7296 17693 7324
rect 17644 7284 17650 7296
rect 17681 7293 17693 7296
rect 17727 7293 17739 7327
rect 17681 7287 17739 7293
rect 17865 7327 17923 7333
rect 17865 7293 17877 7327
rect 17911 7293 17923 7327
rect 17865 7287 17923 7293
rect 16298 7216 16304 7268
rect 16356 7216 16362 7268
rect 16390 7216 16396 7268
rect 16448 7216 16454 7268
rect 16850 7216 16856 7268
rect 16908 7256 16914 7268
rect 17880 7256 17908 7287
rect 17954 7284 17960 7336
rect 18012 7284 18018 7336
rect 18064 7333 18092 7364
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 18693 7327 18751 7333
rect 18693 7293 18705 7327
rect 18739 7293 18751 7327
rect 18791 7324 18819 7364
rect 20717 7361 20729 7395
rect 20763 7392 20775 7395
rect 20763 7364 21220 7392
rect 20763 7361 20775 7364
rect 20717 7355 20775 7361
rect 21192 7333 21220 7364
rect 21284 7333 21312 7432
rect 22462 7420 22468 7472
rect 22520 7420 22526 7472
rect 25866 7420 25872 7472
rect 25924 7420 25930 7472
rect 24762 7392 24768 7404
rect 24044 7364 24768 7392
rect 20165 7327 20223 7333
rect 20165 7324 20177 7327
rect 18791 7296 20177 7324
rect 18693 7287 18751 7293
rect 20165 7293 20177 7296
rect 20211 7293 20223 7327
rect 20165 7287 20223 7293
rect 21080 7327 21138 7333
rect 21080 7293 21092 7327
rect 21126 7293 21138 7327
rect 21080 7287 21138 7293
rect 21177 7327 21235 7333
rect 21177 7293 21189 7327
rect 21223 7293 21235 7327
rect 21177 7287 21235 7293
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7293 21327 7327
rect 21269 7287 21327 7293
rect 21452 7327 21510 7333
rect 21452 7293 21464 7327
rect 21498 7293 21510 7327
rect 21452 7287 21510 7293
rect 18708 7256 18736 7287
rect 16908 7228 17908 7256
rect 17972 7228 18736 7256
rect 18960 7259 19018 7265
rect 16908 7216 16914 7228
rect 17972 7200 18000 7228
rect 18960 7225 18972 7259
rect 19006 7256 19018 7259
rect 19334 7256 19340 7268
rect 19006 7228 19340 7256
rect 19006 7225 19018 7228
rect 18960 7219 19018 7225
rect 19334 7216 19340 7228
rect 19392 7216 19398 7268
rect 15562 7188 15568 7200
rect 14476 7160 15568 7188
rect 15562 7148 15568 7160
rect 15620 7188 15626 7200
rect 16945 7191 17003 7197
rect 16945 7188 16957 7191
rect 15620 7160 16957 7188
rect 15620 7148 15626 7160
rect 16945 7157 16957 7160
rect 16991 7188 17003 7191
rect 17586 7188 17592 7200
rect 16991 7160 17592 7188
rect 16991 7157 17003 7160
rect 16945 7151 17003 7157
rect 17586 7148 17592 7160
rect 17644 7188 17650 7200
rect 17770 7188 17776 7200
rect 17644 7160 17776 7188
rect 17644 7148 17650 7160
rect 17770 7148 17776 7160
rect 17828 7148 17834 7200
rect 17954 7148 17960 7200
rect 18012 7148 18018 7200
rect 18325 7191 18383 7197
rect 18325 7157 18337 7191
rect 18371 7188 18383 7191
rect 19886 7188 19892 7200
rect 18371 7160 19892 7188
rect 18371 7157 18383 7160
rect 18325 7151 18383 7157
rect 19886 7148 19892 7160
rect 19944 7148 19950 7200
rect 21100 7188 21128 7287
rect 21467 7256 21495 7287
rect 21542 7284 21548 7336
rect 21600 7284 21606 7336
rect 21634 7284 21640 7336
rect 21692 7284 21698 7336
rect 24044 7333 24072 7364
rect 24762 7352 24768 7364
rect 24820 7352 24826 7404
rect 25884 7392 25912 7420
rect 24964 7364 25912 7392
rect 22649 7327 22707 7333
rect 22649 7293 22661 7327
rect 22695 7293 22707 7327
rect 22649 7287 22707 7293
rect 24026 7327 24084 7333
rect 24026 7293 24038 7327
rect 24072 7293 24084 7327
rect 24026 7287 24084 7293
rect 24489 7327 24547 7333
rect 24489 7293 24501 7327
rect 24535 7324 24547 7327
rect 24578 7324 24584 7336
rect 24535 7296 24584 7324
rect 24535 7293 24547 7296
rect 24489 7287 24547 7293
rect 22281 7259 22339 7265
rect 22281 7256 22293 7259
rect 21467 7228 22293 7256
rect 22281 7225 22293 7228
rect 22327 7256 22339 7259
rect 22370 7256 22376 7268
rect 22327 7228 22376 7256
rect 22327 7225 22339 7228
rect 22281 7219 22339 7225
rect 22370 7216 22376 7228
rect 22428 7216 22434 7268
rect 22664 7188 22692 7287
rect 24578 7284 24584 7296
rect 24636 7284 24642 7336
rect 24964 7333 24992 7364
rect 24857 7327 24915 7333
rect 24857 7293 24869 7327
rect 24903 7293 24915 7327
rect 24857 7287 24915 7293
rect 24949 7327 25007 7333
rect 24949 7293 24961 7327
rect 24995 7293 25007 7327
rect 24949 7287 25007 7293
rect 24872 7256 24900 7287
rect 25038 7284 25044 7336
rect 25096 7284 25102 7336
rect 25130 7284 25136 7336
rect 25188 7324 25194 7336
rect 25225 7327 25283 7333
rect 25225 7324 25237 7327
rect 25188 7296 25237 7324
rect 25188 7284 25194 7296
rect 25225 7293 25237 7296
rect 25271 7293 25283 7327
rect 25225 7287 25283 7293
rect 25866 7284 25872 7336
rect 25924 7284 25930 7336
rect 26602 7284 26608 7336
rect 26660 7284 26666 7336
rect 25317 7259 25375 7265
rect 25317 7256 25329 7259
rect 24872 7228 25329 7256
rect 25317 7225 25329 7228
rect 25363 7225 25375 7259
rect 25317 7219 25375 7225
rect 23014 7188 23020 7200
rect 21100 7160 23020 7188
rect 23014 7148 23020 7160
rect 23072 7148 23078 7200
rect 24029 7191 24087 7197
rect 24029 7157 24041 7191
rect 24075 7188 24087 7191
rect 24302 7188 24308 7200
rect 24075 7160 24308 7188
rect 24075 7157 24087 7160
rect 24029 7151 24087 7157
rect 24302 7148 24308 7160
rect 24360 7148 24366 7200
rect 24578 7148 24584 7200
rect 24636 7148 24642 7200
rect 552 7098 27576 7120
rect 552 7046 7114 7098
rect 7166 7046 7178 7098
rect 7230 7046 7242 7098
rect 7294 7046 7306 7098
rect 7358 7046 7370 7098
rect 7422 7046 13830 7098
rect 13882 7046 13894 7098
rect 13946 7046 13958 7098
rect 14010 7046 14022 7098
rect 14074 7046 14086 7098
rect 14138 7046 20546 7098
rect 20598 7046 20610 7098
rect 20662 7046 20674 7098
rect 20726 7046 20738 7098
rect 20790 7046 20802 7098
rect 20854 7046 27262 7098
rect 27314 7046 27326 7098
rect 27378 7046 27390 7098
rect 27442 7046 27454 7098
rect 27506 7046 27518 7098
rect 27570 7046 27576 7098
rect 552 7024 27576 7046
rect 5626 6944 5632 6996
rect 5684 6944 5690 6996
rect 5902 6944 5908 6996
rect 5960 6944 5966 6996
rect 8662 6944 8668 6996
rect 8720 6944 8726 6996
rect 8846 6944 8852 6996
rect 8904 6944 8910 6996
rect 9674 6944 9680 6996
rect 9732 6944 9738 6996
rect 10781 6987 10839 6993
rect 10781 6953 10793 6987
rect 10827 6984 10839 6987
rect 10870 6984 10876 6996
rect 10827 6956 10876 6984
rect 10827 6953 10839 6956
rect 10781 6947 10839 6953
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 15286 6984 15292 6996
rect 12584 6956 15292 6984
rect 12584 6944 12590 6956
rect 15286 6944 15292 6956
rect 15344 6944 15350 6996
rect 15933 6987 15991 6993
rect 15933 6953 15945 6987
rect 15979 6984 15991 6987
rect 16390 6984 16396 6996
rect 15979 6956 16396 6984
rect 15979 6953 15991 6956
rect 15933 6947 15991 6953
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 21269 6987 21327 6993
rect 21269 6953 21281 6987
rect 21315 6984 21327 6987
rect 21634 6984 21640 6996
rect 21315 6956 21640 6984
rect 21315 6953 21327 6956
rect 21269 6947 21327 6953
rect 21634 6944 21640 6956
rect 21692 6944 21698 6996
rect 24854 6944 24860 6996
rect 24912 6984 24918 6996
rect 25685 6987 25743 6993
rect 25685 6984 25697 6987
rect 24912 6956 25697 6984
rect 24912 6944 24918 6956
rect 25685 6953 25697 6956
rect 25731 6984 25743 6987
rect 25866 6984 25872 6996
rect 25731 6956 25872 6984
rect 25731 6953 25743 6956
rect 25685 6947 25743 6953
rect 25866 6944 25872 6956
rect 25924 6944 25930 6996
rect 26237 6987 26295 6993
rect 26237 6953 26249 6987
rect 26283 6984 26295 6987
rect 26602 6984 26608 6996
rect 26283 6956 26608 6984
rect 26283 6953 26295 6956
rect 26237 6947 26295 6953
rect 26602 6944 26608 6956
rect 26660 6944 26666 6996
rect 5644 6916 5672 6944
rect 7926 6916 7932 6928
rect 5644 6888 7932 6916
rect 7926 6876 7932 6888
rect 7984 6876 7990 6928
rect 8864 6916 8892 6944
rect 9692 6916 9720 6944
rect 13630 6916 13636 6928
rect 8864 6888 9168 6916
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6848 5503 6851
rect 5534 6848 5540 6860
rect 5491 6820 5540 6848
rect 5491 6817 5503 6820
rect 5445 6811 5503 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6817 5687 6851
rect 5629 6811 5687 6817
rect 5644 6780 5672 6811
rect 5810 6808 5816 6860
rect 5868 6808 5874 6860
rect 5994 6808 6000 6860
rect 6052 6808 6058 6860
rect 8110 6808 8116 6860
rect 8168 6808 8174 6860
rect 8570 6808 8576 6860
rect 8628 6848 8634 6860
rect 8849 6851 8907 6857
rect 8849 6848 8861 6851
rect 8628 6820 8861 6848
rect 8628 6808 8634 6820
rect 8849 6817 8861 6820
rect 8895 6817 8907 6851
rect 8849 6811 8907 6817
rect 9030 6808 9036 6860
rect 9088 6808 9094 6860
rect 9140 6857 9168 6888
rect 9600 6888 9720 6916
rect 12544 6888 13636 6916
rect 9125 6851 9183 6857
rect 9125 6817 9137 6851
rect 9171 6817 9183 6851
rect 9125 6811 9183 6817
rect 9401 6851 9459 6857
rect 9401 6817 9413 6851
rect 9447 6848 9459 6851
rect 9600 6848 9628 6888
rect 9447 6820 9628 6848
rect 9668 6851 9726 6857
rect 9447 6817 9459 6820
rect 9401 6811 9459 6817
rect 9668 6817 9680 6851
rect 9714 6848 9726 6851
rect 10042 6848 10048 6860
rect 9714 6820 10048 6848
rect 9714 6817 9726 6820
rect 9668 6811 9726 6817
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 11882 6808 11888 6860
rect 11940 6808 11946 6860
rect 11974 6808 11980 6860
rect 12032 6808 12038 6860
rect 12158 6808 12164 6860
rect 12216 6808 12222 6860
rect 12544 6857 12572 6888
rect 13630 6876 13636 6888
rect 13688 6876 13694 6928
rect 14752 6888 14964 6916
rect 12529 6851 12587 6857
rect 12529 6817 12541 6851
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 12618 6808 12624 6860
rect 12676 6808 12682 6860
rect 12710 6808 12716 6860
rect 12768 6808 12774 6860
rect 12894 6808 12900 6860
rect 12952 6808 12958 6860
rect 12986 6808 12992 6860
rect 13044 6848 13050 6860
rect 13725 6851 13783 6857
rect 13725 6848 13737 6851
rect 13044 6820 13737 6848
rect 13044 6808 13050 6820
rect 13725 6817 13737 6820
rect 13771 6817 13783 6851
rect 13725 6811 13783 6817
rect 13817 6851 13875 6857
rect 13817 6817 13829 6851
rect 13863 6817 13875 6851
rect 13817 6811 13875 6817
rect 14001 6851 14059 6857
rect 14001 6817 14013 6851
rect 14047 6848 14059 6851
rect 14090 6848 14096 6860
rect 14047 6820 14096 6848
rect 14047 6817 14059 6820
rect 14001 6811 14059 6817
rect 7098 6780 7104 6792
rect 5644 6752 7104 6780
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 11238 6740 11244 6792
rect 11296 6780 11302 6792
rect 11701 6783 11759 6789
rect 11701 6780 11713 6783
rect 11296 6752 11713 6780
rect 11296 6740 11302 6752
rect 11701 6749 11713 6752
rect 11747 6749 11759 6783
rect 11701 6743 11759 6749
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6780 12311 6783
rect 12802 6780 12808 6792
rect 12299 6752 12808 6780
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 13538 6740 13544 6792
rect 13596 6780 13602 6792
rect 13832 6780 13860 6811
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 14185 6851 14243 6857
rect 14185 6817 14197 6851
rect 14231 6848 14243 6851
rect 14752 6848 14780 6888
rect 14826 6857 14832 6860
rect 14231 6820 14780 6848
rect 14231 6817 14243 6820
rect 14185 6811 14243 6817
rect 14820 6811 14832 6857
rect 14826 6808 14832 6811
rect 14884 6808 14890 6860
rect 14936 6848 14964 6888
rect 16408 6848 16436 6944
rect 24578 6925 24584 6928
rect 24572 6916 24584 6925
rect 17788 6888 18092 6916
rect 24539 6888 24584 6916
rect 17788 6857 17816 6888
rect 16669 6851 16727 6857
rect 16669 6848 16681 6851
rect 14936 6820 16068 6848
rect 16408 6820 16681 6848
rect 13596 6752 13860 6780
rect 13596 6740 13602 6752
rect 14550 6740 14556 6792
rect 14608 6740 14614 6792
rect 16040 6780 16068 6820
rect 16669 6817 16681 6820
rect 16715 6817 16727 6851
rect 16669 6811 16727 6817
rect 17773 6851 17831 6857
rect 17773 6817 17785 6851
rect 17819 6817 17831 6851
rect 17773 6811 17831 6817
rect 17865 6851 17923 6857
rect 17865 6817 17877 6851
rect 17911 6848 17923 6851
rect 17954 6848 17960 6860
rect 17911 6820 17960 6848
rect 17911 6817 17923 6820
rect 17865 6811 17923 6817
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 18064 6848 18092 6888
rect 24572 6879 24584 6888
rect 24578 6876 24584 6879
rect 24636 6876 24642 6928
rect 18121 6851 18179 6857
rect 18121 6848 18133 6851
rect 18064 6820 18133 6848
rect 18121 6817 18133 6820
rect 18167 6817 18179 6851
rect 18121 6811 18179 6817
rect 19334 6808 19340 6860
rect 19392 6808 19398 6860
rect 19886 6808 19892 6860
rect 19944 6808 19950 6860
rect 19996 6820 20944 6848
rect 16850 6780 16856 6792
rect 16040 6752 16856 6780
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6780 17279 6783
rect 17678 6780 17684 6792
rect 17267 6752 17684 6780
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 19150 6740 19156 6792
rect 19208 6780 19214 6792
rect 19996 6780 20024 6820
rect 19208 6752 20024 6780
rect 20717 6783 20775 6789
rect 19208 6740 19214 6752
rect 20717 6749 20729 6783
rect 20763 6749 20775 6783
rect 20717 6743 20775 6749
rect 12161 6715 12219 6721
rect 12161 6681 12173 6715
rect 12207 6712 12219 6715
rect 12434 6712 12440 6724
rect 12207 6684 12440 6712
rect 12207 6681 12219 6684
rect 12161 6675 12219 6681
rect 12434 6672 12440 6684
rect 12492 6672 12498 6724
rect 19168 6712 19196 6740
rect 18791 6684 19196 6712
rect 19245 6715 19303 6721
rect 5350 6604 5356 6656
rect 5408 6644 5414 6656
rect 5445 6647 5503 6653
rect 5445 6644 5457 6647
rect 5408 6616 5457 6644
rect 5408 6604 5414 6616
rect 5445 6613 5457 6616
rect 5491 6613 5503 6647
rect 5445 6607 5503 6613
rect 6822 6604 6828 6656
rect 6880 6604 6886 6656
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 11149 6647 11207 6653
rect 11149 6644 11161 6647
rect 11020 6616 11161 6644
rect 11020 6604 11026 6616
rect 11149 6613 11161 6616
rect 11195 6613 11207 6647
rect 11149 6607 11207 6613
rect 12250 6604 12256 6656
rect 12308 6644 12314 6656
rect 12989 6647 13047 6653
rect 12989 6644 13001 6647
rect 12308 6616 13001 6644
rect 12308 6604 12314 6616
rect 12989 6613 13001 6616
rect 13035 6613 13047 6647
rect 12989 6607 13047 6613
rect 15194 6604 15200 6656
rect 15252 6644 15258 6656
rect 16117 6647 16175 6653
rect 16117 6644 16129 6647
rect 15252 6616 16129 6644
rect 15252 6604 15258 6616
rect 16117 6613 16129 6616
rect 16163 6613 16175 6647
rect 16117 6607 16175 6613
rect 16298 6604 16304 6656
rect 16356 6644 16362 6656
rect 18791 6644 18819 6684
rect 19245 6681 19257 6715
rect 19291 6712 19303 6715
rect 20732 6712 20760 6743
rect 20916 6721 20944 6820
rect 20990 6808 20996 6860
rect 21048 6848 21054 6860
rect 21085 6851 21143 6857
rect 21085 6848 21097 6851
rect 21048 6820 21097 6848
rect 21048 6808 21054 6820
rect 21085 6817 21097 6820
rect 21131 6848 21143 6851
rect 21450 6848 21456 6860
rect 21131 6820 21456 6848
rect 21131 6817 21143 6820
rect 21085 6811 21143 6817
rect 21450 6808 21456 6820
rect 21508 6808 21514 6860
rect 22393 6851 22451 6857
rect 22393 6817 22405 6851
rect 22439 6848 22451 6851
rect 22741 6851 22799 6857
rect 22741 6848 22753 6851
rect 22439 6820 22753 6848
rect 22439 6817 22451 6820
rect 22393 6811 22451 6817
rect 22741 6817 22753 6820
rect 22787 6817 22799 6851
rect 22741 6811 22799 6817
rect 25590 6808 25596 6860
rect 25648 6848 25654 6860
rect 25869 6851 25927 6857
rect 25869 6848 25881 6851
rect 25648 6820 25881 6848
rect 25648 6808 25654 6820
rect 25869 6817 25881 6820
rect 25915 6817 25927 6851
rect 25869 6811 25927 6817
rect 26053 6851 26111 6857
rect 26053 6817 26065 6851
rect 26099 6848 26111 6851
rect 26421 6851 26479 6857
rect 26421 6848 26433 6851
rect 26099 6820 26433 6848
rect 26099 6817 26111 6820
rect 26053 6811 26111 6817
rect 26421 6817 26433 6820
rect 26467 6817 26479 6851
rect 26421 6811 26479 6817
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 19291 6684 20760 6712
rect 20901 6715 20959 6721
rect 19291 6681 19303 6684
rect 19245 6675 19303 6681
rect 20901 6681 20913 6715
rect 20947 6681 20959 6715
rect 20901 6675 20959 6681
rect 22664 6712 22692 6743
rect 23290 6740 23296 6792
rect 23348 6740 23354 6792
rect 24302 6780 24308 6792
rect 23952 6752 24308 6780
rect 23952 6712 23980 6752
rect 24302 6740 24308 6752
rect 24360 6740 24366 6792
rect 25777 6783 25835 6789
rect 25777 6749 25789 6783
rect 25823 6780 25835 6783
rect 26786 6780 26792 6792
rect 25823 6752 26792 6780
rect 25823 6749 25835 6752
rect 25777 6743 25835 6749
rect 26786 6740 26792 6752
rect 26844 6740 26850 6792
rect 26970 6740 26976 6792
rect 27028 6740 27034 6792
rect 22664 6684 23980 6712
rect 16356 6616 18819 6644
rect 16356 6604 16362 6616
rect 18966 6604 18972 6656
rect 19024 6644 19030 6656
rect 20073 6647 20131 6653
rect 20073 6644 20085 6647
rect 19024 6616 20085 6644
rect 19024 6604 19030 6616
rect 20073 6613 20085 6616
rect 20119 6613 20131 6647
rect 20073 6607 20131 6613
rect 21726 6604 21732 6656
rect 21784 6644 21790 6656
rect 22664 6644 22692 6684
rect 21784 6616 22692 6644
rect 21784 6604 21790 6616
rect 552 6554 27416 6576
rect 552 6502 3756 6554
rect 3808 6502 3820 6554
rect 3872 6502 3884 6554
rect 3936 6502 3948 6554
rect 4000 6502 4012 6554
rect 4064 6502 10472 6554
rect 10524 6502 10536 6554
rect 10588 6502 10600 6554
rect 10652 6502 10664 6554
rect 10716 6502 10728 6554
rect 10780 6502 17188 6554
rect 17240 6502 17252 6554
rect 17304 6502 17316 6554
rect 17368 6502 17380 6554
rect 17432 6502 17444 6554
rect 17496 6502 23904 6554
rect 23956 6502 23968 6554
rect 24020 6502 24032 6554
rect 24084 6502 24096 6554
rect 24148 6502 24160 6554
rect 24212 6502 27416 6554
rect 552 6480 27416 6502
rect 5534 6400 5540 6452
rect 5592 6400 5598 6452
rect 6086 6400 6092 6452
rect 6144 6440 6150 6452
rect 6457 6443 6515 6449
rect 6457 6440 6469 6443
rect 6144 6412 6469 6440
rect 6144 6400 6150 6412
rect 6457 6409 6469 6412
rect 6503 6409 6515 6443
rect 6457 6403 6515 6409
rect 6638 6400 6644 6452
rect 6696 6400 6702 6452
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 7558 6440 7564 6452
rect 7156 6412 7564 6440
rect 7156 6400 7162 6412
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 13354 6440 13360 6452
rect 7984 6412 13360 6440
rect 7984 6400 7990 6412
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 14826 6400 14832 6452
rect 14884 6440 14890 6452
rect 14921 6443 14979 6449
rect 14921 6440 14933 6443
rect 14884 6412 14933 6440
rect 14884 6400 14890 6412
rect 14921 6409 14933 6412
rect 14967 6409 14979 6443
rect 14921 6403 14979 6409
rect 17678 6400 17684 6452
rect 17736 6440 17742 6452
rect 18693 6443 18751 6449
rect 18693 6440 18705 6443
rect 17736 6412 18705 6440
rect 17736 6400 17742 6412
rect 18693 6409 18705 6412
rect 18739 6409 18751 6443
rect 21266 6440 21272 6452
rect 18693 6403 18751 6409
rect 19306 6412 21272 6440
rect 5445 6375 5503 6381
rect 5445 6341 5457 6375
rect 5491 6372 5503 6375
rect 5994 6372 6000 6384
rect 5491 6344 6000 6372
rect 5491 6341 5503 6344
rect 5445 6335 5503 6341
rect 5994 6332 6000 6344
rect 6052 6372 6058 6384
rect 6052 6344 6132 6372
rect 6052 6332 6058 6344
rect 5626 6264 5632 6316
rect 5684 6264 5690 6316
rect 6104 6313 6132 6344
rect 6270 6332 6276 6384
rect 6328 6372 6334 6384
rect 7009 6375 7067 6381
rect 7009 6372 7021 6375
rect 6328 6344 7021 6372
rect 6328 6332 6334 6344
rect 7009 6341 7021 6344
rect 7055 6341 7067 6375
rect 7009 6335 7067 6341
rect 11974 6332 11980 6384
rect 12032 6372 12038 6384
rect 12345 6375 12403 6381
rect 12345 6372 12357 6375
rect 12032 6344 12357 6372
rect 12032 6332 12038 6344
rect 12345 6341 12357 6344
rect 12391 6341 12403 6375
rect 12345 6335 12403 6341
rect 17586 6332 17592 6384
rect 17644 6372 17650 6384
rect 19306 6372 19334 6412
rect 21266 6400 21272 6412
rect 21324 6440 21330 6452
rect 22465 6443 22523 6449
rect 21324 6412 21864 6440
rect 21324 6400 21330 6412
rect 17644 6344 19334 6372
rect 17644 6332 17650 6344
rect 6089 6307 6147 6313
rect 6089 6273 6101 6307
rect 6135 6304 6147 6307
rect 8294 6304 8300 6316
rect 6135 6276 7328 6304
rect 6135 6273 6147 6276
rect 6089 6267 6147 6273
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6205 4767 6239
rect 4709 6199 4767 6205
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6236 5319 6239
rect 5353 6239 5411 6245
rect 5353 6236 5365 6239
rect 5307 6208 5365 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 5353 6205 5365 6208
rect 5399 6205 5411 6239
rect 5353 6199 5411 6205
rect 4246 6128 4252 6180
rect 4304 6168 4310 6180
rect 4724 6168 4752 6199
rect 5902 6196 5908 6248
rect 5960 6196 5966 6248
rect 5997 6239 6055 6245
rect 5997 6205 6009 6239
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 6181 6239 6239 6245
rect 6181 6205 6193 6239
rect 6227 6236 6239 6239
rect 6914 6236 6920 6248
rect 6227 6208 6920 6236
rect 6227 6205 6239 6208
rect 6181 6199 6239 6205
rect 6012 6168 6040 6199
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 7300 6245 7328 6276
rect 7484 6276 8300 6304
rect 7484 6245 7512 6276
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 8846 6264 8852 6316
rect 8904 6304 8910 6316
rect 11790 6304 11796 6316
rect 8904 6276 11796 6304
rect 8904 6264 8910 6276
rect 11790 6264 11796 6276
rect 11848 6264 11854 6316
rect 12250 6304 12256 6316
rect 12084 6276 12256 6304
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6205 7527 6239
rect 7469 6199 7527 6205
rect 6641 6171 6699 6177
rect 4304 6140 6224 6168
rect 4304 6128 4310 6140
rect 6196 6112 6224 6140
rect 6641 6137 6653 6171
rect 6687 6137 6699 6171
rect 6641 6131 6699 6137
rect 6178 6060 6184 6112
rect 6236 6060 6242 6112
rect 6365 6103 6423 6109
rect 6365 6069 6377 6103
rect 6411 6100 6423 6103
rect 6656 6100 6684 6131
rect 6730 6128 6736 6180
rect 6788 6168 6794 6180
rect 7484 6168 7512 6199
rect 7558 6196 7564 6248
rect 7616 6196 7622 6248
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6236 7803 6239
rect 7791 6208 8064 6236
rect 7791 6205 7803 6208
rect 7745 6199 7803 6205
rect 6788 6140 7512 6168
rect 7576 6168 7604 6196
rect 8036 6177 8064 6208
rect 8662 6196 8668 6248
rect 8720 6196 8726 6248
rect 9401 6239 9459 6245
rect 9401 6205 9413 6239
rect 9447 6236 9459 6239
rect 9493 6239 9551 6245
rect 9493 6236 9505 6239
rect 9447 6208 9505 6236
rect 9447 6205 9459 6208
rect 9401 6199 9459 6205
rect 9493 6205 9505 6208
rect 9539 6205 9551 6239
rect 9493 6199 9551 6205
rect 9858 6196 9864 6248
rect 9916 6196 9922 6248
rect 11514 6196 11520 6248
rect 11572 6236 11578 6248
rect 11882 6236 11888 6248
rect 11572 6208 11888 6236
rect 11572 6196 11578 6208
rect 11882 6196 11888 6208
rect 11940 6196 11946 6248
rect 11974 6196 11980 6248
rect 12032 6196 12038 6248
rect 12084 6245 12112 6276
rect 12250 6264 12256 6276
rect 12308 6264 12314 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12406 6276 12909 6304
rect 12406 6248 12434 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 17034 6264 17040 6316
rect 17092 6304 17098 6316
rect 17092 6276 18276 6304
rect 17092 6264 17098 6276
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6205 12127 6239
rect 12069 6199 12127 6205
rect 12161 6239 12219 6245
rect 12161 6205 12173 6239
rect 12207 6236 12219 6239
rect 12207 6208 12296 6236
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 7837 6171 7895 6177
rect 7837 6168 7849 6171
rect 7576 6140 7849 6168
rect 6788 6128 6794 6140
rect 7837 6137 7849 6140
rect 7883 6137 7895 6171
rect 7837 6131 7895 6137
rect 8021 6171 8079 6177
rect 8021 6137 8033 6171
rect 8067 6168 8079 6171
rect 9030 6168 9036 6180
rect 8067 6140 9036 6168
rect 8067 6137 8079 6140
rect 8021 6131 8079 6137
rect 9030 6128 9036 6140
rect 9088 6128 9094 6180
rect 11330 6128 11336 6180
rect 11388 6168 11394 6180
rect 12084 6168 12112 6199
rect 12268 6180 12296 6208
rect 12342 6196 12348 6248
rect 12400 6208 12434 6248
rect 12400 6196 12406 6208
rect 14366 6196 14372 6248
rect 14424 6196 14430 6248
rect 14642 6196 14648 6248
rect 14700 6196 14706 6248
rect 14918 6196 14924 6248
rect 14976 6236 14982 6248
rect 15473 6239 15531 6245
rect 15473 6236 15485 6239
rect 14976 6208 15485 6236
rect 14976 6196 14982 6208
rect 15473 6205 15485 6208
rect 15519 6205 15531 6239
rect 15473 6199 15531 6205
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6236 15807 6239
rect 16574 6236 16580 6248
rect 15795 6208 16580 6236
rect 15795 6205 15807 6208
rect 15749 6199 15807 6205
rect 11388 6140 12112 6168
rect 11388 6128 11394 6140
rect 12250 6128 12256 6180
rect 12308 6128 12314 6180
rect 14461 6171 14519 6177
rect 14461 6168 14473 6171
rect 12406 6140 14473 6168
rect 6411 6072 6684 6100
rect 6411 6069 6423 6072
rect 6365 6063 6423 6069
rect 7742 6060 7748 6112
rect 7800 6060 7806 6112
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6100 8263 6103
rect 8386 6100 8392 6112
rect 8251 6072 8392 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 8481 6103 8539 6109
rect 8481 6069 8493 6103
rect 8527 6100 8539 6103
rect 8570 6100 8576 6112
rect 8527 6072 8576 6100
rect 8527 6069 8539 6072
rect 8481 6063 8539 6069
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 9582 6060 9588 6112
rect 9640 6060 9646 6112
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 9732 6072 11161 6100
rect 9732 6060 9738 6072
rect 11149 6069 11161 6072
rect 11195 6100 11207 6103
rect 11606 6100 11612 6112
rect 11195 6072 11612 6100
rect 11195 6069 11207 6072
rect 11149 6063 11207 6069
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 11698 6060 11704 6112
rect 11756 6060 11762 6112
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 12406 6100 12434 6140
rect 14461 6137 14473 6140
rect 14507 6137 14519 6171
rect 14461 6131 14519 6137
rect 14550 6128 14556 6180
rect 14608 6168 14614 6180
rect 15764 6168 15792 6199
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 18248 6245 18276 6276
rect 18690 6264 18696 6316
rect 18748 6304 18754 6316
rect 20993 6307 21051 6313
rect 18748 6276 19196 6304
rect 18748 6264 18754 6276
rect 17865 6239 17923 6245
rect 17865 6236 17877 6239
rect 17144 6208 17877 6236
rect 14608 6140 15792 6168
rect 16016 6171 16074 6177
rect 14608 6128 14614 6140
rect 16016 6137 16028 6171
rect 16062 6168 16074 6171
rect 16114 6168 16120 6180
rect 16062 6140 16120 6168
rect 16062 6137 16074 6140
rect 16016 6131 16074 6137
rect 16114 6128 16120 6140
rect 16172 6128 16178 6180
rect 11848 6072 12434 6100
rect 14829 6103 14887 6109
rect 11848 6060 11854 6072
rect 14829 6069 14841 6103
rect 14875 6100 14887 6103
rect 15378 6100 15384 6112
rect 14875 6072 15384 6100
rect 14875 6069 14887 6072
rect 14829 6063 14887 6069
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 17144 6109 17172 6208
rect 17865 6205 17877 6208
rect 17911 6236 17923 6239
rect 18233 6239 18291 6245
rect 17911 6208 18092 6236
rect 17911 6205 17923 6208
rect 17865 6199 17923 6205
rect 18064 6168 18092 6208
rect 18233 6205 18245 6239
rect 18279 6205 18291 6239
rect 18233 6199 18291 6205
rect 18966 6196 18972 6248
rect 19024 6196 19030 6248
rect 19058 6196 19064 6248
rect 19116 6196 19122 6248
rect 19168 6245 19196 6276
rect 20993 6273 21005 6307
rect 21039 6304 21051 6307
rect 21726 6304 21732 6316
rect 21039 6276 21732 6304
rect 21039 6273 21051 6276
rect 20993 6267 21051 6273
rect 21726 6264 21732 6276
rect 21784 6264 21790 6316
rect 19153 6239 19211 6245
rect 19153 6205 19165 6239
rect 19199 6205 19211 6239
rect 19153 6199 19211 6205
rect 19337 6239 19395 6245
rect 19337 6205 19349 6239
rect 19383 6205 19395 6239
rect 19337 6199 19395 6205
rect 19242 6168 19248 6180
rect 18064 6140 19248 6168
rect 19242 6128 19248 6140
rect 19300 6128 19306 6180
rect 19352 6112 19380 6199
rect 21634 6196 21640 6248
rect 21692 6196 21698 6248
rect 21836 6245 21864 6412
rect 22465 6409 22477 6443
rect 22511 6440 22523 6443
rect 23290 6440 23296 6452
rect 22511 6412 23296 6440
rect 22511 6409 22523 6412
rect 22465 6403 22523 6409
rect 23290 6400 23296 6412
rect 23348 6400 23354 6452
rect 25961 6443 26019 6449
rect 25961 6409 25973 6443
rect 26007 6440 26019 6443
rect 26970 6440 26976 6452
rect 26007 6412 26976 6440
rect 26007 6409 26019 6412
rect 25961 6403 26019 6409
rect 26970 6400 26976 6412
rect 27028 6400 27034 6452
rect 21910 6332 21916 6384
rect 21968 6332 21974 6384
rect 22094 6332 22100 6384
rect 22152 6372 22158 6384
rect 22152 6344 23612 6372
rect 22152 6332 22158 6344
rect 21821 6239 21879 6245
rect 21821 6205 21833 6239
rect 21867 6205 21879 6239
rect 21928 6236 21956 6332
rect 22370 6264 22376 6316
rect 22428 6264 22434 6316
rect 21984 6239 22042 6245
rect 21984 6236 21996 6239
rect 21928 6208 21996 6236
rect 21821 6199 21879 6205
rect 21984 6205 21996 6208
rect 22030 6205 22042 6239
rect 21984 6199 22042 6205
rect 22094 6196 22100 6248
rect 22152 6236 22158 6248
rect 22235 6239 22293 6245
rect 22152 6208 22197 6236
rect 22152 6196 22158 6208
rect 22235 6205 22247 6239
rect 22281 6236 22293 6239
rect 22388 6236 22416 6264
rect 23584 6245 23612 6344
rect 24302 6264 24308 6316
rect 24360 6304 24366 6316
rect 24581 6307 24639 6313
rect 24581 6304 24593 6307
rect 24360 6276 24593 6304
rect 24360 6264 24366 6276
rect 24581 6273 24593 6276
rect 24627 6273 24639 6307
rect 24581 6267 24639 6273
rect 22281 6208 22416 6236
rect 22833 6239 22891 6245
rect 22281 6205 22293 6208
rect 22235 6199 22293 6205
rect 22833 6205 22845 6239
rect 22879 6205 22891 6239
rect 22833 6199 22891 6205
rect 23569 6239 23627 6245
rect 23569 6205 23581 6239
rect 23615 6205 23627 6239
rect 23569 6199 23627 6205
rect 20748 6171 20806 6177
rect 20748 6137 20760 6171
rect 20794 6168 20806 6171
rect 21085 6171 21143 6177
rect 21085 6168 21097 6171
rect 20794 6140 21097 6168
rect 20794 6137 20806 6140
rect 20748 6131 20806 6137
rect 21085 6137 21097 6140
rect 21131 6137 21143 6171
rect 21085 6131 21143 6137
rect 22370 6128 22376 6180
rect 22428 6168 22434 6180
rect 22848 6168 22876 6199
rect 24394 6196 24400 6248
rect 24452 6196 24458 6248
rect 24848 6239 24906 6245
rect 24848 6205 24860 6239
rect 24894 6236 24906 6239
rect 25682 6236 25688 6248
rect 24894 6208 25688 6236
rect 24894 6205 24906 6208
rect 24848 6199 24906 6205
rect 25682 6196 25688 6208
rect 25740 6196 25746 6248
rect 22428 6140 22876 6168
rect 22428 6128 22434 6140
rect 17129 6103 17187 6109
rect 17129 6069 17141 6103
rect 17175 6069 17187 6103
rect 17129 6063 17187 6069
rect 17218 6060 17224 6112
rect 17276 6060 17282 6112
rect 18417 6103 18475 6109
rect 18417 6069 18429 6103
rect 18463 6100 18475 6103
rect 19334 6100 19340 6112
rect 18463 6072 19340 6100
rect 18463 6069 18475 6072
rect 18417 6063 18475 6069
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 19613 6103 19671 6109
rect 19613 6069 19625 6103
rect 19659 6100 19671 6103
rect 20346 6100 20352 6112
rect 19659 6072 20352 6100
rect 19659 6069 19671 6072
rect 19613 6063 19671 6069
rect 20346 6060 20352 6072
rect 20404 6060 20410 6112
rect 20438 6060 20444 6112
rect 20496 6100 20502 6112
rect 22186 6100 22192 6112
rect 20496 6072 22192 6100
rect 20496 6060 20502 6072
rect 22186 6060 22192 6072
rect 22244 6100 22250 6112
rect 22649 6103 22707 6109
rect 22649 6100 22661 6103
rect 22244 6072 22661 6100
rect 22244 6060 22250 6072
rect 22649 6069 22661 6072
rect 22695 6069 22707 6103
rect 22649 6063 22707 6069
rect 23198 6060 23204 6112
rect 23256 6100 23262 6112
rect 23385 6103 23443 6109
rect 23385 6100 23397 6103
rect 23256 6072 23397 6100
rect 23256 6060 23262 6072
rect 23385 6069 23397 6072
rect 23431 6069 23443 6103
rect 23385 6063 23443 6069
rect 23474 6060 23480 6112
rect 23532 6100 23538 6112
rect 23845 6103 23903 6109
rect 23845 6100 23857 6103
rect 23532 6072 23857 6100
rect 23532 6060 23538 6072
rect 23845 6069 23857 6072
rect 23891 6069 23903 6103
rect 23845 6063 23903 6069
rect 552 6010 27576 6032
rect 552 5958 7114 6010
rect 7166 5958 7178 6010
rect 7230 5958 7242 6010
rect 7294 5958 7306 6010
rect 7358 5958 7370 6010
rect 7422 5958 13830 6010
rect 13882 5958 13894 6010
rect 13946 5958 13958 6010
rect 14010 5958 14022 6010
rect 14074 5958 14086 6010
rect 14138 5958 20546 6010
rect 20598 5958 20610 6010
rect 20662 5958 20674 6010
rect 20726 5958 20738 6010
rect 20790 5958 20802 6010
rect 20854 5958 27262 6010
rect 27314 5958 27326 6010
rect 27378 5958 27390 6010
rect 27442 5958 27454 6010
rect 27506 5958 27518 6010
rect 27570 5958 27576 6010
rect 552 5936 27576 5958
rect 4246 5856 4252 5908
rect 4304 5856 4310 5908
rect 5994 5856 6000 5908
rect 6052 5896 6058 5908
rect 6365 5899 6423 5905
rect 6365 5896 6377 5899
rect 6052 5868 6377 5896
rect 6052 5856 6058 5868
rect 6365 5865 6377 5868
rect 6411 5865 6423 5899
rect 6365 5859 6423 5865
rect 6457 5899 6515 5905
rect 6457 5865 6469 5899
rect 6503 5896 6515 5899
rect 6730 5896 6736 5908
rect 6503 5868 6736 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 6178 5788 6184 5840
rect 6236 5828 6242 5840
rect 6472 5828 6500 5859
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 8205 5899 8263 5905
rect 8205 5865 8217 5899
rect 8251 5896 8263 5899
rect 8846 5896 8852 5908
rect 8251 5868 8852 5896
rect 8251 5865 8263 5868
rect 8205 5859 8263 5865
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 10134 5856 10140 5908
rect 10192 5856 10198 5908
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 13081 5899 13139 5905
rect 13081 5896 13093 5899
rect 12032 5868 13093 5896
rect 12032 5856 12038 5868
rect 13081 5865 13093 5868
rect 13127 5865 13139 5899
rect 13081 5859 13139 5865
rect 13354 5856 13360 5908
rect 13412 5896 13418 5908
rect 13412 5868 14228 5896
rect 13412 5856 13418 5868
rect 6914 5828 6920 5840
rect 6236 5800 6500 5828
rect 6564 5800 6920 5828
rect 6236 5788 6242 5800
rect 5350 5720 5356 5772
rect 5408 5769 5414 5772
rect 5408 5760 5420 5769
rect 5997 5763 6055 5769
rect 5408 5732 5453 5760
rect 5408 5723 5420 5732
rect 5997 5729 6009 5763
rect 6043 5760 6055 5763
rect 6086 5760 6092 5772
rect 6043 5732 6092 5760
rect 6043 5729 6055 5732
rect 5997 5723 6055 5729
rect 5408 5720 5414 5723
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 6273 5763 6331 5769
rect 6273 5729 6285 5763
rect 6319 5760 6331 5763
rect 6564 5760 6592 5800
rect 6914 5788 6920 5800
rect 6972 5828 6978 5840
rect 8018 5828 8024 5840
rect 6972 5800 8024 5828
rect 6972 5788 6978 5800
rect 8018 5788 8024 5800
rect 8076 5788 8082 5840
rect 9674 5828 9680 5840
rect 8312 5800 9680 5828
rect 6319 5732 6592 5760
rect 7092 5763 7150 5769
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 7092 5729 7104 5763
rect 7138 5760 7150 5763
rect 7374 5760 7380 5772
rect 7138 5732 7380 5760
rect 7138 5729 7150 5732
rect 7092 5723 7150 5729
rect 7374 5720 7380 5732
rect 7432 5720 7438 5772
rect 8312 5769 8340 5800
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 11698 5828 11704 5840
rect 11164 5800 11704 5828
rect 8570 5769 8576 5772
rect 8297 5763 8355 5769
rect 8297 5729 8309 5763
rect 8343 5729 8355 5763
rect 8564 5760 8576 5769
rect 8531 5732 8576 5760
rect 8297 5723 8355 5729
rect 8564 5723 8576 5732
rect 8570 5720 8576 5723
rect 8628 5720 8634 5772
rect 8938 5720 8944 5772
rect 8996 5760 9002 5772
rect 9861 5763 9919 5769
rect 9861 5760 9873 5763
rect 8996 5732 9873 5760
rect 8996 5720 9002 5732
rect 9861 5729 9873 5732
rect 9907 5729 9919 5763
rect 9861 5723 9919 5729
rect 5629 5695 5687 5701
rect 5629 5661 5641 5695
rect 5675 5692 5687 5695
rect 6822 5692 6828 5704
rect 5675 5664 6828 5692
rect 5675 5661 5687 5664
rect 5629 5655 5687 5661
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 6638 5584 6644 5636
rect 6696 5584 6702 5636
rect 9876 5624 9904 5723
rect 10962 5720 10968 5772
rect 11020 5720 11026 5772
rect 11164 5769 11192 5800
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 12066 5788 12072 5840
rect 12124 5788 12130 5840
rect 12158 5788 12164 5840
rect 12216 5828 12222 5840
rect 14093 5831 14151 5837
rect 14093 5828 14105 5831
rect 12216 5800 14105 5828
rect 12216 5788 12222 5800
rect 14093 5797 14105 5800
rect 14139 5797 14151 5831
rect 14093 5791 14151 5797
rect 11149 5763 11207 5769
rect 11149 5729 11161 5763
rect 11195 5729 11207 5763
rect 11149 5723 11207 5729
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5760 11299 5763
rect 11330 5760 11336 5772
rect 11287 5732 11336 5760
rect 11287 5729 11299 5732
rect 11241 5723 11299 5729
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 11422 5720 11428 5772
rect 11480 5720 11486 5772
rect 11514 5720 11520 5772
rect 11572 5720 11578 5772
rect 11606 5720 11612 5772
rect 11664 5720 11670 5772
rect 11865 5763 11923 5769
rect 11865 5760 11877 5763
rect 11716 5732 11877 5760
rect 11057 5695 11115 5701
rect 11057 5661 11069 5695
rect 11103 5692 11115 5695
rect 11716 5692 11744 5732
rect 11865 5729 11877 5732
rect 11911 5729 11923 5763
rect 12084 5760 12112 5788
rect 13817 5763 13875 5769
rect 13817 5760 13829 5763
rect 12084 5732 13829 5760
rect 11865 5723 11923 5729
rect 13817 5729 13829 5732
rect 13863 5729 13875 5763
rect 13817 5723 13875 5729
rect 11103 5664 11744 5692
rect 11103 5661 11115 5664
rect 11057 5655 11115 5661
rect 13630 5652 13636 5704
rect 13688 5652 13694 5704
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5692 14151 5695
rect 14200 5692 14228 5868
rect 14918 5856 14924 5908
rect 14976 5856 14982 5908
rect 16114 5856 16120 5908
rect 16172 5856 16178 5908
rect 17218 5856 17224 5908
rect 17276 5856 17282 5908
rect 19702 5856 19708 5908
rect 19760 5896 19766 5908
rect 20438 5896 20444 5908
rect 19760 5868 20444 5896
rect 19760 5856 19766 5868
rect 20438 5856 20444 5868
rect 20496 5856 20502 5908
rect 21542 5896 21548 5908
rect 21284 5868 21548 5896
rect 16942 5828 16948 5840
rect 15304 5800 16948 5828
rect 15304 5772 15332 5800
rect 16942 5788 16948 5800
rect 17000 5828 17006 5840
rect 17236 5828 17264 5856
rect 19613 5831 19671 5837
rect 19613 5828 19625 5831
rect 17000 5800 17080 5828
rect 17000 5788 17006 5800
rect 14366 5720 14372 5772
rect 14424 5720 14430 5772
rect 14458 5720 14464 5772
rect 14516 5720 14522 5772
rect 14642 5720 14648 5772
rect 14700 5720 14706 5772
rect 15194 5720 15200 5772
rect 15252 5720 15258 5772
rect 15286 5720 15292 5772
rect 15344 5720 15350 5772
rect 15378 5720 15384 5772
rect 15436 5720 15442 5772
rect 15562 5720 15568 5772
rect 15620 5720 15626 5772
rect 14139 5664 14228 5692
rect 16761 5695 16819 5701
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 16761 5661 16773 5695
rect 16807 5692 16819 5695
rect 16853 5695 16911 5701
rect 16853 5692 16865 5695
rect 16807 5664 16865 5692
rect 16807 5661 16819 5664
rect 16761 5655 16819 5661
rect 16853 5661 16865 5664
rect 16899 5661 16911 5695
rect 17052 5692 17080 5800
rect 17144 5800 17264 5828
rect 18248 5800 19625 5828
rect 17144 5769 17172 5800
rect 17129 5763 17187 5769
rect 17129 5729 17141 5763
rect 17175 5729 17187 5763
rect 17129 5723 17187 5729
rect 17221 5763 17279 5769
rect 17221 5729 17233 5763
rect 17267 5729 17279 5763
rect 17221 5723 17279 5729
rect 17313 5763 17371 5769
rect 17313 5729 17325 5763
rect 17359 5729 17371 5763
rect 17313 5723 17371 5729
rect 17236 5692 17264 5723
rect 17052 5664 17264 5692
rect 16853 5655 16911 5661
rect 9876 5596 11192 5624
rect 5810 5516 5816 5568
rect 5868 5516 5874 5568
rect 6089 5559 6147 5565
rect 6089 5525 6101 5559
rect 6135 5556 6147 5559
rect 6270 5556 6276 5568
rect 6135 5528 6276 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 6730 5516 6736 5568
rect 6788 5556 6794 5568
rect 8938 5556 8944 5568
rect 6788 5528 8944 5556
rect 6788 5516 6794 5528
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 9030 5516 9036 5568
rect 9088 5556 9094 5568
rect 9677 5559 9735 5565
rect 9677 5556 9689 5559
rect 9088 5528 9689 5556
rect 9088 5516 9094 5528
rect 9677 5525 9689 5528
rect 9723 5525 9735 5559
rect 11164 5556 11192 5596
rect 11238 5584 11244 5636
rect 11296 5584 11302 5636
rect 13909 5627 13967 5633
rect 13909 5624 13921 5627
rect 12912 5596 13921 5624
rect 11330 5556 11336 5568
rect 11164 5528 11336 5556
rect 9677 5519 9735 5525
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 11514 5516 11520 5568
rect 11572 5556 11578 5568
rect 12912 5556 12940 5596
rect 13909 5593 13921 5596
rect 13955 5593 13967 5627
rect 13909 5587 13967 5593
rect 14829 5627 14887 5633
rect 14829 5593 14841 5627
rect 14875 5624 14887 5627
rect 17328 5624 17356 5723
rect 17494 5720 17500 5772
rect 17552 5720 17558 5772
rect 17586 5720 17592 5772
rect 17644 5760 17650 5772
rect 17865 5763 17923 5769
rect 17865 5760 17877 5763
rect 17644 5732 17877 5760
rect 17644 5720 17650 5732
rect 17865 5729 17877 5732
rect 17911 5729 17923 5763
rect 17865 5723 17923 5729
rect 18046 5720 18052 5772
rect 18104 5720 18110 5772
rect 18138 5720 18144 5772
rect 18196 5720 18202 5772
rect 18248 5769 18276 5800
rect 19613 5797 19625 5800
rect 19659 5797 19671 5831
rect 20898 5828 20904 5840
rect 19613 5791 19671 5797
rect 20272 5800 20904 5828
rect 18233 5763 18291 5769
rect 18233 5729 18245 5763
rect 18279 5729 18291 5763
rect 18233 5723 18291 5729
rect 18877 5763 18935 5769
rect 18877 5729 18889 5763
rect 18923 5729 18935 5763
rect 18877 5723 18935 5729
rect 18892 5692 18920 5723
rect 18966 5720 18972 5772
rect 19024 5760 19030 5772
rect 19024 5732 19069 5760
rect 19024 5720 19030 5732
rect 19150 5720 19156 5772
rect 19208 5720 19214 5772
rect 19242 5720 19248 5772
rect 19300 5720 19306 5772
rect 19383 5763 19441 5769
rect 19383 5729 19395 5763
rect 19429 5760 19441 5763
rect 20272 5760 20300 5800
rect 20898 5788 20904 5800
rect 20956 5788 20962 5840
rect 19429 5732 20300 5760
rect 19429 5729 19441 5732
rect 19383 5723 19441 5729
rect 20346 5720 20352 5772
rect 20404 5720 20410 5772
rect 21284 5769 21312 5868
rect 21542 5856 21548 5868
rect 21600 5856 21606 5908
rect 21910 5856 21916 5908
rect 21968 5856 21974 5908
rect 23385 5899 23443 5905
rect 23385 5896 23397 5899
rect 22112 5868 23397 5896
rect 22112 5828 22140 5868
rect 23385 5865 23397 5868
rect 23431 5896 23443 5899
rect 24394 5896 24400 5908
rect 23431 5868 24400 5896
rect 23431 5865 23443 5868
rect 23385 5859 23443 5865
rect 24394 5856 24400 5868
rect 24452 5856 24458 5908
rect 23750 5828 23756 5840
rect 21432 5800 22140 5828
rect 22572 5800 23756 5828
rect 21432 5769 21460 5800
rect 21269 5763 21327 5769
rect 21269 5729 21281 5763
rect 21315 5729 21327 5763
rect 21269 5723 21327 5729
rect 21417 5763 21475 5769
rect 21417 5729 21429 5763
rect 21463 5729 21475 5763
rect 21417 5723 21475 5729
rect 21542 5720 21548 5772
rect 21600 5720 21606 5772
rect 21818 5769 21824 5772
rect 21637 5763 21695 5769
rect 21637 5729 21649 5763
rect 21683 5729 21695 5763
rect 21637 5723 21695 5729
rect 21775 5763 21824 5769
rect 21775 5729 21787 5763
rect 21821 5729 21824 5763
rect 21775 5723 21824 5729
rect 19702 5692 19708 5704
rect 18892 5664 19708 5692
rect 19702 5652 19708 5664
rect 19760 5652 19766 5704
rect 20070 5652 20076 5704
rect 20128 5692 20134 5704
rect 20165 5695 20223 5701
rect 20165 5692 20177 5695
rect 20128 5664 20177 5692
rect 20128 5652 20134 5664
rect 20165 5661 20177 5664
rect 20211 5692 20223 5695
rect 21652 5692 21680 5723
rect 21818 5720 21824 5723
rect 21876 5720 21882 5772
rect 21993 5763 22051 5769
rect 21993 5760 22005 5763
rect 21928 5732 22005 5760
rect 20211 5664 21680 5692
rect 20211 5661 20223 5664
rect 20165 5655 20223 5661
rect 14875 5596 17356 5624
rect 19521 5627 19579 5633
rect 14875 5593 14887 5596
rect 14829 5587 14887 5593
rect 19521 5593 19533 5627
rect 19567 5624 19579 5627
rect 20254 5624 20260 5636
rect 19567 5596 20260 5624
rect 19567 5593 19579 5596
rect 19521 5587 19579 5593
rect 20254 5584 20260 5596
rect 20312 5584 20318 5636
rect 20364 5596 21128 5624
rect 11572 5528 12940 5556
rect 12989 5559 13047 5565
rect 11572 5516 11578 5528
rect 12989 5525 13001 5559
rect 13035 5556 13047 5559
rect 13538 5556 13544 5568
rect 13035 5528 13544 5556
rect 13035 5525 13047 5528
rect 12989 5519 13047 5525
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 18509 5559 18567 5565
rect 18509 5525 18521 5559
rect 18555 5556 18567 5559
rect 18966 5556 18972 5568
rect 18555 5528 18972 5556
rect 18555 5525 18567 5528
rect 18509 5519 18567 5525
rect 18966 5516 18972 5528
rect 19024 5516 19030 5568
rect 19978 5516 19984 5568
rect 20036 5556 20042 5568
rect 20364 5556 20392 5596
rect 20036 5528 20392 5556
rect 20036 5516 20042 5528
rect 20990 5516 20996 5568
rect 21048 5516 21054 5568
rect 21100 5556 21128 5596
rect 21542 5584 21548 5636
rect 21600 5624 21606 5636
rect 21928 5624 21956 5732
rect 21993 5729 22005 5732
rect 22039 5729 22051 5763
rect 21993 5723 22051 5729
rect 22370 5720 22376 5772
rect 22428 5720 22434 5772
rect 22572 5769 22600 5800
rect 23750 5788 23756 5800
rect 23808 5788 23814 5840
rect 24302 5788 24308 5840
rect 24360 5828 24366 5840
rect 24670 5828 24676 5840
rect 24360 5800 24676 5828
rect 24360 5788 24366 5800
rect 24670 5788 24676 5800
rect 24728 5828 24734 5840
rect 24728 5800 24808 5828
rect 24728 5788 24734 5800
rect 22521 5763 22600 5769
rect 22521 5729 22533 5763
rect 22567 5732 22600 5763
rect 22567 5729 22579 5732
rect 22521 5723 22579 5729
rect 22646 5720 22652 5772
rect 22704 5720 22710 5772
rect 22738 5720 22744 5772
rect 22796 5720 22802 5772
rect 22879 5763 22937 5769
rect 22879 5729 22891 5763
rect 22925 5760 22937 5763
rect 23014 5760 23020 5772
rect 22925 5732 23020 5760
rect 22925 5729 22937 5732
rect 22879 5723 22937 5729
rect 22094 5652 22100 5704
rect 22152 5692 22158 5704
rect 22904 5692 22932 5723
rect 23014 5720 23020 5732
rect 23072 5720 23078 5772
rect 24780 5769 24808 5800
rect 24509 5763 24567 5769
rect 24509 5729 24521 5763
rect 24555 5760 24567 5763
rect 24765 5763 24823 5769
rect 24555 5732 24716 5760
rect 24555 5729 24567 5732
rect 24509 5723 24567 5729
rect 22152 5664 22932 5692
rect 24688 5692 24716 5732
rect 24765 5729 24777 5763
rect 24811 5729 24823 5763
rect 24765 5723 24823 5729
rect 24857 5695 24915 5701
rect 24857 5692 24869 5695
rect 24688 5664 24869 5692
rect 22152 5652 22158 5664
rect 24857 5661 24869 5664
rect 24903 5661 24915 5695
rect 24857 5655 24915 5661
rect 25406 5652 25412 5704
rect 25464 5652 25470 5704
rect 22738 5624 22744 5636
rect 21600 5596 21956 5624
rect 22112 5596 22744 5624
rect 21600 5584 21606 5596
rect 22112 5556 22140 5596
rect 22738 5584 22744 5596
rect 22796 5584 22802 5636
rect 21100 5528 22140 5556
rect 22189 5559 22247 5565
rect 22189 5525 22201 5559
rect 22235 5556 22247 5559
rect 22646 5556 22652 5568
rect 22235 5528 22652 5556
rect 22235 5525 22247 5528
rect 22189 5519 22247 5525
rect 22646 5516 22652 5528
rect 22704 5516 22710 5568
rect 23017 5559 23075 5565
rect 23017 5525 23029 5559
rect 23063 5556 23075 5559
rect 23106 5556 23112 5568
rect 23063 5528 23112 5556
rect 23063 5525 23075 5528
rect 23017 5519 23075 5525
rect 23106 5516 23112 5528
rect 23164 5516 23170 5568
rect 552 5466 27416 5488
rect 552 5414 3756 5466
rect 3808 5414 3820 5466
rect 3872 5414 3884 5466
rect 3936 5414 3948 5466
rect 4000 5414 4012 5466
rect 4064 5414 10472 5466
rect 10524 5414 10536 5466
rect 10588 5414 10600 5466
rect 10652 5414 10664 5466
rect 10716 5414 10728 5466
rect 10780 5414 17188 5466
rect 17240 5414 17252 5466
rect 17304 5414 17316 5466
rect 17368 5414 17380 5466
rect 17432 5414 17444 5466
rect 17496 5414 23904 5466
rect 23956 5414 23968 5466
rect 24020 5414 24032 5466
rect 24084 5414 24096 5466
rect 24148 5414 24160 5466
rect 24212 5414 27416 5466
rect 552 5392 27416 5414
rect 5902 5312 5908 5364
rect 5960 5352 5966 5364
rect 5997 5355 6055 5361
rect 5997 5352 6009 5355
rect 5960 5324 6009 5352
rect 5960 5312 5966 5324
rect 5997 5321 6009 5324
rect 6043 5352 6055 5355
rect 6638 5352 6644 5364
rect 6043 5324 6644 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 7374 5312 7380 5364
rect 7432 5312 7438 5364
rect 8386 5312 8392 5364
rect 8444 5352 8450 5364
rect 8573 5355 8631 5361
rect 8573 5352 8585 5355
rect 8444 5324 8585 5352
rect 8444 5312 8450 5324
rect 8573 5321 8585 5324
rect 8619 5321 8631 5355
rect 8573 5315 8631 5321
rect 8662 5312 8668 5364
rect 8720 5352 8726 5364
rect 8757 5355 8815 5361
rect 8757 5352 8769 5355
rect 8720 5324 8769 5352
rect 8720 5312 8726 5324
rect 8757 5321 8769 5324
rect 8803 5321 8815 5355
rect 8757 5315 8815 5321
rect 11333 5355 11391 5361
rect 11333 5321 11345 5355
rect 11379 5352 11391 5355
rect 11422 5352 11428 5364
rect 11379 5324 11428 5352
rect 11379 5321 11391 5324
rect 11333 5315 11391 5321
rect 11422 5312 11428 5324
rect 11480 5352 11486 5364
rect 12342 5352 12348 5364
rect 11480 5324 12348 5352
rect 11480 5312 11486 5324
rect 12342 5312 12348 5324
rect 12400 5352 12406 5364
rect 13630 5352 13636 5364
rect 12400 5324 13636 5352
rect 12400 5312 12406 5324
rect 6362 5244 6368 5296
rect 6420 5284 6426 5296
rect 6420 5256 11008 5284
rect 6420 5244 6426 5256
rect 8846 5176 8852 5228
rect 8904 5216 8910 5228
rect 9217 5219 9275 5225
rect 9217 5216 9229 5219
rect 8904 5188 9229 5216
rect 8904 5176 8910 5188
rect 9217 5185 9229 5188
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 4614 5108 4620 5160
rect 4672 5108 4678 5160
rect 4884 5151 4942 5157
rect 4884 5117 4896 5151
rect 4930 5148 4942 5151
rect 5810 5148 5816 5160
rect 4930 5120 5816 5148
rect 4930 5117 4942 5120
rect 4884 5111 4942 5117
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 7558 5108 7564 5160
rect 7616 5148 7622 5160
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 7616 5120 7941 5148
rect 7616 5108 7622 5120
rect 7929 5117 7941 5120
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 8018 5108 8024 5160
rect 8076 5148 8082 5160
rect 8076 5120 8892 5148
rect 8076 5108 8082 5120
rect 8386 5040 8392 5092
rect 8444 5040 8450 5092
rect 8864 5089 8892 5120
rect 9030 5108 9036 5160
rect 9088 5108 9094 5160
rect 8849 5083 8907 5089
rect 8849 5049 8861 5083
rect 8895 5049 8907 5083
rect 10980 5080 11008 5256
rect 11146 5244 11152 5296
rect 11204 5284 11210 5296
rect 11698 5284 11704 5296
rect 11204 5256 11704 5284
rect 11204 5244 11210 5256
rect 11698 5244 11704 5256
rect 11756 5244 11762 5296
rect 13556 5225 13584 5324
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 14737 5355 14795 5361
rect 14737 5321 14749 5355
rect 14783 5352 14795 5355
rect 18046 5352 18052 5364
rect 14783 5324 18052 5352
rect 14783 5321 14795 5324
rect 14737 5315 14795 5321
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 19058 5312 19064 5364
rect 19116 5352 19122 5364
rect 19116 5324 19656 5352
rect 19116 5312 19122 5324
rect 19628 5284 19656 5324
rect 20070 5312 20076 5364
rect 20128 5312 20134 5364
rect 20809 5355 20867 5361
rect 20809 5321 20821 5355
rect 20855 5352 20867 5355
rect 21634 5352 21640 5364
rect 20855 5324 21640 5352
rect 20855 5321 20867 5324
rect 20809 5315 20867 5321
rect 21634 5312 21640 5324
rect 21692 5312 21698 5364
rect 23569 5355 23627 5361
rect 23569 5321 23581 5355
rect 23615 5352 23627 5355
rect 25406 5352 25412 5364
rect 23615 5324 25412 5352
rect 23615 5321 23627 5324
rect 23569 5315 23627 5321
rect 25406 5312 25412 5324
rect 25464 5312 25470 5364
rect 19628 5256 20484 5284
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 13630 5176 13636 5228
rect 13688 5216 13694 5228
rect 14090 5216 14096 5228
rect 13688 5188 14096 5216
rect 13688 5176 13694 5188
rect 14090 5176 14096 5188
rect 14148 5216 14154 5228
rect 14148 5188 14596 5216
rect 14148 5176 14154 5188
rect 11606 5108 11612 5160
rect 11664 5148 11670 5160
rect 12713 5151 12771 5157
rect 12713 5148 12725 5151
rect 11664 5120 12725 5148
rect 11664 5108 11670 5120
rect 12713 5117 12725 5120
rect 12759 5117 12771 5151
rect 12713 5111 12771 5117
rect 12986 5108 12992 5160
rect 13044 5148 13050 5160
rect 14568 5157 14596 5188
rect 16574 5176 16580 5228
rect 16632 5216 16638 5228
rect 16632 5188 17172 5216
rect 16632 5176 16638 5188
rect 14277 5151 14335 5157
rect 14277 5148 14289 5151
rect 13044 5120 14289 5148
rect 13044 5108 13050 5120
rect 14277 5117 14289 5120
rect 14323 5117 14335 5151
rect 14277 5111 14335 5117
rect 14553 5151 14611 5157
rect 14553 5117 14565 5151
rect 14599 5148 14611 5151
rect 14829 5151 14887 5157
rect 14829 5148 14841 5151
rect 14599 5120 14841 5148
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 14829 5117 14841 5120
rect 14875 5117 14887 5151
rect 14829 5111 14887 5117
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5117 15991 5151
rect 15933 5111 15991 5117
rect 16485 5151 16543 5157
rect 16485 5117 16497 5151
rect 16531 5148 16543 5151
rect 16850 5148 16856 5160
rect 16531 5120 16856 5148
rect 16531 5117 16543 5120
rect 16485 5111 16543 5117
rect 12250 5080 12256 5092
rect 10980 5052 12256 5080
rect 8849 5043 8907 5049
rect 12250 5040 12256 5052
rect 12308 5040 12314 5092
rect 12434 5040 12440 5092
rect 12492 5089 12498 5092
rect 12492 5043 12504 5089
rect 15948 5080 15976 5111
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 17144 5157 17172 5188
rect 17129 5151 17187 5157
rect 17129 5117 17141 5151
rect 17175 5148 17187 5151
rect 17954 5148 17960 5160
rect 17175 5120 17960 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 17954 5108 17960 5120
rect 18012 5148 18018 5160
rect 18506 5148 18512 5160
rect 18012 5120 18512 5148
rect 18012 5108 18018 5120
rect 18506 5108 18512 5120
rect 18564 5108 18570 5160
rect 18693 5151 18751 5157
rect 18693 5117 18705 5151
rect 18739 5148 18751 5151
rect 19886 5148 19892 5160
rect 18739 5120 19892 5148
rect 18739 5117 18751 5120
rect 18693 5111 18751 5117
rect 19886 5108 19892 5120
rect 19944 5108 19950 5160
rect 20165 5151 20223 5157
rect 20165 5117 20177 5151
rect 20211 5117 20223 5151
rect 20165 5111 20223 5117
rect 16942 5080 16948 5092
rect 14108 5052 16948 5080
rect 12492 5040 12498 5043
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 8589 5015 8647 5021
rect 8589 5012 8601 5015
rect 7800 4984 8601 5012
rect 7800 4972 7806 4984
rect 8589 4981 8601 4984
rect 8635 4981 8647 5015
rect 8589 4975 8647 4981
rect 11330 4972 11336 5024
rect 11388 5012 11394 5024
rect 14108 5012 14136 5052
rect 16942 5040 16948 5052
rect 17000 5040 17006 5092
rect 18966 5089 18972 5092
rect 17037 5083 17095 5089
rect 17037 5049 17049 5083
rect 17083 5080 17095 5083
rect 17374 5083 17432 5089
rect 17374 5080 17386 5083
rect 17083 5052 17386 5080
rect 17083 5049 17095 5052
rect 17037 5043 17095 5049
rect 17374 5049 17386 5052
rect 17420 5049 17432 5083
rect 17374 5043 17432 5049
rect 18960 5043 18972 5089
rect 19024 5080 19030 5092
rect 19024 5052 19060 5080
rect 18966 5040 18972 5043
rect 19024 5040 19030 5052
rect 19334 5040 19340 5092
rect 19392 5080 19398 5092
rect 20180 5080 20208 5111
rect 20254 5108 20260 5160
rect 20312 5148 20318 5160
rect 20456 5157 20484 5256
rect 21726 5244 21732 5296
rect 21784 5284 21790 5296
rect 22373 5287 22431 5293
rect 22373 5284 22385 5287
rect 21784 5256 22385 5284
rect 21784 5244 21790 5256
rect 22373 5253 22385 5256
rect 22419 5253 22431 5287
rect 22373 5247 22431 5253
rect 23750 5244 23756 5296
rect 23808 5284 23814 5296
rect 23845 5287 23903 5293
rect 23845 5284 23857 5287
rect 23808 5256 23857 5284
rect 23808 5244 23814 5256
rect 23845 5253 23857 5256
rect 23891 5253 23903 5287
rect 23845 5247 23903 5253
rect 20349 5151 20407 5157
rect 20349 5148 20361 5151
rect 20312 5120 20361 5148
rect 20312 5108 20318 5120
rect 20349 5117 20361 5120
rect 20395 5117 20407 5151
rect 20349 5111 20407 5117
rect 20441 5151 20499 5157
rect 20441 5117 20453 5151
rect 20487 5117 20499 5151
rect 20441 5111 20499 5117
rect 20533 5151 20591 5157
rect 20533 5117 20545 5151
rect 20579 5148 20591 5151
rect 20990 5148 20996 5160
rect 20579 5120 20996 5148
rect 20579 5117 20591 5120
rect 20533 5111 20591 5117
rect 20990 5108 20996 5120
rect 21048 5108 21054 5160
rect 21082 5108 21088 5160
rect 21140 5108 21146 5160
rect 21266 5108 21272 5160
rect 21324 5148 21330 5160
rect 22922 5148 22928 5160
rect 21324 5120 22928 5148
rect 21324 5108 21330 5120
rect 22922 5108 22928 5120
rect 22980 5108 22986 5160
rect 23106 5108 23112 5160
rect 23164 5108 23170 5160
rect 23198 5108 23204 5160
rect 23256 5108 23262 5160
rect 23293 5151 23351 5157
rect 23293 5117 23305 5151
rect 23339 5148 23351 5151
rect 23474 5148 23480 5160
rect 23339 5120 23480 5148
rect 23339 5117 23351 5120
rect 23293 5111 23351 5117
rect 23474 5108 23480 5120
rect 23532 5108 23538 5160
rect 24670 5108 24676 5160
rect 24728 5148 24734 5160
rect 25225 5151 25283 5157
rect 25225 5148 25237 5151
rect 24728 5120 25237 5148
rect 24728 5108 24734 5120
rect 25225 5117 25237 5120
rect 25271 5117 25283 5151
rect 25225 5111 25283 5117
rect 25866 5108 25872 5160
rect 25924 5108 25930 5160
rect 21358 5080 21364 5092
rect 19392 5052 21364 5080
rect 19392 5040 19398 5052
rect 21358 5040 21364 5052
rect 21416 5040 21422 5092
rect 22370 5040 22376 5092
rect 22428 5080 22434 5092
rect 23216 5080 23244 5108
rect 23566 5080 23572 5092
rect 22428 5052 23572 5080
rect 22428 5040 22434 5052
rect 23566 5040 23572 5052
rect 23624 5040 23630 5092
rect 24980 5083 25038 5089
rect 24980 5049 24992 5083
rect 25026 5080 25038 5083
rect 25317 5083 25375 5089
rect 25317 5080 25329 5083
rect 25026 5052 25329 5080
rect 25026 5049 25038 5052
rect 24980 5043 25038 5049
rect 25317 5049 25329 5052
rect 25363 5049 25375 5083
rect 25317 5043 25375 5049
rect 11388 4984 14136 5012
rect 14185 5015 14243 5021
rect 11388 4972 11394 4984
rect 14185 4981 14197 5015
rect 14231 5012 14243 5015
rect 14369 5015 14427 5021
rect 14369 5012 14381 5015
rect 14231 4984 14381 5012
rect 14231 4981 14243 4984
rect 14185 4975 14243 4981
rect 14369 4981 14381 4984
rect 14415 4981 14427 5015
rect 14369 4975 14427 4981
rect 14458 4972 14464 5024
rect 14516 5012 14522 5024
rect 14642 5012 14648 5024
rect 14516 4984 14648 5012
rect 14516 4972 14522 4984
rect 14642 4972 14648 4984
rect 14700 5012 14706 5024
rect 15013 5015 15071 5021
rect 15013 5012 15025 5015
rect 14700 4984 15025 5012
rect 14700 4972 14706 4984
rect 15013 4981 15025 4984
rect 15059 4981 15071 5015
rect 15013 4975 15071 4981
rect 15562 4972 15568 5024
rect 15620 5012 15626 5024
rect 16117 5015 16175 5021
rect 16117 5012 16129 5015
rect 15620 4984 16129 5012
rect 15620 4972 15626 4984
rect 16117 4981 16129 4984
rect 16163 5012 16175 5015
rect 17494 5012 17500 5024
rect 16163 4984 17500 5012
rect 16163 4981 16175 4984
rect 16117 4975 16175 4981
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 18509 5015 18567 5021
rect 18509 4981 18521 5015
rect 18555 5012 18567 5015
rect 19978 5012 19984 5024
rect 18555 4984 19984 5012
rect 18555 4981 18567 4984
rect 18509 4975 18567 4981
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 20254 4972 20260 5024
rect 20312 5012 20318 5024
rect 20530 5012 20536 5024
rect 20312 4984 20536 5012
rect 20312 4972 20318 4984
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 22830 5012 22836 5024
rect 20956 4984 22836 5012
rect 20956 4972 20962 4984
rect 22830 4972 22836 4984
rect 22888 4972 22894 5024
rect 552 4922 27576 4944
rect 552 4870 7114 4922
rect 7166 4870 7178 4922
rect 7230 4870 7242 4922
rect 7294 4870 7306 4922
rect 7358 4870 7370 4922
rect 7422 4870 13830 4922
rect 13882 4870 13894 4922
rect 13946 4870 13958 4922
rect 14010 4870 14022 4922
rect 14074 4870 14086 4922
rect 14138 4870 20546 4922
rect 20598 4870 20610 4922
rect 20662 4870 20674 4922
rect 20726 4870 20738 4922
rect 20790 4870 20802 4922
rect 20854 4870 27262 4922
rect 27314 4870 27326 4922
rect 27378 4870 27390 4922
rect 27442 4870 27454 4922
rect 27506 4870 27518 4922
rect 27570 4870 27576 4922
rect 552 4848 27576 4870
rect 7558 4768 7564 4820
rect 7616 4768 7622 4820
rect 8294 4768 8300 4820
rect 8352 4808 8358 4820
rect 12989 4811 13047 4817
rect 8352 4780 8800 4808
rect 8352 4768 8358 4780
rect 8113 4743 8171 4749
rect 8113 4740 8125 4743
rect 6104 4712 8125 4740
rect 5258 4632 5264 4684
rect 5316 4632 5322 4684
rect 6104 4681 6132 4712
rect 8113 4709 8125 4712
rect 8159 4740 8171 4743
rect 8772 4740 8800 4780
rect 12989 4777 13001 4811
rect 13035 4808 13047 4811
rect 18598 4808 18604 4820
rect 13035 4780 18604 4808
rect 13035 4777 13047 4780
rect 12989 4771 13047 4777
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 22646 4808 22652 4820
rect 22066 4780 22652 4808
rect 9950 4740 9956 4752
rect 8159 4712 8622 4740
rect 8159 4709 8171 4712
rect 8113 4703 8171 4709
rect 5445 4675 5503 4681
rect 5445 4641 5457 4675
rect 5491 4672 5503 4675
rect 6089 4675 6147 4681
rect 6089 4672 6101 4675
rect 5491 4644 6101 4672
rect 5491 4641 5503 4644
rect 5445 4635 5503 4641
rect 6089 4641 6101 4644
rect 6135 4641 6147 4675
rect 6089 4635 6147 4641
rect 6270 4632 6276 4684
rect 6328 4632 6334 4684
rect 6362 4632 6368 4684
rect 6420 4672 6426 4684
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 6420 4644 7389 4672
rect 6420 4632 6426 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 7466 4632 7472 4684
rect 7524 4632 7530 4684
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4641 7711 4675
rect 7653 4635 7711 4641
rect 7745 4675 7803 4681
rect 7745 4641 7757 4675
rect 7791 4641 7803 4675
rect 7745 4635 7803 4641
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4604 6515 4607
rect 6546 4604 6552 4616
rect 6503 4576 6552 4604
rect 6503 4573 6515 4576
rect 6457 4567 6515 4573
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 7668 4536 7696 4635
rect 7760 4604 7788 4635
rect 7834 4632 7840 4684
rect 7892 4632 7898 4684
rect 8294 4632 8300 4684
rect 8352 4632 8358 4684
rect 8594 4681 8622 4712
rect 8772 4712 9956 4740
rect 8772 4681 8800 4712
rect 9950 4700 9956 4712
rect 10008 4700 10014 4752
rect 11333 4743 11391 4749
rect 11333 4709 11345 4743
rect 11379 4740 11391 4743
rect 12434 4740 12440 4752
rect 11379 4712 12440 4740
rect 11379 4709 11391 4712
rect 11333 4703 11391 4709
rect 12434 4700 12440 4712
rect 12492 4700 12498 4752
rect 12894 4740 12900 4752
rect 12544 4712 12900 4740
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4641 8631 4675
rect 8573 4635 8631 4641
rect 8757 4675 8815 4681
rect 8757 4641 8769 4675
rect 8803 4641 8815 4675
rect 8757 4635 8815 4641
rect 9030 4632 9036 4684
rect 9088 4632 9094 4684
rect 12544 4681 12572 4712
rect 12894 4700 12900 4712
rect 12952 4740 12958 4752
rect 13541 4743 13599 4749
rect 12952 4712 13032 4740
rect 12952 4700 12958 4712
rect 12529 4675 12587 4681
rect 12529 4641 12541 4675
rect 12575 4641 12587 4675
rect 12529 4635 12587 4641
rect 12621 4675 12679 4681
rect 12621 4641 12633 4675
rect 12667 4672 12679 4675
rect 12710 4672 12716 4684
rect 12667 4644 12716 4672
rect 12667 4641 12679 4644
rect 12621 4635 12679 4641
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 12802 4632 12808 4684
rect 12860 4632 12866 4684
rect 13004 4672 13032 4712
rect 13541 4709 13553 4743
rect 13587 4740 13599 4743
rect 13587 4712 17356 4740
rect 13587 4709 13599 4712
rect 13541 4703 13599 4709
rect 13081 4675 13139 4681
rect 13081 4672 13093 4675
rect 13004 4644 13093 4672
rect 13081 4641 13093 4644
rect 13127 4641 13139 4675
rect 13081 4635 13139 4641
rect 13170 4632 13176 4684
rect 13228 4632 13234 4684
rect 13357 4675 13415 4681
rect 13357 4641 13369 4675
rect 13403 4672 13415 4675
rect 13630 4672 13636 4684
rect 13403 4644 13636 4672
rect 13403 4641 13415 4644
rect 13357 4635 13415 4641
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 13998 4632 14004 4684
rect 14056 4632 14062 4684
rect 14093 4675 14151 4681
rect 14093 4641 14105 4675
rect 14139 4641 14151 4675
rect 14093 4635 14151 4641
rect 14277 4675 14335 4681
rect 14277 4641 14289 4675
rect 14323 4672 14335 4675
rect 14458 4672 14464 4684
rect 14323 4644 14464 4672
rect 14323 4641 14335 4644
rect 14277 4635 14335 4641
rect 9582 4604 9588 4616
rect 7760 4576 9588 4604
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 10137 4607 10195 4613
rect 10137 4573 10149 4607
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4604 10839 4607
rect 14108 4604 14136 4635
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 14826 4681 14832 4684
rect 14820 4635 14832 4681
rect 14826 4632 14832 4635
rect 14884 4632 14890 4684
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 16117 4675 16175 4681
rect 16117 4672 16129 4675
rect 15252 4644 16129 4672
rect 15252 4632 15258 4644
rect 16117 4641 16129 4644
rect 16163 4641 16175 4675
rect 16117 4635 16175 4641
rect 17129 4675 17187 4681
rect 17129 4641 17141 4675
rect 17175 4641 17187 4675
rect 17129 4635 17187 4641
rect 10827 4576 14136 4604
rect 10827 4573 10839 4576
rect 10781 4567 10839 4573
rect 8018 4536 8024 4548
rect 7668 4508 8024 4536
rect 8018 4496 8024 4508
rect 8076 4496 8082 4548
rect 9122 4496 9128 4548
rect 9180 4536 9186 4548
rect 10152 4536 10180 4567
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 16761 4607 16819 4613
rect 16761 4573 16773 4607
rect 16807 4573 16819 4607
rect 16761 4567 16819 4573
rect 9180 4508 10180 4536
rect 9180 4496 9186 4508
rect 11514 4496 11520 4548
rect 11572 4536 11578 4548
rect 11701 4539 11759 4545
rect 11701 4536 11713 4539
rect 11572 4508 11713 4536
rect 11572 4496 11578 4508
rect 11701 4505 11713 4508
rect 11747 4536 11759 4539
rect 11790 4536 11796 4548
rect 11747 4508 11796 4536
rect 11747 4505 11759 4508
rect 11701 4499 11759 4505
rect 11790 4496 11796 4508
rect 11848 4496 11854 4548
rect 12802 4496 12808 4548
rect 12860 4536 12866 4548
rect 13630 4536 13636 4548
rect 12860 4508 13636 4536
rect 12860 4496 12866 4508
rect 13630 4496 13636 4508
rect 13688 4496 13694 4548
rect 15933 4539 15991 4545
rect 15933 4505 15945 4539
rect 15979 4536 15991 4539
rect 16776 4536 16804 4567
rect 16850 4564 16856 4616
rect 16908 4564 16914 4616
rect 17144 4604 17172 4635
rect 17218 4632 17224 4684
rect 17276 4632 17282 4684
rect 17328 4681 17356 4712
rect 19426 4700 19432 4752
rect 19484 4700 19490 4752
rect 20533 4743 20591 4749
rect 20533 4709 20545 4743
rect 20579 4740 20591 4743
rect 22066 4740 22094 4780
rect 22646 4768 22652 4780
rect 22704 4768 22710 4820
rect 22922 4768 22928 4820
rect 22980 4808 22986 4820
rect 22980 4780 23520 4808
rect 22980 4768 22986 4780
rect 20579 4712 22094 4740
rect 22296 4712 23428 4740
rect 20579 4709 20591 4712
rect 20533 4703 20591 4709
rect 17313 4675 17371 4681
rect 17313 4641 17325 4675
rect 17359 4641 17371 4675
rect 17313 4635 17371 4641
rect 17494 4632 17500 4684
rect 17552 4632 17558 4684
rect 19978 4632 19984 4684
rect 20036 4672 20042 4684
rect 20073 4675 20131 4681
rect 20073 4672 20085 4675
rect 20036 4644 20085 4672
rect 20036 4632 20042 4644
rect 20073 4641 20085 4644
rect 20119 4641 20131 4675
rect 20073 4635 20131 4641
rect 20254 4632 20260 4684
rect 20312 4632 20318 4684
rect 20346 4632 20352 4684
rect 20404 4672 20410 4684
rect 20625 4675 20683 4681
rect 20404 4644 20449 4672
rect 20404 4632 20410 4644
rect 20625 4641 20637 4675
rect 20671 4641 20683 4675
rect 20625 4635 20683 4641
rect 20763 4675 20821 4681
rect 20763 4641 20775 4675
rect 20809 4672 20821 4675
rect 20898 4672 20904 4684
rect 20809 4644 20904 4672
rect 20809 4641 20821 4644
rect 20763 4635 20821 4641
rect 19521 4607 19579 4613
rect 19521 4604 19533 4607
rect 17144 4576 19533 4604
rect 19521 4573 19533 4576
rect 19567 4573 19579 4607
rect 19521 4567 19579 4573
rect 20640 4536 20668 4635
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 22296 4681 22324 4712
rect 22281 4675 22339 4681
rect 22281 4641 22293 4675
rect 22327 4641 22339 4675
rect 22281 4635 22339 4641
rect 22370 4632 22376 4684
rect 22428 4632 22434 4684
rect 22465 4675 22523 4681
rect 22465 4641 22477 4675
rect 22511 4641 22523 4675
rect 22465 4635 22523 4641
rect 22649 4675 22707 4681
rect 22649 4641 22661 4675
rect 22695 4641 22707 4675
rect 22649 4635 22707 4641
rect 21913 4607 21971 4613
rect 21913 4573 21925 4607
rect 21959 4604 21971 4607
rect 22005 4607 22063 4613
rect 22005 4604 22017 4607
rect 21959 4576 22017 4604
rect 21959 4573 21971 4576
rect 21913 4567 21971 4573
rect 22005 4573 22017 4576
rect 22051 4573 22063 4607
rect 22005 4567 22063 4573
rect 15979 4508 20668 4536
rect 20901 4539 20959 4545
rect 15979 4505 15991 4508
rect 15933 4499 15991 4505
rect 20901 4505 20913 4539
rect 20947 4536 20959 4539
rect 22480 4536 22508 4635
rect 20947 4508 22508 4536
rect 20947 4505 20959 4508
rect 20901 4499 20959 4505
rect 4890 4428 4896 4480
rect 4948 4468 4954 4480
rect 5261 4471 5319 4477
rect 5261 4468 5273 4471
rect 4948 4440 5273 4468
rect 4948 4428 4954 4440
rect 5261 4437 5273 4440
rect 5307 4437 5319 4471
rect 5261 4431 5319 4437
rect 8481 4471 8539 4477
rect 8481 4437 8493 4471
rect 8527 4468 8539 4471
rect 8570 4468 8576 4480
rect 8527 4440 8576 4468
rect 8527 4437 8539 4440
rect 8481 4431 8539 4437
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 8662 4428 8668 4480
rect 8720 4428 8726 4480
rect 9217 4471 9275 4477
rect 9217 4437 9229 4471
rect 9263 4468 9275 4471
rect 9306 4468 9312 4480
rect 9263 4440 9312 4468
rect 9263 4437 9275 4440
rect 9217 4431 9275 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 10870 4428 10876 4480
rect 10928 4468 10934 4480
rect 11149 4471 11207 4477
rect 11149 4468 11161 4471
rect 10928 4440 11161 4468
rect 10928 4428 10934 4440
rect 11149 4437 11161 4440
rect 11195 4437 11207 4471
rect 11149 4431 11207 4437
rect 11330 4428 11336 4480
rect 11388 4428 11394 4480
rect 14461 4471 14519 4477
rect 14461 4437 14473 4471
rect 14507 4468 14519 4471
rect 15286 4468 15292 4480
rect 14507 4440 15292 4468
rect 14507 4437 14519 4440
rect 14461 4431 14519 4437
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 18141 4471 18199 4477
rect 18141 4437 18153 4471
rect 18187 4468 18199 4471
rect 18506 4468 18512 4480
rect 18187 4440 18512 4468
rect 18187 4437 18199 4440
rect 18141 4431 18199 4437
rect 18506 4428 18512 4440
rect 18564 4428 18570 4480
rect 21082 4428 21088 4480
rect 21140 4468 21146 4480
rect 21269 4471 21327 4477
rect 21269 4468 21281 4471
rect 21140 4440 21281 4468
rect 21140 4428 21146 4440
rect 21269 4437 21281 4440
rect 21315 4437 21327 4471
rect 21269 4431 21327 4437
rect 21358 4428 21364 4480
rect 21416 4468 21422 4480
rect 21910 4468 21916 4480
rect 21416 4440 21916 4468
rect 21416 4428 21422 4440
rect 21910 4428 21916 4440
rect 21968 4468 21974 4480
rect 22664 4468 22692 4635
rect 22738 4564 22744 4616
rect 22796 4564 22802 4616
rect 23400 4477 23428 4712
rect 23492 4681 23520 4780
rect 23750 4768 23756 4820
rect 23808 4768 23814 4820
rect 24121 4811 24179 4817
rect 24121 4777 24133 4811
rect 24167 4808 24179 4811
rect 25866 4808 25872 4820
rect 24167 4780 25872 4808
rect 24167 4777 24179 4780
rect 24121 4771 24179 4777
rect 25866 4768 25872 4780
rect 25924 4768 25930 4820
rect 23768 4740 23796 4768
rect 23768 4712 24808 4740
rect 23477 4675 23535 4681
rect 23477 4641 23489 4675
rect 23523 4641 23535 4675
rect 23477 4635 23535 4641
rect 23658 4632 23664 4684
rect 23716 4632 23722 4684
rect 24780 4681 24808 4712
rect 23753 4675 23811 4681
rect 23753 4641 23765 4675
rect 23799 4641 23811 4675
rect 23753 4635 23811 4641
rect 23845 4675 23903 4681
rect 23845 4641 23857 4675
rect 23891 4672 23903 4675
rect 24213 4675 24271 4681
rect 24213 4672 24225 4675
rect 23891 4644 24225 4672
rect 23891 4641 23903 4644
rect 23845 4635 23903 4641
rect 24213 4641 24225 4644
rect 24259 4641 24271 4675
rect 24213 4635 24271 4641
rect 24765 4675 24823 4681
rect 24765 4641 24777 4675
rect 24811 4641 24823 4675
rect 24765 4635 24823 4641
rect 23566 4564 23572 4616
rect 23624 4604 23630 4616
rect 23768 4604 23796 4635
rect 23624 4576 23796 4604
rect 23624 4564 23630 4576
rect 21968 4440 22692 4468
rect 23385 4471 23443 4477
rect 21968 4428 21974 4440
rect 23385 4437 23397 4471
rect 23431 4468 23443 4471
rect 24302 4468 24308 4480
rect 23431 4440 24308 4468
rect 23431 4437 23443 4440
rect 23385 4431 23443 4437
rect 24302 4428 24308 4440
rect 24360 4428 24366 4480
rect 552 4378 27416 4400
rect 552 4326 3756 4378
rect 3808 4326 3820 4378
rect 3872 4326 3884 4378
rect 3936 4326 3948 4378
rect 4000 4326 4012 4378
rect 4064 4326 10472 4378
rect 10524 4326 10536 4378
rect 10588 4326 10600 4378
rect 10652 4326 10664 4378
rect 10716 4326 10728 4378
rect 10780 4326 17188 4378
rect 17240 4326 17252 4378
rect 17304 4326 17316 4378
rect 17368 4326 17380 4378
rect 17432 4326 17444 4378
rect 17496 4326 23904 4378
rect 23956 4326 23968 4378
rect 24020 4326 24032 4378
rect 24084 4326 24096 4378
rect 24148 4326 24160 4378
rect 24212 4326 27416 4378
rect 552 4304 27416 4326
rect 8570 4224 8576 4276
rect 8628 4224 8634 4276
rect 8757 4267 8815 4273
rect 8757 4233 8769 4267
rect 8803 4264 8815 4267
rect 9030 4264 9036 4276
rect 8803 4236 9036 4264
rect 8803 4233 8815 4236
rect 8757 4227 8815 4233
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 9950 4224 9956 4276
rect 10008 4264 10014 4276
rect 10413 4267 10471 4273
rect 10413 4264 10425 4267
rect 10008 4236 10425 4264
rect 10008 4224 10014 4236
rect 10413 4233 10425 4236
rect 10459 4264 10471 4267
rect 12437 4267 12495 4273
rect 10459 4236 12112 4264
rect 10459 4233 10471 4236
rect 10413 4227 10471 4233
rect 5997 4199 6055 4205
rect 5997 4165 6009 4199
rect 6043 4165 6055 4199
rect 5997 4159 6055 4165
rect 6012 4128 6040 4159
rect 8110 4156 8116 4208
rect 8168 4156 8174 4208
rect 6546 4128 6552 4140
rect 6012 4100 6552 4128
rect 6546 4088 6552 4100
rect 6604 4128 6610 4140
rect 6604 4100 7696 4128
rect 6604 4088 6610 4100
rect 4614 4020 4620 4072
rect 4672 4060 4678 4072
rect 4672 4032 5304 4060
rect 4672 4020 4678 4032
rect 4890 4001 4896 4004
rect 4884 3992 4896 4001
rect 4851 3964 4896 3992
rect 4884 3955 4896 3964
rect 4890 3952 4896 3955
rect 4948 3952 4954 4004
rect 5276 3992 5304 4032
rect 6362 4020 6368 4072
rect 6420 4060 6426 4072
rect 6457 4063 6515 4069
rect 6457 4060 6469 4063
rect 6420 4032 6469 4060
rect 6420 4020 6426 4032
rect 6457 4029 6469 4032
rect 6503 4029 6515 4063
rect 6457 4023 6515 4029
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4060 7343 4063
rect 7466 4060 7472 4072
rect 7331 4032 7472 4060
rect 7331 4029 7343 4032
rect 7285 4023 7343 4029
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 7668 4069 7696 4100
rect 7926 4088 7932 4140
rect 7984 4088 7990 4140
rect 12084 4128 12112 4236
rect 12437 4233 12449 4267
rect 12483 4264 12495 4267
rect 12526 4264 12532 4276
rect 12483 4236 12532 4264
rect 12483 4233 12495 4236
rect 12437 4227 12495 4233
rect 12526 4224 12532 4236
rect 12584 4264 12590 4276
rect 13170 4264 13176 4276
rect 12584 4236 13176 4264
rect 12584 4224 12590 4236
rect 13170 4224 13176 4236
rect 13228 4224 13234 4276
rect 14826 4224 14832 4276
rect 14884 4224 14890 4276
rect 21726 4264 21732 4276
rect 20824 4236 21732 4264
rect 12250 4156 12256 4208
rect 12308 4196 12314 4208
rect 13538 4196 13544 4208
rect 12308 4168 13544 4196
rect 12308 4156 12314 4168
rect 13538 4156 13544 4168
rect 13596 4156 13602 4208
rect 15212 4168 15792 4196
rect 8036 4100 9168 4128
rect 12084 4100 12434 4128
rect 7653 4063 7711 4069
rect 7653 4029 7665 4063
rect 7699 4060 7711 4063
rect 8036 4060 8064 4100
rect 9140 4072 9168 4100
rect 7699 4032 8064 4060
rect 8205 4063 8263 4069
rect 7699 4029 7711 4032
rect 7653 4023 7711 4029
rect 8205 4029 8217 4063
rect 8251 4060 8263 4063
rect 8294 4060 8300 4072
rect 8251 4032 8300 4060
rect 8251 4029 8263 4032
rect 8205 4023 8263 4029
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 9033 4063 9091 4069
rect 9033 4029 9045 4063
rect 9079 4029 9091 4063
rect 9033 4023 9091 4029
rect 6822 3992 6828 4004
rect 5276 3964 6828 3992
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 7742 3992 7748 4004
rect 7484 3964 7748 3992
rect 7006 3884 7012 3936
rect 7064 3924 7070 3936
rect 7484 3933 7512 3964
rect 7742 3952 7748 3964
rect 7800 3952 7806 4004
rect 7837 3995 7895 4001
rect 7837 3961 7849 3995
rect 7883 3992 7895 3995
rect 7883 3964 8248 3992
rect 7883 3961 7895 3964
rect 7837 3955 7895 3961
rect 8220 3936 8248 3964
rect 8386 3952 8392 4004
rect 8444 3952 8450 4004
rect 7101 3927 7159 3933
rect 7101 3924 7113 3927
rect 7064 3896 7113 3924
rect 7064 3884 7070 3896
rect 7101 3893 7113 3896
rect 7147 3893 7159 3927
rect 7101 3887 7159 3893
rect 7469 3927 7527 3933
rect 7469 3893 7481 3927
rect 7515 3893 7527 3927
rect 7469 3887 7527 3893
rect 7558 3884 7564 3936
rect 7616 3884 7622 3936
rect 7926 3884 7932 3936
rect 7984 3884 7990 3936
rect 8202 3884 8208 3936
rect 8260 3884 8266 3936
rect 8570 3884 8576 3936
rect 8628 3933 8634 3936
rect 8628 3927 8647 3933
rect 8635 3893 8647 3927
rect 9048 3924 9076 4023
rect 9122 4020 9128 4072
rect 9180 4020 9186 4072
rect 9306 4069 9312 4072
rect 9300 4023 9312 4069
rect 9364 4060 9370 4072
rect 10781 4063 10839 4069
rect 9364 4032 9400 4060
rect 9306 4020 9312 4023
rect 9364 4020 9370 4032
rect 10781 4029 10793 4063
rect 10827 4060 10839 4063
rect 10870 4060 10876 4072
rect 10827 4032 10876 4060
rect 10827 4029 10839 4032
rect 10781 4023 10839 4029
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 11057 4063 11115 4069
rect 11057 4029 11069 4063
rect 11103 4060 11115 4063
rect 11606 4060 11612 4072
rect 11103 4032 11612 4060
rect 11103 4029 11115 4032
rect 11057 4023 11115 4029
rect 11072 3992 11100 4023
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 11302 3995 11360 4001
rect 11302 3992 11314 3995
rect 9416 3964 11100 3992
rect 11164 3964 11314 3992
rect 9416 3924 9444 3964
rect 9048 3896 9444 3924
rect 10965 3927 11023 3933
rect 8628 3887 8647 3893
rect 10965 3893 10977 3927
rect 11011 3924 11023 3927
rect 11164 3924 11192 3964
rect 11302 3961 11314 3964
rect 11348 3961 11360 3995
rect 12406 3992 12434 4100
rect 12710 4020 12716 4072
rect 12768 4060 12774 4072
rect 13541 4063 13599 4069
rect 13541 4060 13553 4063
rect 12768 4032 13553 4060
rect 12768 4020 12774 4032
rect 13541 4029 13553 4032
rect 13587 4029 13599 4063
rect 13541 4023 13599 4029
rect 13630 4020 13636 4072
rect 13688 4060 13694 4072
rect 14093 4063 14151 4069
rect 14093 4060 14105 4063
rect 13688 4032 14105 4060
rect 13688 4020 13694 4032
rect 14093 4029 14105 4032
rect 14139 4029 14151 4063
rect 14093 4023 14151 4029
rect 14182 4020 14188 4072
rect 14240 4060 14246 4072
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 14240 4032 14289 4060
rect 14240 4020 14246 4032
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 14277 4023 14335 4029
rect 14458 4020 14464 4072
rect 14516 4060 14522 4072
rect 14553 4063 14611 4069
rect 14553 4060 14565 4063
rect 14516 4032 14565 4060
rect 14516 4020 14522 4032
rect 14553 4029 14565 4032
rect 14599 4060 14611 4063
rect 15010 4060 15016 4072
rect 14599 4032 15016 4060
rect 14599 4029 14611 4032
rect 14553 4023 14611 4029
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 15102 4020 15108 4072
rect 15160 4020 15166 4072
rect 15212 4069 15240 4168
rect 15396 4140 15424 4168
rect 15378 4088 15384 4140
rect 15436 4088 15442 4140
rect 15654 4128 15660 4140
rect 15488 4100 15660 4128
rect 15197 4063 15255 4069
rect 15197 4029 15209 4063
rect 15243 4029 15255 4063
rect 15197 4023 15255 4029
rect 15286 4020 15292 4072
rect 15344 4020 15350 4072
rect 15488 4069 15516 4100
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 15764 4128 15792 4168
rect 15764 4100 16252 4128
rect 15473 4063 15531 4069
rect 15473 4029 15485 4063
rect 15519 4029 15531 4063
rect 15473 4023 15531 4029
rect 15562 4020 15568 4072
rect 15620 4060 15626 4072
rect 16224 4069 16252 4100
rect 19978 4088 19984 4140
rect 20036 4128 20042 4140
rect 20824 4137 20852 4236
rect 21726 4224 21732 4236
rect 21784 4224 21790 4276
rect 22189 4267 22247 4273
rect 22189 4233 22201 4267
rect 22235 4264 22247 4267
rect 22738 4264 22744 4276
rect 22235 4236 22744 4264
rect 22235 4233 22247 4236
rect 22189 4227 22247 4233
rect 22738 4224 22744 4236
rect 22796 4224 22802 4276
rect 22830 4224 22836 4276
rect 22888 4264 22894 4276
rect 23290 4264 23296 4276
rect 22888 4236 23296 4264
rect 22888 4224 22894 4236
rect 23290 4224 23296 4236
rect 23348 4224 23354 4276
rect 22646 4156 22652 4208
rect 22704 4196 22710 4208
rect 22704 4168 23796 4196
rect 22704 4156 22710 4168
rect 20809 4131 20867 4137
rect 20809 4128 20821 4131
rect 20036 4100 20821 4128
rect 20036 4088 20042 4100
rect 20809 4097 20821 4100
rect 20855 4097 20867 4131
rect 20809 4091 20867 4097
rect 23198 4088 23204 4140
rect 23256 4128 23262 4140
rect 23658 4128 23664 4140
rect 23256 4100 23664 4128
rect 23256 4088 23262 4100
rect 23658 4088 23664 4100
rect 23716 4088 23722 4140
rect 23768 4128 23796 4168
rect 23768 4100 24256 4128
rect 15933 4063 15991 4069
rect 15933 4060 15945 4063
rect 15620 4032 15945 4060
rect 15620 4020 15626 4032
rect 15933 4029 15945 4032
rect 15979 4029 15991 4063
rect 15933 4023 15991 4029
rect 16117 4063 16175 4069
rect 16117 4029 16129 4063
rect 16163 4029 16175 4063
rect 16117 4023 16175 4029
rect 16209 4063 16267 4069
rect 16209 4029 16221 4063
rect 16255 4029 16267 4063
rect 16209 4023 16267 4029
rect 16301 4063 16359 4069
rect 16301 4029 16313 4063
rect 16347 4029 16359 4063
rect 16301 4023 16359 4029
rect 14369 3995 14427 4001
rect 14369 3992 14381 3995
rect 12406 3964 14381 3992
rect 11302 3955 11360 3961
rect 14369 3961 14381 3964
rect 14415 3961 14427 3995
rect 14369 3955 14427 3961
rect 14737 3995 14795 4001
rect 14737 3961 14749 3995
rect 14783 3992 14795 3995
rect 16132 3992 16160 4023
rect 14783 3964 16160 3992
rect 16316 3992 16344 4023
rect 16482 4020 16488 4072
rect 16540 4060 16546 4072
rect 16669 4063 16727 4069
rect 16669 4060 16681 4063
rect 16540 4032 16681 4060
rect 16540 4020 16546 4032
rect 16669 4029 16681 4032
rect 16715 4060 16727 4063
rect 18506 4060 18512 4072
rect 16715 4032 18512 4060
rect 16715 4029 16727 4032
rect 16669 4023 16727 4029
rect 18506 4020 18512 4032
rect 18564 4060 18570 4072
rect 21082 4069 21088 4072
rect 18969 4063 19027 4069
rect 18969 4060 18981 4063
rect 18564 4032 18981 4060
rect 18564 4020 18570 4032
rect 18969 4029 18981 4032
rect 19015 4029 19027 4063
rect 21076 4060 21088 4069
rect 21043 4032 21088 4060
rect 18969 4023 19027 4029
rect 21076 4023 21088 4032
rect 21082 4020 21088 4023
rect 21140 4020 21146 4072
rect 22186 4020 22192 4072
rect 22244 4060 22250 4072
rect 22554 4069 22560 4072
rect 22373 4063 22431 4069
rect 22373 4060 22385 4063
rect 22244 4032 22385 4060
rect 22244 4020 22250 4032
rect 22373 4029 22385 4032
rect 22419 4029 22431 4063
rect 22373 4023 22431 4029
rect 22521 4063 22560 4069
rect 22521 4029 22533 4063
rect 22521 4023 22560 4029
rect 22554 4020 22560 4023
rect 22612 4020 22618 4072
rect 22830 4020 22836 4072
rect 22888 4069 22894 4072
rect 22888 4060 22896 4069
rect 22888 4032 22933 4060
rect 22888 4023 22896 4032
rect 22888 4020 22894 4023
rect 23014 4020 23020 4072
rect 23072 4060 23078 4072
rect 23109 4063 23167 4069
rect 23109 4060 23121 4063
rect 23072 4032 23121 4060
rect 23072 4020 23078 4032
rect 23109 4029 23121 4032
rect 23155 4029 23167 4063
rect 23109 4023 23167 4029
rect 23290 4020 23296 4072
rect 23348 4060 23354 4072
rect 23983 4063 24041 4069
rect 23983 4060 23995 4063
rect 23348 4032 23995 4060
rect 23348 4020 23354 4032
rect 23983 4029 23995 4032
rect 24029 4029 24041 4063
rect 23983 4023 24041 4029
rect 24118 4020 24124 4072
rect 24176 4020 24182 4072
rect 24228 4069 24256 4100
rect 24213 4063 24271 4069
rect 24213 4029 24225 4063
rect 24259 4029 24271 4063
rect 24213 4023 24271 4029
rect 24302 4020 24308 4072
rect 24360 4069 24366 4072
rect 24360 4063 24399 4069
rect 24387 4029 24399 4063
rect 24360 4023 24399 4029
rect 24489 4063 24547 4069
rect 24489 4029 24501 4063
rect 24535 4029 24547 4063
rect 24489 4023 24547 4029
rect 24360 4020 24366 4023
rect 16758 3992 16764 4004
rect 16316 3964 16764 3992
rect 14783 3961 14795 3964
rect 14737 3955 14795 3961
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 16936 3995 16994 4001
rect 16936 3961 16948 3995
rect 16982 3992 16994 3995
rect 17586 3992 17592 4004
rect 16982 3964 17592 3992
rect 16982 3961 16994 3964
rect 16936 3955 16994 3961
rect 17586 3952 17592 3964
rect 17644 3952 17650 4004
rect 19058 3952 19064 4004
rect 19116 3992 19122 4004
rect 19214 3995 19272 4001
rect 19214 3992 19226 3995
rect 19116 3964 19226 3992
rect 19116 3952 19122 3964
rect 19214 3961 19226 3964
rect 19260 3961 19272 3995
rect 19214 3955 19272 3961
rect 22646 3952 22652 4004
rect 22704 3952 22710 4004
rect 22741 3995 22799 4001
rect 22741 3961 22753 3995
rect 22787 3961 22799 3995
rect 22741 3955 22799 3961
rect 11011 3896 11192 3924
rect 12621 3927 12679 3933
rect 11011 3893 11023 3896
rect 10965 3887 11023 3893
rect 12621 3893 12633 3927
rect 12667 3924 12679 3927
rect 13170 3924 13176 3936
rect 12667 3896 13176 3924
rect 12667 3893 12679 3896
rect 12621 3887 12679 3893
rect 8628 3884 8634 3887
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 14918 3884 14924 3936
rect 14976 3924 14982 3936
rect 15470 3924 15476 3936
rect 14976 3896 15476 3924
rect 14976 3884 14982 3896
rect 15470 3884 15476 3896
rect 15528 3884 15534 3936
rect 16577 3927 16635 3933
rect 16577 3893 16589 3927
rect 16623 3924 16635 3927
rect 17954 3924 17960 3936
rect 16623 3896 17960 3924
rect 16623 3893 16635 3896
rect 16577 3887 16635 3893
rect 17954 3884 17960 3896
rect 18012 3884 18018 3936
rect 18049 3927 18107 3933
rect 18049 3893 18061 3927
rect 18095 3924 18107 3927
rect 18138 3924 18144 3936
rect 18095 3896 18144 3924
rect 18095 3893 18107 3896
rect 18049 3887 18107 3893
rect 18138 3884 18144 3896
rect 18196 3924 18202 3936
rect 20070 3924 20076 3936
rect 18196 3896 20076 3924
rect 18196 3884 18202 3896
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20254 3884 20260 3936
rect 20312 3924 20318 3936
rect 20349 3927 20407 3933
rect 20349 3924 20361 3927
rect 20312 3896 20361 3924
rect 20312 3884 20318 3896
rect 20349 3893 20361 3896
rect 20395 3924 20407 3927
rect 22756 3924 22784 3955
rect 20395 3896 22784 3924
rect 23017 3927 23075 3933
rect 20395 3893 20407 3896
rect 20349 3887 20407 3893
rect 23017 3893 23029 3927
rect 23063 3924 23075 3927
rect 23198 3924 23204 3936
rect 23063 3896 23204 3924
rect 23063 3893 23075 3896
rect 23017 3887 23075 3893
rect 23198 3884 23204 3896
rect 23256 3884 23262 3936
rect 23382 3884 23388 3936
rect 23440 3924 23446 3936
rect 23845 3927 23903 3933
rect 23845 3924 23857 3927
rect 23440 3896 23857 3924
rect 23440 3884 23446 3896
rect 23845 3893 23857 3896
rect 23891 3893 23903 3927
rect 23845 3887 23903 3893
rect 24394 3884 24400 3936
rect 24452 3924 24458 3936
rect 24504 3924 24532 4023
rect 25130 4020 25136 4072
rect 25188 4020 25194 4072
rect 24452 3896 24532 3924
rect 24581 3927 24639 3933
rect 24452 3884 24458 3896
rect 24581 3893 24593 3927
rect 24627 3924 24639 3927
rect 24670 3924 24676 3936
rect 24627 3896 24676 3924
rect 24627 3893 24639 3896
rect 24581 3887 24639 3893
rect 24670 3884 24676 3896
rect 24728 3884 24734 3936
rect 552 3834 27576 3856
rect 552 3782 7114 3834
rect 7166 3782 7178 3834
rect 7230 3782 7242 3834
rect 7294 3782 7306 3834
rect 7358 3782 7370 3834
rect 7422 3782 13830 3834
rect 13882 3782 13894 3834
rect 13946 3782 13958 3834
rect 14010 3782 14022 3834
rect 14074 3782 14086 3834
rect 14138 3782 20546 3834
rect 20598 3782 20610 3834
rect 20662 3782 20674 3834
rect 20726 3782 20738 3834
rect 20790 3782 20802 3834
rect 20854 3782 27262 3834
rect 27314 3782 27326 3834
rect 27378 3782 27390 3834
rect 27442 3782 27454 3834
rect 27506 3782 27518 3834
rect 27570 3782 27576 3834
rect 552 3760 27576 3782
rect 5258 3680 5264 3732
rect 5316 3720 5322 3732
rect 5353 3723 5411 3729
rect 5353 3720 5365 3723
rect 5316 3692 5365 3720
rect 5316 3680 5322 3692
rect 5353 3689 5365 3692
rect 5399 3689 5411 3723
rect 6270 3720 6276 3732
rect 5353 3683 5411 3689
rect 5552 3692 6276 3720
rect 5552 3593 5580 3692
rect 6270 3680 6276 3692
rect 6328 3720 6334 3732
rect 6328 3692 7604 3720
rect 6328 3680 6334 3692
rect 7576 3664 7604 3692
rect 8294 3680 8300 3732
rect 8352 3680 8358 3732
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 12308 3692 13308 3720
rect 12308 3680 12314 3692
rect 7098 3661 7104 3664
rect 7092 3615 7104 3661
rect 7156 3652 7162 3664
rect 7156 3624 7192 3652
rect 7098 3612 7104 3615
rect 7156 3612 7162 3624
rect 7558 3612 7564 3664
rect 7616 3652 7622 3664
rect 8662 3652 8668 3664
rect 7616 3624 8668 3652
rect 7616 3612 7622 3624
rect 8662 3612 8668 3624
rect 8720 3612 8726 3664
rect 12986 3652 12992 3664
rect 8956 3624 12992 3652
rect 5537 3587 5595 3593
rect 5537 3553 5549 3587
rect 5583 3553 5595 3587
rect 5537 3547 5595 3553
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3584 5687 3587
rect 5813 3587 5871 3593
rect 5813 3584 5825 3587
rect 5675 3556 5825 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 5813 3553 5825 3556
rect 5859 3553 5871 3587
rect 5813 3547 5871 3553
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3584 6515 3587
rect 6546 3584 6552 3596
rect 6503 3556 6552 3584
rect 6503 3553 6515 3556
rect 6457 3547 6515 3553
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 8202 3544 8208 3596
rect 8260 3584 8266 3596
rect 8956 3593 8984 3624
rect 12986 3612 12992 3624
rect 13044 3612 13050 3664
rect 13170 3612 13176 3664
rect 13228 3612 13234 3664
rect 13280 3661 13308 3692
rect 15378 3680 15384 3732
rect 15436 3720 15442 3732
rect 15436 3692 15608 3720
rect 15436 3680 15442 3692
rect 13265 3655 13323 3661
rect 13265 3621 13277 3655
rect 13311 3621 13323 3655
rect 13265 3615 13323 3621
rect 15197 3655 15255 3661
rect 15197 3621 15209 3655
rect 15243 3652 15255 3655
rect 15243 3624 15516 3652
rect 15243 3621 15255 3624
rect 15197 3615 15255 3621
rect 8941 3587 8999 3593
rect 8941 3584 8953 3587
rect 8260 3556 8953 3584
rect 8260 3544 8266 3556
rect 8941 3553 8953 3556
rect 8987 3553 8999 3587
rect 8941 3547 8999 3553
rect 9950 3544 9956 3596
rect 10008 3544 10014 3596
rect 11517 3587 11575 3593
rect 11517 3553 11529 3587
rect 11563 3584 11575 3587
rect 11606 3584 11612 3596
rect 11563 3556 11612 3584
rect 11563 3553 11575 3556
rect 11517 3547 11575 3553
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 11784 3587 11842 3593
rect 11784 3553 11796 3587
rect 11830 3584 11842 3587
rect 13081 3587 13139 3593
rect 11830 3556 13032 3584
rect 11830 3553 11842 3556
rect 11784 3547 11842 3553
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 5399 3488 5672 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 5644 3460 5672 3488
rect 6822 3476 6828 3528
rect 6880 3476 6886 3528
rect 13004 3525 13032 3556
rect 13081 3553 13093 3587
rect 13127 3584 13139 3587
rect 13127 3556 13308 3584
rect 13127 3553 13139 3556
rect 13081 3547 13139 3553
rect 13280 3528 13308 3556
rect 13446 3544 13452 3596
rect 13504 3544 13510 3596
rect 13538 3544 13544 3596
rect 13596 3544 13602 3596
rect 14182 3544 14188 3596
rect 14240 3584 14246 3596
rect 14734 3584 14740 3596
rect 14240 3556 14740 3584
rect 14240 3544 14246 3556
rect 14734 3544 14740 3556
rect 14792 3544 14798 3596
rect 14829 3587 14887 3593
rect 14829 3553 14841 3587
rect 14875 3553 14887 3587
rect 14829 3547 14887 3553
rect 9033 3519 9091 3525
rect 9033 3485 9045 3519
rect 9079 3516 9091 3519
rect 10137 3519 10195 3525
rect 10137 3516 10149 3519
rect 9079 3488 10149 3516
rect 9079 3485 9091 3488
rect 9033 3479 9091 3485
rect 10137 3485 10149 3488
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 5626 3408 5632 3460
rect 5684 3408 5690 3460
rect 8205 3451 8263 3457
rect 8205 3417 8217 3451
rect 8251 3448 8263 3451
rect 9048 3448 9076 3479
rect 13262 3476 13268 3528
rect 13320 3476 13326 3528
rect 8251 3420 9076 3448
rect 8251 3417 8263 3420
rect 8205 3411 8263 3417
rect 9674 3408 9680 3460
rect 9732 3448 9738 3460
rect 14844 3448 14872 3547
rect 15010 3544 15016 3596
rect 15068 3544 15074 3596
rect 15286 3544 15292 3596
rect 15344 3544 15350 3596
rect 15488 3593 15516 3624
rect 15580 3593 15608 3692
rect 17586 3680 17592 3732
rect 17644 3680 17650 3732
rect 18414 3680 18420 3732
rect 18472 3680 18478 3732
rect 19058 3680 19064 3732
rect 19116 3680 19122 3732
rect 22649 3723 22707 3729
rect 22649 3689 22661 3723
rect 22695 3720 22707 3723
rect 25130 3720 25136 3732
rect 22695 3692 25136 3720
rect 22695 3689 22707 3692
rect 22649 3683 22707 3689
rect 25130 3680 25136 3692
rect 25188 3680 25194 3732
rect 25590 3680 25596 3732
rect 25648 3680 25654 3732
rect 16482 3652 16488 3664
rect 16132 3624 16488 3652
rect 15473 3587 15531 3593
rect 15473 3553 15485 3587
rect 15519 3553 15531 3587
rect 15473 3547 15531 3553
rect 15565 3587 15623 3593
rect 15565 3553 15577 3587
rect 15611 3553 15623 3587
rect 15565 3547 15623 3553
rect 15654 3544 15660 3596
rect 15712 3544 15718 3596
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 16132 3593 16160 3624
rect 16482 3612 16488 3624
rect 16540 3612 16546 3664
rect 18046 3612 18052 3664
rect 18104 3652 18110 3664
rect 18432 3652 18460 3680
rect 23382 3652 23388 3664
rect 18104 3624 18736 3652
rect 18104 3612 18110 3624
rect 16117 3587 16175 3593
rect 16117 3584 16129 3587
rect 16080 3556 16129 3584
rect 16080 3544 16086 3556
rect 16117 3553 16129 3556
rect 16163 3553 16175 3587
rect 16373 3587 16431 3593
rect 16373 3584 16385 3587
rect 16117 3547 16175 3553
rect 16224 3556 16385 3584
rect 15933 3519 15991 3525
rect 15933 3485 15945 3519
rect 15979 3516 15991 3519
rect 16224 3516 16252 3556
rect 16373 3553 16385 3556
rect 16419 3553 16431 3587
rect 16373 3547 16431 3553
rect 17954 3544 17960 3596
rect 18012 3584 18018 3596
rect 18141 3587 18199 3593
rect 18141 3584 18153 3587
rect 18012 3556 18153 3584
rect 18012 3544 18018 3556
rect 18141 3553 18153 3556
rect 18187 3553 18199 3587
rect 18141 3547 18199 3553
rect 18417 3587 18475 3593
rect 18417 3553 18429 3587
rect 18463 3553 18475 3587
rect 18417 3547 18475 3553
rect 15979 3488 16252 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 18432 3516 18460 3547
rect 18598 3544 18604 3596
rect 18656 3544 18662 3596
rect 18708 3593 18736 3624
rect 22204 3624 23388 3652
rect 18693 3587 18751 3593
rect 18693 3553 18705 3587
rect 18739 3553 18751 3587
rect 18693 3547 18751 3553
rect 18785 3587 18843 3593
rect 18785 3553 18797 3587
rect 18831 3584 18843 3587
rect 19613 3587 19671 3593
rect 19613 3584 19625 3587
rect 18831 3556 19625 3584
rect 18831 3553 18843 3556
rect 18785 3547 18843 3553
rect 19613 3553 19625 3556
rect 19659 3553 19671 3587
rect 19613 3547 19671 3553
rect 20254 3544 20260 3596
rect 20312 3544 20318 3596
rect 21542 3544 21548 3596
rect 21600 3544 21606 3596
rect 21637 3587 21695 3593
rect 21637 3553 21649 3587
rect 21683 3553 21695 3587
rect 21637 3547 21695 3553
rect 17920 3488 18460 3516
rect 20993 3519 21051 3525
rect 17920 3476 17926 3488
rect 20993 3485 21005 3519
rect 21039 3516 21051 3519
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 21039 3488 21281 3516
rect 21039 3485 21051 3488
rect 20993 3479 21051 3485
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21652 3516 21680 3547
rect 21726 3544 21732 3596
rect 21784 3544 21790 3596
rect 21910 3544 21916 3596
rect 21968 3584 21974 3596
rect 22204 3593 22232 3624
rect 23382 3612 23388 3624
rect 23440 3612 23446 3664
rect 23876 3655 23934 3661
rect 23876 3621 23888 3655
rect 23922 3652 23934 3655
rect 24670 3652 24676 3664
rect 23922 3624 24676 3652
rect 23922 3621 23934 3624
rect 23876 3615 23934 3621
rect 24670 3612 24676 3624
rect 24728 3612 24734 3664
rect 22005 3587 22063 3593
rect 22005 3584 22017 3587
rect 21968 3556 22017 3584
rect 21968 3544 21974 3556
rect 22005 3553 22017 3556
rect 22051 3553 22063 3587
rect 22005 3547 22063 3553
rect 22189 3587 22247 3593
rect 22189 3553 22201 3587
rect 22235 3553 22247 3587
rect 22189 3547 22247 3553
rect 22281 3587 22339 3593
rect 22281 3553 22293 3587
rect 22327 3553 22339 3587
rect 22281 3547 22339 3553
rect 22296 3516 22324 3547
rect 22370 3544 22376 3596
rect 22428 3544 22434 3596
rect 24486 3593 24492 3596
rect 24480 3547 24492 3593
rect 24486 3544 24492 3547
rect 24544 3544 24550 3596
rect 22462 3516 22468 3528
rect 21652 3488 22468 3516
rect 21269 3479 21327 3485
rect 22462 3476 22468 3488
rect 22520 3516 22526 3528
rect 23106 3516 23112 3528
rect 22520 3488 23112 3516
rect 22520 3476 22526 3488
rect 23106 3476 23112 3488
rect 23164 3476 23170 3528
rect 24121 3519 24179 3525
rect 24121 3485 24133 3519
rect 24167 3485 24179 3519
rect 24121 3479 24179 3485
rect 24213 3519 24271 3525
rect 24213 3485 24225 3519
rect 24259 3485 24271 3519
rect 24213 3479 24271 3485
rect 9732 3420 10272 3448
rect 9732 3408 9738 3420
rect 7742 3340 7748 3392
rect 7800 3380 7806 3392
rect 9769 3383 9827 3389
rect 9769 3380 9781 3383
rect 7800 3352 9781 3380
rect 7800 3340 7806 3352
rect 9769 3349 9781 3352
rect 9815 3349 9827 3383
rect 10244 3380 10272 3420
rect 12820 3420 14872 3448
rect 12820 3380 12848 3420
rect 21818 3408 21824 3460
rect 21876 3448 21882 3460
rect 22741 3451 22799 3457
rect 22741 3448 22753 3451
rect 21876 3420 22753 3448
rect 21876 3408 21882 3420
rect 22741 3417 22753 3420
rect 22787 3417 22799 3451
rect 22741 3411 22799 3417
rect 24136 3448 24164 3479
rect 24219 3448 24247 3479
rect 24136 3420 24247 3448
rect 10244 3352 12848 3380
rect 9769 3343 9827 3349
rect 12894 3340 12900 3392
rect 12952 3380 12958 3392
rect 13630 3380 13636 3392
rect 12952 3352 13636 3380
rect 12952 3340 12958 3352
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 17497 3383 17555 3389
rect 17497 3349 17509 3383
rect 17543 3380 17555 3383
rect 18046 3380 18052 3392
rect 17543 3352 18052 3380
rect 17543 3349 17555 3352
rect 17497 3343 17555 3349
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 20346 3340 20352 3392
rect 20404 3340 20410 3392
rect 21910 3340 21916 3392
rect 21968 3380 21974 3392
rect 22278 3380 22284 3392
rect 21968 3352 22284 3380
rect 21968 3340 21974 3352
rect 22278 3340 22284 3352
rect 22336 3340 22342 3392
rect 23750 3340 23756 3392
rect 23808 3380 23814 3392
rect 24136 3380 24164 3420
rect 23808 3352 24164 3380
rect 23808 3340 23814 3352
rect 552 3290 27416 3312
rect 552 3238 3756 3290
rect 3808 3238 3820 3290
rect 3872 3238 3884 3290
rect 3936 3238 3948 3290
rect 4000 3238 4012 3290
rect 4064 3238 10472 3290
rect 10524 3238 10536 3290
rect 10588 3238 10600 3290
rect 10652 3238 10664 3290
rect 10716 3238 10728 3290
rect 10780 3238 17188 3290
rect 17240 3238 17252 3290
rect 17304 3238 17316 3290
rect 17368 3238 17380 3290
rect 17432 3238 17444 3290
rect 17496 3238 23904 3290
rect 23956 3238 23968 3290
rect 24020 3238 24032 3290
rect 24084 3238 24096 3290
rect 24148 3238 24160 3290
rect 24212 3238 27416 3290
rect 552 3216 27416 3238
rect 6362 3136 6368 3188
rect 6420 3136 6426 3188
rect 8570 3176 8576 3188
rect 6564 3148 8576 3176
rect 6454 3068 6460 3120
rect 6512 3068 6518 3120
rect 2590 3000 2596 3052
rect 2648 3040 2654 3052
rect 4522 3040 4528 3052
rect 2648 3012 4528 3040
rect 2648 3000 2654 3012
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3040 6423 3043
rect 6472 3040 6500 3068
rect 6411 3012 6500 3040
rect 6411 3009 6423 3012
rect 6365 3003 6423 3009
rect 6457 2975 6515 2981
rect 6457 2941 6469 2975
rect 6503 2941 6515 2975
rect 6457 2935 6515 2941
rect 6472 2836 6500 2935
rect 6564 2904 6592 3148
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8662 3136 8668 3188
rect 8720 3176 8726 3188
rect 8941 3179 8999 3185
rect 8941 3176 8953 3179
rect 8720 3148 8953 3176
rect 8720 3136 8726 3148
rect 8941 3145 8953 3148
rect 8987 3145 8999 3179
rect 8941 3139 8999 3145
rect 11790 3136 11796 3188
rect 11848 3136 11854 3188
rect 12434 3136 12440 3188
rect 12492 3136 12498 3188
rect 12986 3136 12992 3188
rect 13044 3176 13050 3188
rect 14182 3176 14188 3188
rect 13044 3148 14188 3176
rect 13044 3136 13050 3148
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 15654 3136 15660 3188
rect 15712 3176 15718 3188
rect 16669 3179 16727 3185
rect 16669 3176 16681 3179
rect 15712 3148 16681 3176
rect 15712 3136 15718 3148
rect 16669 3145 16681 3148
rect 16715 3145 16727 3179
rect 16669 3139 16727 3145
rect 16758 3136 16764 3188
rect 16816 3176 16822 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 16816 3148 17417 3176
rect 16816 3136 16822 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17405 3139 17463 3145
rect 21361 3179 21419 3185
rect 21361 3145 21373 3179
rect 21407 3176 21419 3179
rect 21542 3176 21548 3188
rect 21407 3148 21548 3176
rect 21407 3145 21419 3148
rect 21361 3139 21419 3145
rect 21542 3136 21548 3148
rect 21600 3136 21606 3188
rect 21634 3136 21640 3188
rect 21692 3176 21698 3188
rect 21692 3148 22048 3176
rect 21692 3136 21698 3148
rect 22020 3120 22048 3148
rect 22370 3136 22376 3188
rect 22428 3176 22434 3188
rect 22649 3179 22707 3185
rect 22649 3176 22661 3179
rect 22428 3148 22661 3176
rect 22428 3136 22434 3148
rect 22649 3145 22661 3148
rect 22695 3145 22707 3179
rect 22649 3139 22707 3145
rect 23290 3136 23296 3188
rect 23348 3176 23354 3188
rect 23348 3148 24164 3176
rect 23348 3136 23354 3148
rect 8202 3068 8208 3120
rect 8260 3068 8266 3120
rect 11609 3111 11667 3117
rect 11609 3077 11621 3111
rect 11655 3108 11667 3111
rect 13173 3111 13231 3117
rect 13173 3108 13185 3111
rect 11655 3080 13185 3108
rect 11655 3077 11667 3080
rect 11609 3071 11667 3077
rect 13173 3077 13185 3080
rect 13219 3108 13231 3111
rect 13446 3108 13452 3120
rect 13219 3080 13452 3108
rect 13219 3077 13231 3080
rect 13173 3071 13231 3077
rect 13446 3068 13452 3080
rect 13504 3068 13510 3120
rect 21269 3111 21327 3117
rect 21269 3077 21281 3111
rect 21315 3108 21327 3111
rect 21315 3080 21956 3108
rect 21315 3077 21327 3080
rect 21269 3071 21327 3077
rect 6822 3000 6828 3052
rect 6880 3000 6886 3052
rect 12345 3043 12403 3049
rect 12345 3009 12357 3043
rect 12391 3040 12403 3043
rect 12526 3040 12532 3052
rect 12391 3012 12532 3040
rect 12391 3009 12403 3012
rect 12345 3003 12403 3009
rect 12526 3000 12532 3012
rect 12584 3040 12590 3052
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 12584 3012 12909 3040
rect 12584 3000 12590 3012
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13354 3000 13360 3052
rect 13412 3000 13418 3052
rect 17313 3043 17371 3049
rect 17313 3009 17325 3043
rect 17359 3040 17371 3043
rect 18046 3040 18052 3052
rect 17359 3012 18052 3040
rect 17359 3009 17371 3012
rect 17313 3003 17371 3009
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 21928 3049 21956 3080
rect 22002 3068 22008 3120
rect 22060 3108 22066 3120
rect 24136 3108 24164 3148
rect 24486 3136 24492 3188
rect 24544 3176 24550 3188
rect 24581 3179 24639 3185
rect 24581 3176 24593 3179
rect 24544 3148 24593 3176
rect 24544 3136 24550 3148
rect 24581 3145 24593 3148
rect 24627 3145 24639 3179
rect 24581 3139 24639 3145
rect 25590 3108 25596 3120
rect 22060 3080 23888 3108
rect 22060 3068 22066 3080
rect 21913 3043 21971 3049
rect 21913 3009 21925 3043
rect 21959 3040 21971 3043
rect 22462 3040 22468 3052
rect 21959 3012 22468 3040
rect 21959 3009 21971 3012
rect 21913 3003 21971 3009
rect 22462 3000 22468 3012
rect 22520 3000 22526 3052
rect 6641 2975 6699 2981
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 8481 2975 8539 2981
rect 8481 2972 8493 2975
rect 6687 2944 8493 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 8481 2941 8493 2944
rect 8527 2941 8539 2975
rect 8481 2935 8539 2941
rect 8573 2975 8631 2981
rect 8573 2941 8585 2975
rect 8619 2972 8631 2975
rect 9674 2972 9680 2984
rect 8619 2944 9680 2972
rect 8619 2941 8631 2944
rect 8573 2935 8631 2941
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 11333 2975 11391 2981
rect 11333 2941 11345 2975
rect 11379 2941 11391 2975
rect 11333 2935 11391 2941
rect 6733 2907 6791 2913
rect 6733 2904 6745 2907
rect 6564 2876 6745 2904
rect 6733 2873 6745 2876
rect 6779 2873 6791 2907
rect 6733 2867 6791 2873
rect 7092 2907 7150 2913
rect 7092 2873 7104 2907
rect 7138 2904 7150 2907
rect 7558 2904 7564 2916
rect 7138 2876 7564 2904
rect 7138 2873 7150 2876
rect 7092 2867 7150 2873
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 7742 2864 7748 2916
rect 7800 2904 7806 2916
rect 8909 2907 8967 2913
rect 8909 2904 8921 2907
rect 7800 2876 8921 2904
rect 7800 2864 7806 2876
rect 8909 2873 8921 2876
rect 8955 2873 8967 2907
rect 8909 2867 8967 2873
rect 9122 2864 9128 2916
rect 9180 2864 9186 2916
rect 11348 2848 11376 2935
rect 11422 2932 11428 2984
rect 11480 2932 11486 2984
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2972 12035 2975
rect 12250 2972 12256 2984
rect 12023 2944 12256 2972
rect 12023 2941 12035 2944
rect 11977 2935 12035 2941
rect 12250 2932 12256 2944
rect 12308 2972 12314 2984
rect 12621 2975 12679 2981
rect 12621 2972 12633 2975
rect 12308 2944 12633 2972
rect 12308 2932 12314 2944
rect 12621 2941 12633 2944
rect 12667 2941 12679 2975
rect 12621 2935 12679 2941
rect 12713 2975 12771 2981
rect 12713 2941 12725 2975
rect 12759 2941 12771 2975
rect 12713 2935 12771 2941
rect 12805 2975 12863 2981
rect 12805 2941 12817 2975
rect 12851 2941 12863 2975
rect 12805 2935 12863 2941
rect 11440 2904 11468 2932
rect 12069 2907 12127 2913
rect 12069 2904 12081 2907
rect 11440 2876 12081 2904
rect 12069 2873 12081 2876
rect 12115 2904 12127 2907
rect 12728 2904 12756 2935
rect 12115 2876 12756 2904
rect 12820 2904 12848 2935
rect 12986 2932 12992 2984
rect 13044 2972 13050 2984
rect 13081 2975 13139 2981
rect 13081 2972 13093 2975
rect 13044 2944 13093 2972
rect 13044 2932 13050 2944
rect 13081 2941 13093 2944
rect 13127 2941 13139 2975
rect 13081 2935 13139 2941
rect 15286 2932 15292 2984
rect 15344 2972 15350 2984
rect 17862 2972 17868 2984
rect 15344 2944 17868 2972
rect 15344 2932 15350 2944
rect 17862 2932 17868 2944
rect 17920 2932 17926 2984
rect 17957 2975 18015 2981
rect 17957 2941 17969 2975
rect 18003 2972 18015 2975
rect 18138 2972 18144 2984
rect 18003 2944 18144 2972
rect 18003 2941 18015 2944
rect 17957 2935 18015 2941
rect 18138 2932 18144 2944
rect 18196 2932 18202 2984
rect 18414 2932 18420 2984
rect 18472 2932 18478 2984
rect 18690 2932 18696 2984
rect 18748 2932 18754 2984
rect 19889 2975 19947 2981
rect 19889 2941 19901 2975
rect 19935 2972 19947 2975
rect 19978 2972 19984 2984
rect 19935 2944 19984 2972
rect 19935 2941 19947 2944
rect 19889 2935 19947 2941
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 21818 2932 21824 2984
rect 21876 2972 21882 2984
rect 23860 2981 23888 3080
rect 24136 3080 25596 3108
rect 23201 2975 23259 2981
rect 23201 2972 23213 2975
rect 21876 2944 23213 2972
rect 21876 2932 21882 2944
rect 23201 2941 23213 2944
rect 23247 2941 23259 2975
rect 23201 2935 23259 2941
rect 23845 2975 23903 2981
rect 23845 2941 23857 2975
rect 23891 2941 23903 2975
rect 23845 2935 23903 2941
rect 20156 2907 20214 2913
rect 12820 2876 13216 2904
rect 12115 2873 12127 2876
rect 12069 2867 12127 2873
rect 8110 2836 8116 2848
rect 6472 2808 8116 2836
rect 8110 2796 8116 2808
rect 8168 2836 8174 2848
rect 8757 2839 8815 2845
rect 8757 2836 8769 2839
rect 8168 2808 8769 2836
rect 8168 2796 8174 2808
rect 8757 2805 8769 2808
rect 8803 2805 8815 2839
rect 8757 2799 8815 2805
rect 10042 2796 10048 2848
rect 10100 2836 10106 2848
rect 11330 2836 11336 2848
rect 10100 2808 11336 2836
rect 10100 2796 10106 2808
rect 11330 2796 11336 2808
rect 11388 2836 11394 2848
rect 12161 2839 12219 2845
rect 12161 2836 12173 2839
rect 11388 2808 12173 2836
rect 11388 2796 11394 2808
rect 12161 2805 12173 2808
rect 12207 2836 12219 2839
rect 12820 2836 12848 2876
rect 13188 2848 13216 2876
rect 20156 2873 20168 2907
rect 20202 2904 20214 2907
rect 20346 2904 20352 2916
rect 20202 2876 20352 2904
rect 20202 2873 20214 2876
rect 20156 2867 20214 2873
rect 20346 2864 20352 2876
rect 20404 2864 20410 2916
rect 23860 2904 23888 2935
rect 24026 2932 24032 2984
rect 24084 2932 24090 2984
rect 24136 2981 24164 3080
rect 25590 3068 25596 3080
rect 25648 3068 25654 3120
rect 24489 3043 24547 3049
rect 24489 3009 24501 3043
rect 24535 3040 24547 3043
rect 25133 3043 25191 3049
rect 25133 3040 25145 3043
rect 24535 3012 25145 3040
rect 24535 3009 24547 3012
rect 24489 3003 24547 3009
rect 25133 3009 25145 3012
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 25682 3000 25688 3052
rect 25740 3040 25746 3052
rect 25869 3043 25927 3049
rect 25869 3040 25881 3043
rect 25740 3012 25881 3040
rect 25740 3000 25746 3012
rect 25869 3009 25881 3012
rect 25915 3009 25927 3043
rect 25869 3003 25927 3009
rect 24121 2975 24179 2981
rect 24121 2941 24133 2975
rect 24167 2941 24179 2975
rect 24121 2935 24179 2941
rect 24213 2975 24271 2981
rect 24213 2941 24225 2975
rect 24259 2972 24271 2975
rect 25317 2975 25375 2981
rect 25317 2972 25329 2975
rect 24259 2944 25329 2972
rect 24259 2941 24271 2944
rect 24213 2935 24271 2941
rect 25317 2941 25329 2944
rect 25363 2941 25375 2975
rect 25317 2935 25375 2941
rect 25222 2904 25228 2916
rect 23860 2876 25228 2904
rect 25222 2864 25228 2876
rect 25280 2864 25286 2916
rect 12207 2808 12848 2836
rect 12207 2805 12219 2808
rect 12161 2799 12219 2805
rect 13170 2796 13176 2848
rect 13228 2796 13234 2848
rect 13357 2839 13415 2845
rect 13357 2805 13369 2839
rect 13403 2836 13415 2839
rect 13722 2836 13728 2848
rect 13403 2808 13728 2836
rect 13403 2805 13415 2808
rect 13357 2799 13415 2805
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 16114 2836 16120 2848
rect 15252 2808 16120 2836
rect 15252 2796 15258 2808
rect 16114 2796 16120 2808
rect 16172 2796 16178 2848
rect 17218 2796 17224 2848
rect 17276 2836 17282 2848
rect 18233 2839 18291 2845
rect 18233 2836 18245 2839
rect 17276 2808 18245 2836
rect 17276 2796 17282 2808
rect 18233 2805 18245 2808
rect 18279 2805 18291 2839
rect 18233 2799 18291 2805
rect 19334 2796 19340 2848
rect 19392 2796 19398 2848
rect 21450 2796 21456 2848
rect 21508 2836 21514 2848
rect 22186 2836 22192 2848
rect 21508 2808 22192 2836
rect 21508 2796 21514 2808
rect 22186 2796 22192 2808
rect 22244 2836 22250 2848
rect 22830 2836 22836 2848
rect 22244 2808 22836 2836
rect 22244 2796 22250 2808
rect 22830 2796 22836 2808
rect 22888 2836 22894 2848
rect 23198 2836 23204 2848
rect 22888 2808 23204 2836
rect 22888 2796 22894 2808
rect 23198 2796 23204 2808
rect 23256 2796 23262 2848
rect 23382 2796 23388 2848
rect 23440 2836 23446 2848
rect 24486 2836 24492 2848
rect 23440 2808 24492 2836
rect 23440 2796 23446 2808
rect 24486 2796 24492 2808
rect 24544 2796 24550 2848
rect 552 2746 27576 2768
rect 552 2694 7114 2746
rect 7166 2694 7178 2746
rect 7230 2694 7242 2746
rect 7294 2694 7306 2746
rect 7358 2694 7370 2746
rect 7422 2694 13830 2746
rect 13882 2694 13894 2746
rect 13946 2694 13958 2746
rect 14010 2694 14022 2746
rect 14074 2694 14086 2746
rect 14138 2694 20546 2746
rect 20598 2694 20610 2746
rect 20662 2694 20674 2746
rect 20726 2694 20738 2746
rect 20790 2694 20802 2746
rect 20854 2694 27262 2746
rect 27314 2694 27326 2746
rect 27378 2694 27390 2746
rect 27442 2694 27454 2746
rect 27506 2694 27518 2746
rect 27570 2694 27576 2746
rect 552 2672 27576 2694
rect 7558 2592 7564 2644
rect 7616 2592 7622 2644
rect 11238 2632 11244 2644
rect 10244 2604 11244 2632
rect 9953 2567 10011 2573
rect 9953 2564 9965 2567
rect 7484 2536 9965 2564
rect 7484 2508 7512 2536
rect 9953 2533 9965 2536
rect 9999 2564 10011 2567
rect 10244 2564 10272 2604
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 11333 2635 11391 2641
rect 11333 2601 11345 2635
rect 11379 2632 11391 2635
rect 11514 2632 11520 2644
rect 11379 2604 11520 2632
rect 11379 2601 11391 2604
rect 11333 2595 11391 2601
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 11977 2635 12035 2641
rect 11977 2601 11989 2635
rect 12023 2632 12035 2635
rect 12250 2632 12256 2644
rect 12023 2604 12256 2632
rect 12023 2601 12035 2604
rect 11977 2595 12035 2601
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 13412 2604 13676 2632
rect 13412 2592 13418 2604
rect 9999 2536 10272 2564
rect 9999 2533 10011 2536
rect 9953 2527 10011 2533
rect 7466 2456 7472 2508
rect 7524 2456 7530 2508
rect 7653 2499 7711 2505
rect 7653 2465 7665 2499
rect 7699 2496 7711 2499
rect 7926 2496 7932 2508
rect 7699 2468 7932 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 7926 2456 7932 2468
rect 7984 2456 7990 2508
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 10042 2496 10048 2508
rect 9815 2468 10048 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 10244 2505 10272 2536
rect 11072 2536 11836 2564
rect 11072 2508 11100 2536
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2465 10287 2499
rect 10229 2459 10287 2465
rect 10413 2499 10471 2505
rect 10413 2465 10425 2499
rect 10459 2496 10471 2499
rect 10459 2468 10640 2496
rect 10459 2465 10471 2468
rect 10413 2459 10471 2465
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2397 10563 2431
rect 10612 2428 10640 2468
rect 11054 2456 11060 2508
rect 11112 2456 11118 2508
rect 11241 2499 11299 2505
rect 11241 2465 11253 2499
rect 11287 2465 11299 2499
rect 11241 2459 11299 2465
rect 10962 2428 10968 2440
rect 10612 2400 10968 2428
rect 10505 2391 10563 2397
rect 10318 2320 10324 2372
rect 10376 2360 10382 2372
rect 10520 2360 10548 2391
rect 10962 2388 10968 2400
rect 11020 2428 11026 2440
rect 11149 2431 11207 2437
rect 11149 2428 11161 2431
rect 11020 2400 11161 2428
rect 11020 2388 11026 2400
rect 11149 2397 11161 2400
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 10376 2332 10548 2360
rect 11256 2360 11284 2459
rect 11422 2456 11428 2508
rect 11480 2496 11486 2508
rect 11808 2505 11836 2536
rect 12526 2524 12532 2576
rect 12584 2524 12590 2576
rect 13262 2524 13268 2576
rect 13320 2564 13326 2576
rect 13509 2567 13567 2573
rect 13509 2564 13521 2567
rect 13320 2536 13521 2564
rect 13320 2524 13326 2536
rect 13509 2533 13521 2536
rect 13555 2533 13567 2567
rect 13648 2564 13676 2604
rect 14182 2592 14188 2644
rect 14240 2632 14246 2644
rect 14829 2635 14887 2641
rect 14829 2632 14841 2635
rect 14240 2604 14841 2632
rect 14240 2592 14246 2604
rect 14829 2601 14841 2604
rect 14875 2601 14887 2635
rect 14829 2595 14887 2601
rect 16114 2592 16120 2644
rect 16172 2632 16178 2644
rect 17218 2632 17224 2644
rect 16172 2604 17224 2632
rect 16172 2592 16178 2604
rect 17218 2592 17224 2604
rect 17276 2592 17282 2644
rect 17862 2632 17868 2644
rect 17512 2604 17868 2632
rect 13725 2567 13783 2573
rect 13725 2564 13737 2567
rect 13648 2536 13737 2564
rect 13509 2527 13567 2533
rect 13725 2533 13737 2536
rect 13771 2533 13783 2567
rect 13725 2527 13783 2533
rect 13817 2567 13875 2573
rect 13817 2533 13829 2567
rect 13863 2564 13875 2567
rect 13906 2564 13912 2576
rect 13863 2536 13912 2564
rect 13863 2533 13875 2536
rect 13817 2527 13875 2533
rect 13906 2524 13912 2536
rect 13964 2524 13970 2576
rect 14274 2524 14280 2576
rect 14332 2564 14338 2576
rect 14332 2536 17356 2564
rect 14332 2524 14338 2536
rect 11517 2499 11575 2505
rect 11517 2496 11529 2499
rect 11480 2468 11529 2496
rect 11480 2456 11486 2468
rect 11517 2465 11529 2468
rect 11563 2465 11575 2499
rect 11517 2459 11575 2465
rect 11793 2499 11851 2505
rect 11793 2465 11805 2499
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 12161 2499 12219 2505
rect 12161 2465 12173 2499
rect 12207 2465 12219 2499
rect 12161 2459 12219 2465
rect 11330 2388 11336 2440
rect 11388 2428 11394 2440
rect 11609 2431 11667 2437
rect 11609 2428 11621 2431
rect 11388 2400 11621 2428
rect 11388 2388 11394 2400
rect 11609 2397 11621 2400
rect 11655 2397 11667 2431
rect 11609 2391 11667 2397
rect 11701 2431 11759 2437
rect 11701 2397 11713 2431
rect 11747 2428 11759 2431
rect 11974 2428 11980 2440
rect 11747 2400 11980 2428
rect 11747 2397 11759 2400
rect 11701 2391 11759 2397
rect 11974 2388 11980 2400
rect 12032 2428 12038 2440
rect 12176 2428 12204 2459
rect 12250 2456 12256 2508
rect 12308 2456 12314 2508
rect 12345 2499 12403 2505
rect 12345 2465 12357 2499
rect 12391 2496 12403 2499
rect 12710 2496 12716 2508
rect 12391 2468 12716 2496
rect 12391 2465 12403 2468
rect 12345 2459 12403 2465
rect 12710 2456 12716 2468
rect 12768 2456 12774 2508
rect 12986 2456 12992 2508
rect 13044 2496 13050 2508
rect 14001 2499 14059 2505
rect 14001 2496 14013 2499
rect 13044 2468 14013 2496
rect 13044 2456 13050 2468
rect 14001 2465 14013 2468
rect 14047 2465 14059 2499
rect 14001 2459 14059 2465
rect 14090 2456 14096 2508
rect 14148 2456 14154 2508
rect 14734 2456 14740 2508
rect 14792 2456 14798 2508
rect 15010 2456 15016 2508
rect 15068 2456 15074 2508
rect 15289 2499 15347 2505
rect 15289 2465 15301 2499
rect 15335 2465 15347 2499
rect 15289 2459 15347 2465
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 12032 2400 13277 2428
rect 12032 2388 12038 2400
rect 13265 2397 13277 2400
rect 13311 2428 13323 2431
rect 13311 2400 14044 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 12621 2363 12679 2369
rect 12621 2360 12633 2363
rect 11256 2332 12633 2360
rect 10376 2320 10382 2332
rect 12621 2329 12633 2332
rect 12667 2360 12679 2363
rect 12986 2360 12992 2372
rect 12667 2332 12992 2360
rect 12667 2329 12679 2332
rect 12621 2323 12679 2329
rect 12986 2320 12992 2332
rect 13044 2320 13050 2372
rect 9585 2295 9643 2301
rect 9585 2261 9597 2295
rect 9631 2292 9643 2295
rect 9674 2292 9680 2304
rect 9631 2264 9680 2292
rect 9631 2261 9643 2264
rect 9585 2255 9643 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 10134 2252 10140 2304
rect 10192 2292 10198 2304
rect 10413 2295 10471 2301
rect 10413 2292 10425 2295
rect 10192 2264 10425 2292
rect 10192 2252 10198 2264
rect 10413 2261 10425 2264
rect 10459 2261 10471 2295
rect 10413 2255 10471 2261
rect 10781 2295 10839 2301
rect 10781 2261 10793 2295
rect 10827 2292 10839 2295
rect 13262 2292 13268 2304
rect 10827 2264 13268 2292
rect 10827 2261 10839 2264
rect 10781 2255 10839 2261
rect 13262 2252 13268 2264
rect 13320 2252 13326 2304
rect 13354 2252 13360 2304
rect 13412 2252 13418 2304
rect 13538 2252 13544 2304
rect 13596 2252 13602 2304
rect 13630 2252 13636 2304
rect 13688 2292 13694 2304
rect 13817 2295 13875 2301
rect 13817 2292 13829 2295
rect 13688 2264 13829 2292
rect 13688 2252 13694 2264
rect 13817 2261 13829 2264
rect 13863 2261 13875 2295
rect 14016 2292 14044 2400
rect 14366 2388 14372 2440
rect 14424 2428 14430 2440
rect 14752 2428 14780 2456
rect 15304 2428 15332 2459
rect 15378 2456 15384 2508
rect 15436 2456 15442 2508
rect 15565 2499 15623 2505
rect 15565 2465 15577 2499
rect 15611 2465 15623 2499
rect 15565 2459 15623 2465
rect 17129 2499 17187 2505
rect 17129 2465 17141 2499
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 15580 2428 15608 2459
rect 14424 2400 15332 2428
rect 15488 2400 15608 2428
rect 14424 2388 14430 2400
rect 14642 2320 14648 2372
rect 14700 2360 14706 2372
rect 15010 2360 15016 2372
rect 14700 2332 15016 2360
rect 14700 2320 14706 2332
rect 15010 2320 15016 2332
rect 15068 2360 15074 2372
rect 15488 2360 15516 2400
rect 16666 2388 16672 2440
rect 16724 2388 16730 2440
rect 17144 2428 17172 2459
rect 17218 2456 17224 2508
rect 17276 2456 17282 2508
rect 17328 2505 17356 2536
rect 17512 2505 17540 2604
rect 17862 2592 17868 2604
rect 17920 2632 17926 2644
rect 19426 2632 19432 2644
rect 17920 2604 19432 2632
rect 17920 2592 17926 2604
rect 19426 2592 19432 2604
rect 19484 2592 19490 2644
rect 19889 2635 19947 2641
rect 19889 2601 19901 2635
rect 19935 2601 19947 2635
rect 19889 2595 19947 2601
rect 21269 2635 21327 2641
rect 21269 2601 21281 2635
rect 21315 2632 21327 2635
rect 21726 2632 21732 2644
rect 21315 2604 21732 2632
rect 21315 2601 21327 2604
rect 21269 2595 21327 2601
rect 18776 2567 18834 2573
rect 18776 2533 18788 2567
rect 18822 2564 18834 2567
rect 19334 2564 19340 2576
rect 18822 2536 19340 2564
rect 18822 2533 18834 2536
rect 18776 2527 18834 2533
rect 19334 2524 19340 2536
rect 19392 2524 19398 2576
rect 19904 2564 19932 2595
rect 21726 2592 21732 2604
rect 21784 2592 21790 2644
rect 22370 2592 22376 2644
rect 22428 2632 22434 2644
rect 22646 2632 22652 2644
rect 22428 2604 22652 2632
rect 22428 2592 22434 2604
rect 22646 2592 22652 2604
rect 22704 2632 22710 2644
rect 23014 2632 23020 2644
rect 22704 2604 23020 2632
rect 22704 2592 22710 2604
rect 23014 2592 23020 2604
rect 23072 2592 23078 2644
rect 23385 2635 23443 2641
rect 23385 2601 23397 2635
rect 23431 2632 23443 2635
rect 24026 2632 24032 2644
rect 23431 2604 24032 2632
rect 23431 2601 23443 2604
rect 23385 2595 23443 2601
rect 24026 2592 24032 2604
rect 24084 2592 24090 2644
rect 23109 2567 23167 2573
rect 23109 2564 23121 2567
rect 19904 2536 23121 2564
rect 17313 2499 17371 2505
rect 17313 2465 17325 2499
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 17497 2499 17555 2505
rect 17497 2465 17509 2499
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 18046 2456 18052 2508
rect 18104 2496 18110 2508
rect 20640 2505 20668 2536
rect 23109 2533 23121 2536
rect 23155 2533 23167 2567
rect 25682 2564 25688 2576
rect 23109 2527 23167 2533
rect 23676 2536 25688 2564
rect 21450 2505 21456 2508
rect 20625 2499 20683 2505
rect 18104 2468 19564 2496
rect 18104 2456 18110 2468
rect 17589 2431 17647 2437
rect 17589 2428 17601 2431
rect 17144 2400 17601 2428
rect 17589 2397 17601 2400
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2397 18291 2431
rect 18233 2391 18291 2397
rect 15068 2332 15516 2360
rect 15749 2363 15807 2369
rect 15068 2320 15074 2332
rect 15749 2329 15761 2363
rect 15795 2360 15807 2363
rect 18046 2360 18052 2372
rect 15795 2332 18052 2360
rect 15795 2329 15807 2332
rect 15749 2323 15807 2329
rect 18046 2320 18052 2332
rect 18104 2320 18110 2372
rect 14458 2292 14464 2304
rect 14016 2264 14464 2292
rect 13817 2255 13875 2261
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 15102 2252 15108 2304
rect 15160 2292 15166 2304
rect 15197 2295 15255 2301
rect 15197 2292 15209 2295
rect 15160 2264 15209 2292
rect 15160 2252 15166 2264
rect 15197 2261 15209 2264
rect 15243 2261 15255 2295
rect 15197 2255 15255 2261
rect 15930 2252 15936 2304
rect 15988 2292 15994 2304
rect 16117 2295 16175 2301
rect 16117 2292 16129 2295
rect 15988 2264 16129 2292
rect 15988 2252 15994 2264
rect 16117 2261 16129 2264
rect 16163 2261 16175 2295
rect 16117 2255 16175 2261
rect 16850 2252 16856 2304
rect 16908 2252 16914 2304
rect 17586 2252 17592 2304
rect 17644 2292 17650 2304
rect 18248 2292 18276 2391
rect 18506 2388 18512 2440
rect 18564 2388 18570 2440
rect 19536 2428 19564 2468
rect 20625 2465 20637 2499
rect 20671 2465 20683 2499
rect 21448 2496 21456 2505
rect 21411 2468 21456 2496
rect 20625 2459 20683 2465
rect 21448 2459 21456 2468
rect 21450 2456 21456 2459
rect 21508 2456 21514 2508
rect 21545 2499 21603 2505
rect 21545 2465 21557 2499
rect 21591 2465 21603 2499
rect 21545 2459 21603 2465
rect 21637 2499 21695 2505
rect 21637 2465 21649 2499
rect 21683 2465 21695 2499
rect 21637 2459 21695 2465
rect 21560 2428 21588 2459
rect 19536 2400 21588 2428
rect 21652 2428 21680 2459
rect 21818 2456 21824 2508
rect 21876 2456 21882 2508
rect 21913 2499 21971 2505
rect 21913 2465 21925 2499
rect 21959 2496 21971 2499
rect 22002 2496 22008 2508
rect 21959 2468 22008 2496
rect 21959 2465 21971 2468
rect 21913 2459 21971 2465
rect 22002 2456 22008 2468
rect 22060 2456 22066 2508
rect 22186 2505 22192 2508
rect 22184 2496 22192 2505
rect 22147 2468 22192 2496
rect 22184 2459 22192 2468
rect 22186 2456 22192 2459
rect 22244 2456 22250 2508
rect 22278 2456 22284 2508
rect 22336 2456 22342 2508
rect 22370 2456 22376 2508
rect 22428 2456 22434 2508
rect 22462 2456 22468 2508
rect 22520 2505 22526 2508
rect 22520 2499 22559 2505
rect 22547 2465 22559 2499
rect 22520 2459 22559 2465
rect 22649 2499 22707 2505
rect 22649 2465 22661 2499
rect 22695 2496 22707 2499
rect 22741 2499 22799 2505
rect 22741 2496 22753 2499
rect 22695 2468 22753 2496
rect 22695 2465 22707 2468
rect 22649 2459 22707 2465
rect 22741 2465 22753 2468
rect 22787 2465 22799 2499
rect 22741 2459 22799 2465
rect 22889 2499 22947 2505
rect 22889 2465 22901 2499
rect 22935 2496 22947 2499
rect 22935 2465 22968 2496
rect 22889 2459 22968 2465
rect 22520 2456 22526 2459
rect 22388 2428 22416 2456
rect 21652 2400 22416 2428
rect 22646 2360 22652 2372
rect 19444 2332 22652 2360
rect 19444 2292 19472 2332
rect 22646 2320 22652 2332
rect 22704 2320 22710 2372
rect 22756 2360 22784 2459
rect 22940 2428 22968 2459
rect 23014 2456 23020 2508
rect 23072 2456 23078 2508
rect 23198 2456 23204 2508
rect 23256 2505 23262 2508
rect 23256 2496 23264 2505
rect 23256 2468 23301 2496
rect 23256 2459 23264 2468
rect 23256 2456 23262 2459
rect 23676 2428 23704 2536
rect 25682 2524 25688 2536
rect 25740 2564 25746 2576
rect 26053 2567 26111 2573
rect 26053 2564 26065 2567
rect 25740 2536 26065 2564
rect 25740 2524 25746 2536
rect 26053 2533 26065 2536
rect 26099 2533 26111 2567
rect 26053 2527 26111 2533
rect 24204 2499 24262 2505
rect 24204 2465 24216 2499
rect 24250 2496 24262 2499
rect 26421 2499 26479 2505
rect 26421 2496 26433 2499
rect 24250 2468 26433 2496
rect 24250 2465 24262 2468
rect 24204 2459 24262 2465
rect 26421 2465 26433 2468
rect 26467 2465 26479 2499
rect 26421 2459 26479 2465
rect 22940 2400 23704 2428
rect 23750 2388 23756 2440
rect 23808 2428 23814 2440
rect 23937 2431 23995 2437
rect 23937 2428 23949 2431
rect 23808 2400 23949 2428
rect 23808 2388 23814 2400
rect 23937 2397 23949 2400
rect 23983 2397 23995 2431
rect 23937 2391 23995 2397
rect 25409 2431 25467 2437
rect 25409 2397 25421 2431
rect 25455 2397 25467 2431
rect 25409 2391 25467 2397
rect 23382 2360 23388 2372
rect 22756 2332 23388 2360
rect 17644 2264 19472 2292
rect 17644 2252 17650 2264
rect 19978 2252 19984 2304
rect 20036 2252 20042 2304
rect 21726 2252 21732 2304
rect 21784 2292 21790 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21784 2264 22017 2292
rect 21784 2252 21790 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 22094 2252 22100 2304
rect 22152 2292 22158 2304
rect 22756 2292 22784 2332
rect 23382 2320 23388 2332
rect 23440 2320 23446 2372
rect 25317 2363 25375 2369
rect 25317 2329 25329 2363
rect 25363 2360 25375 2363
rect 25424 2360 25452 2391
rect 25958 2388 25964 2440
rect 26016 2428 26022 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26016 2400 26985 2428
rect 26016 2388 26022 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 25363 2332 25452 2360
rect 25363 2329 25375 2332
rect 25317 2323 25375 2329
rect 22152 2264 22784 2292
rect 22152 2252 22158 2264
rect 23014 2252 23020 2304
rect 23072 2292 23078 2304
rect 24302 2292 24308 2304
rect 23072 2264 24308 2292
rect 23072 2252 23078 2264
rect 24302 2252 24308 2264
rect 24360 2252 24366 2304
rect 25222 2252 25228 2304
rect 25280 2292 25286 2304
rect 25866 2292 25872 2304
rect 25280 2264 25872 2292
rect 25280 2252 25286 2264
rect 25866 2252 25872 2264
rect 25924 2252 25930 2304
rect 552 2202 27416 2224
rect 552 2150 3756 2202
rect 3808 2150 3820 2202
rect 3872 2150 3884 2202
rect 3936 2150 3948 2202
rect 4000 2150 4012 2202
rect 4064 2150 10472 2202
rect 10524 2150 10536 2202
rect 10588 2150 10600 2202
rect 10652 2150 10664 2202
rect 10716 2150 10728 2202
rect 10780 2150 17188 2202
rect 17240 2150 17252 2202
rect 17304 2150 17316 2202
rect 17368 2150 17380 2202
rect 17432 2150 17444 2202
rect 17496 2150 23904 2202
rect 23956 2150 23968 2202
rect 24020 2150 24032 2202
rect 24084 2150 24096 2202
rect 24148 2150 24160 2202
rect 24212 2150 27416 2202
rect 552 2128 27416 2150
rect 9674 2048 9680 2100
rect 9732 2048 9738 2100
rect 10229 2091 10287 2097
rect 10229 2057 10241 2091
rect 10275 2088 10287 2091
rect 10962 2088 10968 2100
rect 10275 2060 10968 2088
rect 10275 2057 10287 2060
rect 10229 2051 10287 2057
rect 9401 1887 9459 1893
rect 9401 1853 9413 1887
rect 9447 1884 9459 1887
rect 10134 1884 10140 1896
rect 9447 1856 9536 1884
rect 9646 1859 10140 1884
rect 9447 1853 9459 1856
rect 9401 1847 9459 1853
rect 9214 1708 9220 1760
rect 9272 1708 9278 1760
rect 9508 1757 9536 1856
rect 9631 1856 10140 1859
rect 9631 1853 9689 1856
rect 9631 1819 9643 1853
rect 9677 1819 9689 1853
rect 10134 1844 10140 1856
rect 10192 1844 10198 1896
rect 10138 1831 10150 1844
rect 10184 1831 10196 1844
rect 9631 1813 9689 1819
rect 9858 1776 9864 1828
rect 9916 1776 9922 1828
rect 10138 1825 10196 1831
rect 9493 1751 9551 1757
rect 9493 1717 9505 1751
rect 9539 1717 9551 1751
rect 10152 1748 10180 1825
rect 10244 1816 10272 2051
rect 10962 2048 10968 2060
rect 11020 2048 11026 2100
rect 11054 2048 11060 2100
rect 11112 2088 11118 2100
rect 11241 2091 11299 2097
rect 11241 2088 11253 2091
rect 11112 2060 11253 2088
rect 11112 2048 11118 2060
rect 11241 2057 11253 2060
rect 11287 2057 11299 2091
rect 13538 2088 13544 2100
rect 11241 2051 11299 2057
rect 11992 2060 13544 2088
rect 10321 2023 10379 2029
rect 10321 1989 10333 2023
rect 10367 2020 10379 2023
rect 11992 2020 12020 2060
rect 13538 2048 13544 2060
rect 13596 2048 13602 2100
rect 14274 2048 14280 2100
rect 14332 2048 14338 2100
rect 15565 2091 15623 2097
rect 15565 2057 15577 2091
rect 15611 2088 15623 2091
rect 16666 2088 16672 2100
rect 15611 2060 16672 2088
rect 15611 2057 15623 2060
rect 15565 2051 15623 2057
rect 16666 2048 16672 2060
rect 16724 2048 16730 2100
rect 18509 2091 18567 2097
rect 18509 2057 18521 2091
rect 18555 2088 18567 2091
rect 18690 2088 18696 2100
rect 18555 2060 18696 2088
rect 18555 2057 18567 2060
rect 18509 2051 18567 2057
rect 18690 2048 18696 2060
rect 18748 2048 18754 2100
rect 22278 2088 22284 2100
rect 18800 2060 22284 2088
rect 10367 1992 12020 2020
rect 17037 2023 17095 2029
rect 10367 1989 10379 1992
rect 10321 1983 10379 1989
rect 17037 1989 17049 2023
rect 17083 2020 17095 2023
rect 17083 1992 17816 2020
rect 17083 1989 17095 1992
rect 17037 1983 17095 1989
rect 10413 1955 10471 1961
rect 10413 1921 10425 1955
rect 10459 1952 10471 1955
rect 10594 1952 10600 1964
rect 10459 1924 10600 1952
rect 10459 1921 10471 1924
rect 10413 1915 10471 1921
rect 10594 1912 10600 1924
rect 10652 1912 10658 1964
rect 11514 1952 11520 1964
rect 10704 1924 11520 1952
rect 10502 1844 10508 1896
rect 10560 1844 10566 1896
rect 10704 1893 10732 1924
rect 11514 1912 11520 1924
rect 11572 1912 11578 1964
rect 13357 1955 13415 1961
rect 13357 1921 13369 1955
rect 13403 1952 13415 1955
rect 15654 1952 15660 1964
rect 13403 1924 15660 1952
rect 13403 1921 13415 1924
rect 13357 1915 13415 1921
rect 15654 1912 15660 1924
rect 15712 1912 15718 1964
rect 17788 1961 17816 1992
rect 18138 1980 18144 2032
rect 18196 2020 18202 2032
rect 18414 2020 18420 2032
rect 18196 1992 18420 2020
rect 18196 1980 18202 1992
rect 18414 1980 18420 1992
rect 18472 1980 18478 2032
rect 17773 1955 17831 1961
rect 17773 1921 17785 1955
rect 17819 1952 17831 1955
rect 18800 1952 18828 2060
rect 22278 2048 22284 2060
rect 22336 2048 22342 2100
rect 22370 2048 22376 2100
rect 22428 2088 22434 2100
rect 22428 2060 24992 2088
rect 22428 2048 22434 2060
rect 19978 2020 19984 2032
rect 17819 1924 18828 1952
rect 18892 1992 19984 2020
rect 17819 1921 17831 1924
rect 17773 1915 17831 1921
rect 10689 1887 10747 1893
rect 10689 1853 10701 1887
rect 10735 1853 10747 1887
rect 10689 1847 10747 1853
rect 10781 1887 10839 1893
rect 10781 1853 10793 1887
rect 10827 1853 10839 1887
rect 10781 1847 10839 1853
rect 10873 1887 10931 1893
rect 10873 1853 10885 1887
rect 10919 1853 10931 1887
rect 10873 1847 10931 1853
rect 11885 1887 11943 1893
rect 11885 1853 11897 1887
rect 11931 1884 11943 1887
rect 12342 1884 12348 1896
rect 11931 1856 12348 1884
rect 11931 1853 11943 1856
rect 11885 1847 11943 1853
rect 10796 1816 10824 1847
rect 10244 1788 10824 1816
rect 10888 1748 10916 1847
rect 12342 1844 12348 1856
rect 12400 1844 12406 1896
rect 13101 1887 13159 1893
rect 13101 1853 13113 1887
rect 13147 1884 13159 1887
rect 13630 1884 13636 1896
rect 13147 1856 13636 1884
rect 13147 1853 13159 1856
rect 13101 1847 13159 1853
rect 13630 1844 13636 1856
rect 13688 1844 13694 1896
rect 13817 1887 13875 1893
rect 13817 1853 13829 1887
rect 13863 1884 13875 1887
rect 14093 1887 14151 1893
rect 13863 1856 14044 1884
rect 13863 1853 13875 1856
rect 13817 1847 13875 1853
rect 10152 1720 10916 1748
rect 9493 1711 9551 1717
rect 11146 1708 11152 1760
rect 11204 1708 11210 1760
rect 11974 1708 11980 1760
rect 12032 1708 12038 1760
rect 13170 1708 13176 1760
rect 13228 1748 13234 1760
rect 13909 1751 13967 1757
rect 13909 1748 13921 1751
rect 13228 1720 13921 1748
rect 13228 1708 13234 1720
rect 13909 1717 13921 1720
rect 13955 1717 13967 1751
rect 14016 1748 14044 1856
rect 14093 1853 14105 1887
rect 14139 1853 14151 1887
rect 14093 1847 14151 1853
rect 14108 1816 14136 1847
rect 14366 1844 14372 1896
rect 14424 1844 14430 1896
rect 14458 1844 14464 1896
rect 14516 1844 14522 1896
rect 14642 1844 14648 1896
rect 14700 1844 14706 1896
rect 14921 1887 14979 1893
rect 14921 1853 14933 1887
rect 14967 1853 14979 1887
rect 14921 1847 14979 1853
rect 14660 1816 14688 1844
rect 14108 1788 14688 1816
rect 14366 1748 14372 1760
rect 14016 1720 14372 1748
rect 13909 1711 13967 1717
rect 14366 1708 14372 1720
rect 14424 1708 14430 1760
rect 14826 1708 14832 1760
rect 14884 1708 14890 1760
rect 14936 1748 14964 1847
rect 15102 1844 15108 1896
rect 15160 1844 15166 1896
rect 15194 1844 15200 1896
rect 15252 1844 15258 1896
rect 15930 1893 15936 1896
rect 15289 1887 15347 1893
rect 15289 1853 15301 1887
rect 15335 1853 15347 1887
rect 15924 1884 15936 1893
rect 15891 1856 15936 1884
rect 15289 1847 15347 1853
rect 15924 1847 15936 1856
rect 15304 1816 15332 1847
rect 15930 1844 15936 1847
rect 15988 1844 15994 1896
rect 17862 1844 17868 1896
rect 17920 1844 17926 1896
rect 18046 1844 18052 1896
rect 18104 1844 18110 1896
rect 18138 1844 18144 1896
rect 18196 1844 18202 1896
rect 18233 1887 18291 1893
rect 18233 1853 18245 1887
rect 18279 1884 18291 1887
rect 18892 1884 18920 1992
rect 19978 1980 19984 1992
rect 20036 1980 20042 2032
rect 21453 2023 21511 2029
rect 21453 1989 21465 2023
rect 21499 2020 21511 2023
rect 24302 2020 24308 2032
rect 21499 1992 22564 2020
rect 21499 1989 21511 1992
rect 21453 1983 21511 1989
rect 19886 1912 19892 1964
rect 19944 1952 19950 1964
rect 20073 1955 20131 1961
rect 20073 1952 20085 1955
rect 19944 1924 20085 1952
rect 19944 1912 19950 1924
rect 20073 1921 20085 1924
rect 20119 1921 20131 1955
rect 20073 1915 20131 1921
rect 22186 1912 22192 1964
rect 22244 1952 22250 1964
rect 22370 1952 22376 1964
rect 22244 1924 22376 1952
rect 22244 1912 22250 1924
rect 22370 1912 22376 1924
rect 22428 1912 22434 1964
rect 22536 1952 22564 1992
rect 24228 1992 24308 2020
rect 23569 1955 23627 1961
rect 23569 1952 23581 1955
rect 22536 1924 23581 1952
rect 23569 1921 23581 1924
rect 23615 1921 23627 1955
rect 23569 1915 23627 1921
rect 18279 1856 18920 1884
rect 18279 1853 18291 1856
rect 18233 1847 18291 1853
rect 18966 1844 18972 1896
rect 19024 1844 19030 1896
rect 19058 1844 19064 1896
rect 19116 1844 19122 1896
rect 19153 1887 19211 1893
rect 19153 1853 19165 1887
rect 19199 1853 19211 1887
rect 19153 1847 19211 1853
rect 19337 1887 19395 1893
rect 19337 1853 19349 1887
rect 19383 1884 19395 1887
rect 19426 1884 19432 1896
rect 19383 1856 19432 1884
rect 19383 1853 19395 1856
rect 19337 1847 19395 1853
rect 17129 1819 17187 1825
rect 17129 1816 17141 1819
rect 15304 1788 17141 1816
rect 17129 1785 17141 1788
rect 17175 1785 17187 1819
rect 17129 1779 17187 1785
rect 17954 1776 17960 1828
rect 18012 1816 18018 1828
rect 19168 1816 19196 1847
rect 19426 1844 19432 1856
rect 19484 1844 19490 1896
rect 20898 1844 20904 1896
rect 20956 1884 20962 1896
rect 21545 1887 21603 1893
rect 21545 1884 21557 1887
rect 20956 1856 21557 1884
rect 20956 1844 20962 1856
rect 21545 1853 21557 1856
rect 21591 1853 21603 1887
rect 21545 1847 21603 1853
rect 22830 1844 22836 1896
rect 22888 1844 22894 1896
rect 23382 1844 23388 1896
rect 23440 1884 23446 1896
rect 23845 1887 23903 1893
rect 23845 1884 23857 1887
rect 23440 1856 23857 1884
rect 23440 1844 23446 1856
rect 23845 1853 23857 1856
rect 23891 1853 23903 1887
rect 23845 1847 23903 1853
rect 23938 1887 23996 1893
rect 23938 1853 23950 1887
rect 23984 1853 23996 1887
rect 24228 1884 24256 1992
rect 24302 1980 24308 1992
rect 24360 2020 24366 2032
rect 24360 1992 24900 2020
rect 24360 1980 24366 1992
rect 23938 1847 23996 1853
rect 24136 1856 24256 1884
rect 24310 1887 24368 1893
rect 18012 1788 19196 1816
rect 20340 1819 20398 1825
rect 18012 1776 18018 1788
rect 20340 1785 20352 1819
rect 20386 1816 20398 1819
rect 22281 1819 22339 1825
rect 22281 1816 22293 1819
rect 20386 1788 22293 1816
rect 20386 1785 20398 1788
rect 20340 1779 20398 1785
rect 22281 1785 22293 1788
rect 22327 1785 22339 1819
rect 22281 1779 22339 1785
rect 23474 1776 23480 1828
rect 23532 1816 23538 1828
rect 23952 1816 23980 1847
rect 24136 1825 24164 1856
rect 24310 1853 24322 1887
rect 24356 1853 24368 1887
rect 24310 1847 24368 1853
rect 23532 1788 23980 1816
rect 24121 1819 24179 1825
rect 23532 1776 23538 1788
rect 24121 1785 24133 1819
rect 24167 1785 24179 1819
rect 24121 1779 24179 1785
rect 24210 1776 24216 1828
rect 24268 1776 24274 1828
rect 24320 1816 24348 1847
rect 24486 1844 24492 1896
rect 24544 1884 24550 1896
rect 24762 1893 24768 1896
rect 24581 1887 24639 1893
rect 24581 1884 24593 1887
rect 24544 1856 24593 1884
rect 24544 1844 24550 1856
rect 24581 1853 24593 1856
rect 24627 1853 24639 1887
rect 24581 1847 24639 1853
rect 24729 1887 24768 1893
rect 24729 1853 24741 1887
rect 24729 1847 24768 1853
rect 24762 1844 24768 1847
rect 24820 1844 24826 1896
rect 24872 1893 24900 1992
rect 24964 1893 24992 2060
rect 25958 2048 25964 2100
rect 26016 2048 26022 2100
rect 25225 2023 25283 2029
rect 25225 1989 25237 2023
rect 25271 1989 25283 2023
rect 25225 1983 25283 1989
rect 25240 1952 25268 1983
rect 25240 1924 26280 1952
rect 24857 1887 24915 1893
rect 24857 1853 24869 1887
rect 24903 1853 24915 1887
rect 24857 1847 24915 1853
rect 24949 1887 25007 1893
rect 24949 1853 24961 1887
rect 24995 1853 25007 1887
rect 24949 1847 25007 1853
rect 25046 1887 25104 1893
rect 25046 1853 25058 1887
rect 25092 1853 25104 1887
rect 25046 1847 25104 1853
rect 25056 1816 25084 1847
rect 25222 1844 25228 1896
rect 25280 1884 25286 1896
rect 25317 1887 25375 1893
rect 25317 1884 25329 1887
rect 25280 1856 25329 1884
rect 25280 1844 25286 1856
rect 25317 1853 25329 1856
rect 25363 1853 25375 1887
rect 25317 1847 25375 1853
rect 25501 1887 25559 1893
rect 25501 1853 25513 1887
rect 25547 1853 25559 1887
rect 25501 1847 25559 1853
rect 24320 1788 25084 1816
rect 15286 1748 15292 1760
rect 14936 1720 15292 1748
rect 15286 1708 15292 1720
rect 15344 1708 15350 1760
rect 18690 1708 18696 1760
rect 18748 1708 18754 1760
rect 22462 1708 22468 1760
rect 22520 1748 22526 1760
rect 23017 1751 23075 1757
rect 23017 1748 23029 1751
rect 22520 1720 23029 1748
rect 22520 1708 22526 1720
rect 23017 1717 23029 1720
rect 23063 1717 23075 1751
rect 23017 1711 23075 1717
rect 23106 1708 23112 1760
rect 23164 1748 23170 1760
rect 24320 1748 24348 1788
rect 23164 1720 24348 1748
rect 24489 1751 24547 1757
rect 23164 1708 23170 1720
rect 24489 1717 24501 1751
rect 24535 1748 24547 1751
rect 25516 1748 25544 1847
rect 25590 1844 25596 1896
rect 25648 1844 25654 1896
rect 25682 1844 25688 1896
rect 25740 1844 25746 1896
rect 25866 1844 25872 1896
rect 25924 1884 25930 1896
rect 26252 1893 26280 1924
rect 26053 1887 26111 1893
rect 26053 1884 26065 1887
rect 25924 1856 26065 1884
rect 25924 1844 25930 1856
rect 26053 1853 26065 1856
rect 26099 1853 26111 1887
rect 26053 1847 26111 1853
rect 26237 1887 26295 1893
rect 26237 1853 26249 1887
rect 26283 1853 26295 1887
rect 26237 1847 26295 1853
rect 26329 1887 26387 1893
rect 26329 1853 26341 1887
rect 26375 1853 26387 1887
rect 26329 1847 26387 1853
rect 26421 1887 26479 1893
rect 26421 1853 26433 1887
rect 26467 1853 26479 1887
rect 26421 1847 26479 1853
rect 25608 1816 25636 1844
rect 26344 1816 26372 1847
rect 25608 1788 26372 1816
rect 24535 1720 25544 1748
rect 24535 1717 24547 1720
rect 24489 1711 24547 1717
rect 25774 1708 25780 1760
rect 25832 1748 25838 1760
rect 26436 1748 26464 1847
rect 25832 1720 26464 1748
rect 25832 1708 25838 1720
rect 26694 1708 26700 1760
rect 26752 1708 26758 1760
rect 552 1658 27576 1680
rect 552 1606 7114 1658
rect 7166 1606 7178 1658
rect 7230 1606 7242 1658
rect 7294 1606 7306 1658
rect 7358 1606 7370 1658
rect 7422 1606 13830 1658
rect 13882 1606 13894 1658
rect 13946 1606 13958 1658
rect 14010 1606 14022 1658
rect 14074 1606 14086 1658
rect 14138 1606 20546 1658
rect 20598 1606 20610 1658
rect 20662 1606 20674 1658
rect 20726 1606 20738 1658
rect 20790 1606 20802 1658
rect 20854 1606 27262 1658
rect 27314 1606 27326 1658
rect 27378 1606 27390 1658
rect 27442 1606 27454 1658
rect 27506 1606 27518 1658
rect 27570 1606 27576 1658
rect 552 1584 27576 1606
rect 8386 1504 8392 1556
rect 8444 1544 8450 1556
rect 9858 1544 9864 1556
rect 8444 1516 9864 1544
rect 8444 1504 8450 1516
rect 9858 1504 9864 1516
rect 9916 1504 9922 1556
rect 10042 1504 10048 1556
rect 10100 1544 10106 1556
rect 10137 1547 10195 1553
rect 10137 1544 10149 1547
rect 10100 1516 10149 1544
rect 10100 1504 10106 1516
rect 10137 1513 10149 1516
rect 10183 1513 10195 1547
rect 10137 1507 10195 1513
rect 10594 1504 10600 1556
rect 10652 1544 10658 1556
rect 14093 1547 14151 1553
rect 10652 1516 11376 1544
rect 10652 1504 10658 1516
rect 9024 1479 9082 1485
rect 9024 1445 9036 1479
rect 9070 1476 9082 1479
rect 9214 1476 9220 1488
rect 9070 1448 9220 1476
rect 9070 1445 9082 1448
rect 9024 1439 9082 1445
rect 9214 1436 9220 1448
rect 9272 1436 9278 1488
rect 11146 1436 11152 1488
rect 11204 1476 11210 1488
rect 11204 1448 11284 1476
rect 11204 1436 11210 1448
rect 11256 1417 11284 1448
rect 11232 1411 11290 1417
rect 11232 1377 11244 1411
rect 11278 1377 11290 1411
rect 11348 1408 11376 1516
rect 14093 1513 14105 1547
rect 14139 1513 14151 1547
rect 14093 1507 14151 1513
rect 12710 1436 12716 1488
rect 12768 1476 12774 1488
rect 14108 1476 14136 1507
rect 14826 1504 14832 1556
rect 14884 1544 14890 1556
rect 19610 1544 19616 1556
rect 14884 1516 19616 1544
rect 14884 1504 14890 1516
rect 19610 1504 19616 1516
rect 19668 1504 19674 1556
rect 20533 1547 20591 1553
rect 20533 1513 20545 1547
rect 20579 1544 20591 1547
rect 22186 1544 22192 1556
rect 20579 1516 22192 1544
rect 20579 1513 20591 1516
rect 20533 1507 20591 1513
rect 22186 1504 22192 1516
rect 22244 1504 22250 1556
rect 23293 1547 23351 1553
rect 23293 1513 23305 1547
rect 23339 1513 23351 1547
rect 23293 1507 23351 1513
rect 15378 1476 15384 1488
rect 12768 1448 15384 1476
rect 12768 1436 12774 1448
rect 15378 1436 15384 1448
rect 15436 1436 15442 1488
rect 16384 1479 16442 1485
rect 16384 1445 16396 1479
rect 16430 1476 16442 1479
rect 16850 1476 16856 1488
rect 16430 1448 16856 1476
rect 16430 1445 16442 1448
rect 16384 1439 16442 1445
rect 16850 1436 16856 1448
rect 16908 1436 16914 1488
rect 18506 1436 18512 1488
rect 18564 1476 18570 1488
rect 18564 1448 19104 1476
rect 18564 1436 18570 1448
rect 12529 1411 12587 1417
rect 12529 1408 12541 1411
rect 11348 1380 12541 1408
rect 11232 1371 11290 1377
rect 12529 1377 12541 1380
rect 12575 1377 12587 1411
rect 12529 1371 12587 1377
rect 12629 1411 12687 1417
rect 12629 1377 12641 1411
rect 12675 1408 12687 1411
rect 12728 1408 12756 1436
rect 12675 1380 12756 1408
rect 12675 1377 12687 1380
rect 12629 1371 12687 1377
rect 12802 1368 12808 1420
rect 12860 1408 12866 1420
rect 12969 1411 13027 1417
rect 12969 1408 12981 1411
rect 12860 1380 12981 1408
rect 12860 1368 12866 1380
rect 12969 1377 12981 1380
rect 13015 1377 13027 1411
rect 12969 1371 13027 1377
rect 14366 1368 14372 1420
rect 14424 1408 14430 1420
rect 14645 1411 14703 1417
rect 14645 1408 14657 1411
rect 14424 1380 14657 1408
rect 14424 1368 14430 1380
rect 14645 1377 14657 1380
rect 14691 1377 14703 1411
rect 14645 1371 14703 1377
rect 14737 1411 14795 1417
rect 14737 1377 14749 1411
rect 14783 1377 14795 1411
rect 14737 1371 14795 1377
rect 14921 1411 14979 1417
rect 14921 1377 14933 1411
rect 14967 1408 14979 1411
rect 15010 1408 15016 1420
rect 14967 1380 15016 1408
rect 14967 1377 14979 1380
rect 14921 1371 14979 1377
rect 8757 1343 8815 1349
rect 8757 1309 8769 1343
rect 8803 1309 8815 1343
rect 8757 1303 8815 1309
rect 10965 1343 11023 1349
rect 10965 1309 10977 1343
rect 11011 1309 11023 1343
rect 12713 1343 12771 1349
rect 12713 1340 12725 1343
rect 10965 1303 11023 1309
rect 11992 1312 12725 1340
rect 8772 1204 8800 1303
rect 10980 1204 11008 1303
rect 11606 1204 11612 1216
rect 8772 1176 11612 1204
rect 11606 1164 11612 1176
rect 11664 1204 11670 1216
rect 11992 1204 12020 1312
rect 12713 1309 12725 1312
rect 12759 1309 12771 1343
rect 12713 1303 12771 1309
rect 11664 1176 12020 1204
rect 11664 1164 11670 1176
rect 12342 1164 12348 1216
rect 12400 1204 12406 1216
rect 14752 1204 14780 1371
rect 15010 1368 15016 1380
rect 15068 1368 15074 1420
rect 15654 1368 15660 1420
rect 15712 1408 15718 1420
rect 16022 1408 16028 1420
rect 15712 1380 16028 1408
rect 15712 1368 15718 1380
rect 16022 1368 16028 1380
rect 16080 1408 16086 1420
rect 19076 1417 19104 1448
rect 16117 1411 16175 1417
rect 16117 1408 16129 1411
rect 16080 1380 16129 1408
rect 16080 1368 16086 1380
rect 16117 1377 16129 1380
rect 16163 1377 16175 1411
rect 16117 1371 16175 1377
rect 18805 1411 18863 1417
rect 18805 1377 18817 1411
rect 18851 1408 18863 1411
rect 19061 1411 19119 1417
rect 18851 1380 19012 1408
rect 18851 1377 18863 1380
rect 18805 1371 18863 1377
rect 18984 1340 19012 1380
rect 19061 1377 19073 1411
rect 19107 1408 19119 1411
rect 19153 1411 19211 1417
rect 19153 1408 19165 1411
rect 19107 1380 19165 1408
rect 19107 1377 19119 1380
rect 19061 1371 19119 1377
rect 19153 1377 19165 1380
rect 19199 1377 19211 1411
rect 19153 1371 19211 1377
rect 19420 1411 19478 1417
rect 19420 1377 19432 1411
rect 19466 1408 19478 1411
rect 19794 1408 19800 1420
rect 19466 1380 19800 1408
rect 19466 1377 19478 1380
rect 19420 1371 19478 1377
rect 19794 1368 19800 1380
rect 19852 1368 19858 1420
rect 19886 1368 19892 1420
rect 19944 1408 19950 1420
rect 22180 1411 22238 1417
rect 19944 1380 20760 1408
rect 19944 1368 19950 1380
rect 20732 1340 20760 1380
rect 22180 1377 22192 1411
rect 22226 1408 22238 1411
rect 23198 1408 23204 1420
rect 22226 1380 23204 1408
rect 22226 1377 22238 1380
rect 22180 1371 22238 1377
rect 23198 1368 23204 1380
rect 23256 1368 23262 1420
rect 23308 1408 23336 1507
rect 24762 1504 24768 1556
rect 24820 1544 24826 1556
rect 24857 1547 24915 1553
rect 24857 1544 24869 1547
rect 24820 1516 24869 1544
rect 24820 1504 24826 1516
rect 24857 1513 24869 1516
rect 24903 1513 24915 1547
rect 24857 1507 24915 1513
rect 24520 1479 24578 1485
rect 24520 1445 24532 1479
rect 24566 1476 24578 1479
rect 25593 1479 25651 1485
rect 25593 1476 25605 1479
rect 24566 1448 25605 1476
rect 24566 1445 24578 1448
rect 24520 1439 24578 1445
rect 25593 1445 25605 1448
rect 25639 1445 25651 1479
rect 25593 1439 25651 1445
rect 26237 1411 26295 1417
rect 23308 1380 25452 1408
rect 25424 1349 25452 1380
rect 26237 1377 26249 1411
rect 26283 1408 26295 1411
rect 26694 1408 26700 1420
rect 26283 1380 26700 1408
rect 26283 1377 26295 1380
rect 26237 1371 26295 1377
rect 26694 1368 26700 1380
rect 26752 1368 26758 1420
rect 21913 1343 21971 1349
rect 21913 1340 21925 1343
rect 18984 1312 19196 1340
rect 20732 1312 21925 1340
rect 17954 1272 17960 1284
rect 17420 1244 17960 1272
rect 12400 1176 14780 1204
rect 15105 1207 15163 1213
rect 12400 1164 12406 1176
rect 15105 1173 15117 1207
rect 15151 1204 15163 1207
rect 17420 1204 17448 1244
rect 17954 1232 17960 1244
rect 18012 1232 18018 1284
rect 15151 1176 17448 1204
rect 17497 1207 17555 1213
rect 15151 1173 15163 1176
rect 15105 1167 15163 1173
rect 17497 1173 17509 1207
rect 17543 1204 17555 1207
rect 17586 1204 17592 1216
rect 17543 1176 17592 1204
rect 17543 1173 17555 1176
rect 17497 1167 17555 1173
rect 17586 1164 17592 1176
rect 17644 1164 17650 1216
rect 17678 1164 17684 1216
rect 17736 1164 17742 1216
rect 19168 1204 19196 1312
rect 21913 1309 21925 1312
rect 21959 1309 21971 1343
rect 21913 1303 21971 1309
rect 24765 1343 24823 1349
rect 24765 1309 24777 1343
rect 24811 1309 24823 1343
rect 24765 1303 24823 1309
rect 25409 1343 25467 1349
rect 25409 1309 25421 1343
rect 25455 1309 25467 1343
rect 25409 1303 25467 1309
rect 19334 1204 19340 1216
rect 19168 1176 19340 1204
rect 19334 1164 19340 1176
rect 19392 1164 19398 1216
rect 21928 1204 21956 1303
rect 23750 1272 23756 1284
rect 23216 1244 23756 1272
rect 23216 1204 23244 1244
rect 23750 1232 23756 1244
rect 23808 1272 23814 1284
rect 23808 1244 23888 1272
rect 23808 1232 23814 1244
rect 21928 1176 23244 1204
rect 23385 1207 23443 1213
rect 23385 1173 23397 1207
rect 23431 1204 23443 1207
rect 23474 1204 23480 1216
rect 23431 1176 23480 1204
rect 23431 1173 23443 1176
rect 23385 1167 23443 1173
rect 23474 1164 23480 1176
rect 23532 1164 23538 1216
rect 23860 1204 23888 1244
rect 24780 1204 24808 1303
rect 23860 1176 24808 1204
rect 552 1114 27416 1136
rect 552 1062 3756 1114
rect 3808 1062 3820 1114
rect 3872 1062 3884 1114
rect 3936 1062 3948 1114
rect 4000 1062 4012 1114
rect 4064 1062 10472 1114
rect 10524 1062 10536 1114
rect 10588 1062 10600 1114
rect 10652 1062 10664 1114
rect 10716 1062 10728 1114
rect 10780 1062 17188 1114
rect 17240 1062 17252 1114
rect 17304 1062 17316 1114
rect 17368 1062 17380 1114
rect 17432 1062 17444 1114
rect 17496 1062 23904 1114
rect 23956 1062 23968 1114
rect 24020 1062 24032 1114
rect 24084 1062 24096 1114
rect 24148 1062 24160 1114
rect 24212 1062 27416 1114
rect 552 1040 27416 1062
rect 12621 1003 12679 1009
rect 12621 969 12633 1003
rect 12667 1000 12679 1003
rect 12802 1000 12808 1012
rect 12667 972 12808 1000
rect 12667 969 12679 972
rect 12621 963 12679 969
rect 12802 960 12808 972
rect 12860 960 12866 1012
rect 18509 1003 18567 1009
rect 18509 969 18521 1003
rect 18555 1000 18567 1003
rect 18966 1000 18972 1012
rect 18555 972 18972 1000
rect 18555 969 18567 972
rect 18509 963 18567 969
rect 18966 960 18972 972
rect 19024 960 19030 1012
rect 19334 960 19340 1012
rect 19392 960 19398 1012
rect 19794 960 19800 1012
rect 19852 1000 19858 1012
rect 20073 1003 20131 1009
rect 20073 1000 20085 1003
rect 19852 972 20085 1000
rect 19852 960 19858 972
rect 20073 969 20085 972
rect 20119 969 20131 1003
rect 20073 963 20131 969
rect 22189 1003 22247 1009
rect 22189 969 22201 1003
rect 22235 1000 22247 1003
rect 22830 1000 22836 1012
rect 22235 972 22836 1000
rect 22235 969 22247 972
rect 22189 963 22247 969
rect 22830 960 22836 972
rect 22888 960 22894 1012
rect 23198 960 23204 1012
rect 23256 1000 23262 1012
rect 23845 1003 23903 1009
rect 23845 1000 23857 1003
rect 23256 972 23857 1000
rect 23256 960 23262 972
rect 23845 969 23857 972
rect 23891 969 23903 1003
rect 23845 963 23903 969
rect 25225 1003 25283 1009
rect 25225 969 25237 1003
rect 25271 1000 25283 1003
rect 25774 1000 25780 1012
rect 25271 972 25780 1000
rect 25271 969 25283 972
rect 25225 963 25283 969
rect 25774 960 25780 972
rect 25832 960 25838 1012
rect 22738 892 22744 944
rect 22796 932 22802 944
rect 23290 932 23296 944
rect 22796 904 23296 932
rect 22796 892 22802 904
rect 23290 892 23296 904
rect 23348 892 23354 944
rect 24762 932 24768 944
rect 23400 904 24768 932
rect 17678 824 17684 876
rect 17736 864 17742 876
rect 17865 867 17923 873
rect 17865 864 17877 867
rect 17736 836 17877 864
rect 17736 824 17742 836
rect 17865 833 17877 836
rect 17911 833 17923 867
rect 17865 827 17923 833
rect 18690 824 18696 876
rect 18748 824 18754 876
rect 19058 824 19064 876
rect 19116 864 19122 876
rect 19116 836 19748 864
rect 19116 824 19122 836
rect 12437 799 12495 805
rect 12437 765 12449 799
rect 12483 796 12495 799
rect 13354 796 13360 808
rect 12483 768 13360 796
rect 12483 765 12495 768
rect 12437 759 12495 765
rect 13354 756 13360 768
rect 13412 756 13418 808
rect 19426 756 19432 808
rect 19484 756 19490 808
rect 19610 756 19616 808
rect 19668 756 19674 808
rect 19720 805 19748 836
rect 21652 836 23060 864
rect 21652 808 21680 836
rect 19705 799 19763 805
rect 19705 765 19717 799
rect 19751 765 19763 799
rect 19705 759 19763 765
rect 19797 799 19855 805
rect 19797 765 19809 799
rect 19843 796 19855 799
rect 20898 796 20904 808
rect 19843 768 20904 796
rect 19843 765 19855 768
rect 19797 759 19855 765
rect 20898 756 20904 768
rect 20956 756 20962 808
rect 21545 799 21603 805
rect 21545 765 21557 799
rect 21591 796 21603 799
rect 21634 796 21640 808
rect 21591 768 21640 796
rect 21591 765 21603 768
rect 21545 759 21603 765
rect 21634 756 21640 768
rect 21692 756 21698 808
rect 21726 756 21732 808
rect 21784 756 21790 808
rect 21821 799 21879 805
rect 21821 765 21833 799
rect 21867 765 21879 799
rect 21821 759 21879 765
rect 21913 799 21971 805
rect 21913 765 21925 799
rect 21959 765 21971 799
rect 21913 759 21971 765
rect 21836 660 21864 759
rect 21928 728 21956 759
rect 22094 756 22100 808
rect 22152 796 22158 808
rect 22462 805 22468 808
rect 22281 799 22339 805
rect 22281 796 22293 799
rect 22152 768 22293 796
rect 22152 756 22158 768
rect 22281 765 22293 768
rect 22327 765 22339 799
rect 22281 759 22339 765
rect 22429 799 22468 805
rect 22429 765 22441 799
rect 22429 759 22468 765
rect 22444 756 22468 759
rect 22520 756 22526 808
rect 22554 756 22560 808
rect 22612 756 22618 808
rect 22646 756 22652 808
rect 22704 756 22710 808
rect 22787 799 22845 805
rect 22787 765 22799 799
rect 22833 796 22845 799
rect 22922 796 22928 808
rect 22833 768 22928 796
rect 22833 765 22845 768
rect 22787 759 22845 765
rect 22922 756 22928 768
rect 22980 756 22986 808
rect 23032 805 23060 836
rect 23017 799 23075 805
rect 23017 765 23029 799
rect 23063 765 23075 799
rect 23017 759 23075 765
rect 23201 799 23259 805
rect 23201 765 23213 799
rect 23247 765 23259 799
rect 23201 759 23259 765
rect 22444 728 22472 756
rect 23216 728 23244 759
rect 23290 756 23296 808
rect 23348 756 23354 808
rect 23400 805 23428 904
rect 24762 892 24768 904
rect 24820 892 24826 944
rect 23661 867 23719 873
rect 23661 833 23673 867
rect 23707 864 23719 867
rect 24397 867 24455 873
rect 24397 864 24409 867
rect 23707 836 24409 864
rect 23707 833 23719 836
rect 23661 827 23719 833
rect 24397 833 24409 836
rect 24443 833 24455 867
rect 24397 827 24455 833
rect 23385 799 23443 805
rect 23385 765 23397 799
rect 23431 765 23443 799
rect 23385 759 23443 765
rect 23474 756 23480 808
rect 23532 796 23538 808
rect 24581 799 24639 805
rect 24581 796 24593 799
rect 23532 768 24593 796
rect 23532 756 23538 768
rect 24581 765 24593 768
rect 24627 765 24639 799
rect 24581 759 24639 765
rect 21928 700 22472 728
rect 22940 700 23244 728
rect 22738 660 22744 672
rect 21836 632 22744 660
rect 22738 620 22744 632
rect 22796 620 22802 672
rect 22940 669 22968 700
rect 22925 663 22983 669
rect 22925 629 22937 663
rect 22971 629 22983 663
rect 22925 623 22983 629
rect 552 570 27576 592
rect 552 518 7114 570
rect 7166 518 7178 570
rect 7230 518 7242 570
rect 7294 518 7306 570
rect 7358 518 7370 570
rect 7422 518 13830 570
rect 13882 518 13894 570
rect 13946 518 13958 570
rect 14010 518 14022 570
rect 14074 518 14086 570
rect 14138 518 20546 570
rect 20598 518 20610 570
rect 20662 518 20674 570
rect 20726 518 20738 570
rect 20790 518 20802 570
rect 20854 518 27262 570
rect 27314 518 27326 570
rect 27378 518 27390 570
rect 27442 518 27454 570
rect 27506 518 27518 570
rect 27570 518 27576 570
rect 552 496 27576 518
<< via1 >>
rect 3608 17484 3660 17536
rect 3976 17484 4028 17536
rect 5632 17484 5684 17536
rect 15476 17688 15528 17740
rect 10692 17620 10744 17672
rect 18696 17620 18748 17672
rect 9956 17552 10008 17604
rect 16672 17552 16724 17604
rect 10324 17484 10376 17536
rect 23204 17484 23256 17536
rect 23940 17484 23992 17536
rect 24308 17484 24360 17536
rect 3756 17382 3808 17434
rect 3820 17382 3872 17434
rect 3884 17382 3936 17434
rect 3948 17382 4000 17434
rect 4012 17382 4064 17434
rect 10472 17382 10524 17434
rect 10536 17382 10588 17434
rect 10600 17382 10652 17434
rect 10664 17382 10716 17434
rect 10728 17382 10780 17434
rect 17188 17382 17240 17434
rect 17252 17382 17304 17434
rect 17316 17382 17368 17434
rect 17380 17382 17432 17434
rect 17444 17382 17496 17434
rect 23904 17382 23956 17434
rect 23968 17382 24020 17434
rect 24032 17382 24084 17434
rect 24096 17382 24148 17434
rect 24160 17382 24212 17434
rect 2136 17323 2188 17332
rect 2136 17289 2145 17323
rect 2145 17289 2179 17323
rect 2179 17289 2188 17323
rect 2136 17280 2188 17289
rect 2688 17280 2740 17332
rect 3608 17280 3660 17332
rect 7288 17323 7340 17332
rect 7288 17289 7297 17323
rect 7297 17289 7331 17323
rect 7331 17289 7340 17323
rect 7288 17280 7340 17289
rect 7840 17280 7892 17332
rect 9128 17280 9180 17332
rect 9772 17280 9824 17332
rect 12348 17280 12400 17332
rect 12992 17280 13044 17332
rect 6736 17212 6788 17264
rect 15936 17212 15988 17264
rect 3424 17187 3476 17196
rect 3424 17153 3433 17187
rect 3433 17153 3467 17187
rect 3467 17153 3476 17187
rect 3424 17144 3476 17153
rect 4620 17144 4672 17196
rect 5264 17144 5316 17196
rect 7472 17144 7524 17196
rect 6552 17076 6604 17128
rect 9956 17144 10008 17196
rect 14924 17144 14976 17196
rect 16120 17212 16172 17264
rect 19616 17212 19668 17264
rect 16856 17144 16908 17196
rect 10324 17119 10376 17128
rect 10324 17085 10333 17119
rect 10333 17085 10367 17119
rect 10367 17085 10376 17119
rect 10324 17076 10376 17085
rect 12072 17119 12124 17128
rect 12072 17085 12081 17119
rect 12081 17085 12115 17119
rect 12115 17085 12124 17119
rect 12072 17076 12124 17085
rect 12348 17076 12400 17128
rect 12716 17119 12768 17128
rect 12716 17085 12725 17119
rect 12725 17085 12759 17119
rect 12759 17085 12768 17119
rect 12716 17076 12768 17085
rect 4160 16940 4212 16992
rect 6736 16940 6788 16992
rect 8944 16983 8996 16992
rect 8944 16949 8953 16983
rect 8953 16949 8987 16983
rect 8987 16949 8996 16983
rect 8944 16940 8996 16949
rect 9404 17008 9456 17060
rect 15476 17051 15528 17060
rect 15476 17017 15485 17051
rect 15485 17017 15519 17051
rect 15519 17017 15528 17051
rect 15476 17008 15528 17017
rect 16672 17076 16724 17128
rect 17592 17076 17644 17128
rect 18236 17119 18288 17128
rect 18236 17085 18245 17119
rect 18245 17085 18279 17119
rect 18279 17085 18288 17119
rect 18236 17076 18288 17085
rect 19432 17076 19484 17128
rect 21640 17119 21692 17128
rect 21640 17085 21649 17119
rect 21649 17085 21683 17119
rect 21683 17085 21692 17119
rect 21640 17076 21692 17085
rect 22008 17076 22060 17128
rect 23296 17144 23348 17196
rect 23112 17119 23164 17128
rect 23112 17085 23121 17119
rect 23121 17085 23155 17119
rect 23155 17085 23164 17119
rect 23112 17076 23164 17085
rect 22652 17008 22704 17060
rect 24308 17119 24360 17128
rect 24308 17085 24317 17119
rect 24317 17085 24351 17119
rect 24351 17085 24360 17119
rect 24308 17076 24360 17085
rect 24584 17076 24636 17128
rect 25228 17076 25280 17128
rect 25872 17076 25924 17128
rect 26792 17119 26844 17128
rect 26792 17085 26801 17119
rect 26801 17085 26835 17119
rect 26835 17085 26844 17119
rect 26792 17076 26844 17085
rect 23664 17008 23716 17060
rect 9864 16940 9916 16992
rect 11888 16983 11940 16992
rect 11888 16949 11897 16983
rect 11897 16949 11931 16983
rect 11931 16949 11940 16983
rect 11888 16940 11940 16949
rect 15108 16983 15160 16992
rect 15108 16949 15117 16983
rect 15117 16949 15151 16983
rect 15151 16949 15160 16983
rect 15108 16940 15160 16949
rect 15752 16940 15804 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 16764 16940 16816 16992
rect 17500 16940 17552 16992
rect 17684 16983 17736 16992
rect 17684 16949 17693 16983
rect 17693 16949 17727 16983
rect 17727 16949 17736 16983
rect 17684 16940 17736 16949
rect 20168 16940 20220 16992
rect 21456 16983 21508 16992
rect 21456 16949 21465 16983
rect 21465 16949 21499 16983
rect 21499 16949 21508 16983
rect 21456 16940 21508 16949
rect 22100 16983 22152 16992
rect 22100 16949 22109 16983
rect 22109 16949 22143 16983
rect 22143 16949 22152 16983
rect 22100 16940 22152 16949
rect 22744 16940 22796 16992
rect 22928 16940 22980 16992
rect 23572 16940 23624 16992
rect 26608 17051 26660 17060
rect 26608 17017 26617 17051
rect 26617 17017 26651 17051
rect 26651 17017 26660 17051
rect 26608 17008 26660 17017
rect 25320 16983 25372 16992
rect 25320 16949 25329 16983
rect 25329 16949 25363 16983
rect 25363 16949 25372 16983
rect 25320 16940 25372 16949
rect 25964 16983 26016 16992
rect 25964 16949 25973 16983
rect 25973 16949 26007 16983
rect 26007 16949 26016 16983
rect 25964 16940 26016 16949
rect 7114 16838 7166 16890
rect 7178 16838 7230 16890
rect 7242 16838 7294 16890
rect 7306 16838 7358 16890
rect 7370 16838 7422 16890
rect 13830 16838 13882 16890
rect 13894 16838 13946 16890
rect 13958 16838 14010 16890
rect 14022 16838 14074 16890
rect 14086 16838 14138 16890
rect 20546 16838 20598 16890
rect 20610 16838 20662 16890
rect 20674 16838 20726 16890
rect 20738 16838 20790 16890
rect 20802 16838 20854 16890
rect 27262 16838 27314 16890
rect 27326 16838 27378 16890
rect 27390 16838 27442 16890
rect 27454 16838 27506 16890
rect 27518 16838 27570 16890
rect 756 16736 808 16788
rect 5632 16779 5684 16788
rect 5632 16745 5641 16779
rect 5641 16745 5675 16779
rect 5675 16745 5684 16779
rect 5632 16736 5684 16745
rect 5908 16736 5960 16788
rect 9404 16779 9456 16788
rect 9404 16745 9413 16779
rect 9413 16745 9447 16779
rect 9447 16745 9456 16779
rect 9404 16736 9456 16745
rect 9864 16779 9916 16788
rect 9864 16745 9873 16779
rect 9873 16745 9907 16779
rect 9907 16745 9916 16779
rect 9864 16736 9916 16745
rect 11060 16736 11112 16788
rect 11704 16736 11756 16788
rect 13636 16736 13688 16788
rect 14096 16736 14148 16788
rect 4160 16668 4212 16720
rect 3240 16532 3292 16584
rect 6000 16643 6052 16652
rect 6000 16609 6009 16643
rect 6009 16609 6043 16643
rect 6043 16609 6052 16643
rect 6000 16600 6052 16609
rect 6736 16643 6788 16652
rect 6736 16609 6745 16643
rect 6745 16609 6779 16643
rect 6779 16609 6788 16643
rect 6736 16600 6788 16609
rect 6828 16600 6880 16652
rect 7472 16600 7524 16652
rect 8668 16600 8720 16652
rect 10232 16668 10284 16720
rect 8024 16575 8076 16584
rect 8024 16541 8033 16575
rect 8033 16541 8067 16575
rect 8067 16541 8076 16575
rect 8024 16532 8076 16541
rect 11336 16643 11388 16652
rect 11336 16609 11345 16643
rect 11345 16609 11379 16643
rect 11379 16609 11388 16643
rect 11336 16600 11388 16609
rect 11704 16643 11756 16652
rect 11704 16609 11713 16643
rect 11713 16609 11747 16643
rect 11747 16609 11756 16643
rect 11704 16600 11756 16609
rect 11888 16668 11940 16720
rect 13912 16600 13964 16652
rect 14188 16600 14240 16652
rect 14648 16668 14700 16720
rect 15108 16736 15160 16788
rect 15568 16736 15620 16788
rect 16948 16779 17000 16788
rect 16948 16745 16957 16779
rect 16957 16745 16991 16779
rect 16991 16745 17000 16779
rect 16948 16736 17000 16745
rect 17316 16736 17368 16788
rect 17500 16779 17552 16788
rect 17500 16745 17509 16779
rect 17509 16745 17543 16779
rect 17543 16745 17552 16779
rect 17500 16736 17552 16745
rect 15108 16643 15160 16652
rect 15108 16609 15117 16643
rect 15117 16609 15151 16643
rect 15151 16609 15160 16643
rect 15108 16600 15160 16609
rect 15660 16600 15712 16652
rect 16764 16711 16816 16720
rect 16764 16677 16773 16711
rect 16773 16677 16807 16711
rect 16807 16677 16816 16711
rect 16764 16668 16816 16677
rect 16120 16643 16172 16652
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 16580 16600 16632 16652
rect 17684 16668 17736 16720
rect 15292 16575 15344 16584
rect 15292 16541 15301 16575
rect 15301 16541 15335 16575
rect 15335 16541 15344 16575
rect 15292 16532 15344 16541
rect 17316 16532 17368 16584
rect 23480 16736 23532 16788
rect 19616 16668 19668 16720
rect 18512 16600 18564 16652
rect 20812 16643 20864 16652
rect 20812 16609 20830 16643
rect 20830 16609 20864 16643
rect 20812 16600 20864 16609
rect 19524 16575 19576 16584
rect 19524 16541 19533 16575
rect 19533 16541 19567 16575
rect 19567 16541 19576 16575
rect 19524 16532 19576 16541
rect 21088 16575 21140 16584
rect 21088 16541 21097 16575
rect 21097 16541 21131 16575
rect 21131 16541 21140 16575
rect 21088 16532 21140 16541
rect 22284 16668 22336 16720
rect 21456 16643 21508 16652
rect 21456 16609 21465 16643
rect 21465 16609 21499 16643
rect 21499 16609 21508 16643
rect 21456 16600 21508 16609
rect 21640 16643 21692 16652
rect 21640 16609 21649 16643
rect 21649 16609 21683 16643
rect 21683 16609 21692 16643
rect 21640 16600 21692 16609
rect 21916 16643 21968 16652
rect 21916 16609 21925 16643
rect 21925 16609 21959 16643
rect 21959 16609 21968 16643
rect 21916 16600 21968 16609
rect 22100 16643 22152 16652
rect 22100 16609 22109 16643
rect 22109 16609 22143 16643
rect 22143 16609 22152 16643
rect 22100 16600 22152 16609
rect 22468 16643 22520 16652
rect 22468 16609 22477 16643
rect 22477 16609 22511 16643
rect 22511 16609 22520 16643
rect 22468 16600 22520 16609
rect 22928 16600 22980 16652
rect 23572 16600 23624 16652
rect 25320 16668 25372 16720
rect 23756 16600 23808 16652
rect 24676 16600 24728 16652
rect 25044 16600 25096 16652
rect 23020 16532 23072 16584
rect 17132 16464 17184 16516
rect 17776 16464 17828 16516
rect 7564 16396 7616 16448
rect 9956 16396 10008 16448
rect 10048 16439 10100 16448
rect 10048 16405 10057 16439
rect 10057 16405 10091 16439
rect 10091 16405 10100 16439
rect 10048 16396 10100 16405
rect 11612 16396 11664 16448
rect 13544 16396 13596 16448
rect 16764 16396 16816 16448
rect 17684 16396 17736 16448
rect 17960 16439 18012 16448
rect 17960 16405 17969 16439
rect 17969 16405 18003 16439
rect 18003 16405 18012 16439
rect 17960 16396 18012 16405
rect 24584 16396 24636 16448
rect 3756 16294 3808 16346
rect 3820 16294 3872 16346
rect 3884 16294 3936 16346
rect 3948 16294 4000 16346
rect 4012 16294 4064 16346
rect 10472 16294 10524 16346
rect 10536 16294 10588 16346
rect 10600 16294 10652 16346
rect 10664 16294 10716 16346
rect 10728 16294 10780 16346
rect 17188 16294 17240 16346
rect 17252 16294 17304 16346
rect 17316 16294 17368 16346
rect 17380 16294 17432 16346
rect 17444 16294 17496 16346
rect 23904 16294 23956 16346
rect 23968 16294 24020 16346
rect 24032 16294 24084 16346
rect 24096 16294 24148 16346
rect 24160 16294 24212 16346
rect 5540 16192 5592 16244
rect 6828 16192 6880 16244
rect 4804 16124 4856 16176
rect 6644 16124 6696 16176
rect 8116 16192 8168 16244
rect 8668 16235 8720 16244
rect 8668 16201 8677 16235
rect 8677 16201 8711 16235
rect 8711 16201 8720 16235
rect 8668 16192 8720 16201
rect 8944 16192 8996 16244
rect 11704 16192 11756 16244
rect 13912 16235 13964 16244
rect 13912 16201 13921 16235
rect 13921 16201 13955 16235
rect 13955 16201 13964 16235
rect 13912 16192 13964 16201
rect 18512 16235 18564 16244
rect 18512 16201 18521 16235
rect 18521 16201 18555 16235
rect 18555 16201 18564 16235
rect 18512 16192 18564 16201
rect 20812 16192 20864 16244
rect 16672 16124 16724 16176
rect 3240 16099 3292 16108
rect 3240 16065 3249 16099
rect 3249 16065 3283 16099
rect 3283 16065 3292 16099
rect 3240 16056 3292 16065
rect 3332 15988 3384 16040
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 5632 16031 5684 16040
rect 5632 15997 5641 16031
rect 5641 15997 5675 16031
rect 5675 15997 5684 16031
rect 5632 15988 5684 15997
rect 6276 16031 6328 16040
rect 6276 15997 6285 16031
rect 6285 15997 6319 16031
rect 6319 15997 6328 16031
rect 6276 15988 6328 15997
rect 8024 16056 8076 16108
rect 8760 16056 8812 16108
rect 8300 15988 8352 16040
rect 9680 16056 9732 16108
rect 10232 16099 10284 16108
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 11980 16056 12032 16108
rect 7472 15920 7524 15972
rect 11612 15988 11664 16040
rect 13084 16056 13136 16108
rect 15292 16056 15344 16108
rect 15752 16056 15804 16108
rect 16580 15988 16632 16040
rect 16948 16056 17000 16108
rect 17040 16056 17092 16108
rect 16856 15988 16908 16040
rect 17316 15988 17368 16040
rect 9312 15920 9364 15972
rect 10324 15920 10376 15972
rect 11520 15920 11572 15972
rect 11980 15963 12032 15972
rect 11980 15929 11989 15963
rect 11989 15929 12023 15963
rect 12023 15929 12032 15963
rect 11980 15920 12032 15929
rect 12164 15920 12216 15972
rect 15016 15963 15068 15972
rect 15016 15929 15025 15963
rect 15025 15929 15059 15963
rect 15059 15929 15068 15963
rect 15016 15920 15068 15929
rect 17592 16031 17644 16040
rect 17592 15997 17601 16031
rect 17601 15997 17635 16031
rect 17635 15997 17644 16031
rect 17592 15988 17644 15997
rect 17776 15988 17828 16040
rect 18144 16056 18196 16108
rect 19616 16031 19668 16040
rect 19616 15997 19625 16031
rect 19625 15997 19659 16031
rect 19659 15997 19668 16031
rect 19616 15988 19668 15997
rect 5908 15852 5960 15904
rect 12256 15895 12308 15904
rect 12256 15861 12265 15895
rect 12265 15861 12299 15895
rect 12299 15861 12308 15895
rect 12256 15852 12308 15861
rect 13176 15852 13228 15904
rect 13728 15852 13780 15904
rect 14464 15852 14516 15904
rect 16212 15895 16264 15904
rect 16212 15861 16221 15895
rect 16221 15861 16255 15895
rect 16255 15861 16264 15895
rect 16212 15852 16264 15861
rect 16948 15895 17000 15904
rect 16948 15861 16957 15895
rect 16957 15861 16991 15895
rect 16991 15861 17000 15895
rect 18880 15920 18932 15972
rect 19340 15920 19392 15972
rect 20444 15988 20496 16040
rect 23572 16192 23624 16244
rect 25964 16124 26016 16176
rect 23664 16056 23716 16108
rect 23020 16031 23072 16040
rect 23020 15997 23029 16031
rect 23029 15997 23063 16031
rect 23063 15997 23072 16031
rect 23020 15988 23072 15997
rect 23112 15988 23164 16040
rect 26608 15988 26660 16040
rect 16948 15852 17000 15861
rect 17868 15852 17920 15904
rect 21272 15852 21324 15904
rect 22744 15895 22796 15904
rect 22744 15861 22753 15895
rect 22753 15861 22787 15895
rect 22787 15861 22796 15895
rect 22744 15852 22796 15861
rect 23664 15852 23716 15904
rect 7114 15750 7166 15802
rect 7178 15750 7230 15802
rect 7242 15750 7294 15802
rect 7306 15750 7358 15802
rect 7370 15750 7422 15802
rect 13830 15750 13882 15802
rect 13894 15750 13946 15802
rect 13958 15750 14010 15802
rect 14022 15750 14074 15802
rect 14086 15750 14138 15802
rect 20546 15750 20598 15802
rect 20610 15750 20662 15802
rect 20674 15750 20726 15802
rect 20738 15750 20790 15802
rect 20802 15750 20854 15802
rect 27262 15750 27314 15802
rect 27326 15750 27378 15802
rect 27390 15750 27442 15802
rect 27454 15750 27506 15802
rect 27518 15750 27570 15802
rect 3332 15691 3384 15700
rect 3332 15657 3341 15691
rect 3341 15657 3375 15691
rect 3375 15657 3384 15691
rect 3332 15648 3384 15657
rect 6276 15648 6328 15700
rect 7472 15648 7524 15700
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 13176 15691 13228 15700
rect 13176 15657 13185 15691
rect 13185 15657 13219 15691
rect 13219 15657 13228 15691
rect 13176 15648 13228 15657
rect 13544 15691 13596 15700
rect 13544 15657 13553 15691
rect 13553 15657 13587 15691
rect 13587 15657 13596 15691
rect 13544 15648 13596 15657
rect 14464 15691 14516 15700
rect 14464 15657 14473 15691
rect 14473 15657 14507 15691
rect 14507 15657 14516 15691
rect 14464 15648 14516 15657
rect 15936 15648 15988 15700
rect 4988 15580 5040 15632
rect 5540 15580 5592 15632
rect 3608 15444 3660 15496
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 4804 15555 4856 15564
rect 4804 15521 4813 15555
rect 4813 15521 4847 15555
rect 4847 15521 4856 15555
rect 4804 15512 4856 15521
rect 4988 15376 5040 15428
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 8024 15580 8076 15632
rect 8116 15580 8168 15632
rect 15292 15623 15344 15632
rect 15292 15589 15301 15623
rect 15301 15589 15335 15623
rect 15335 15589 15344 15623
rect 15292 15580 15344 15589
rect 17868 15580 17920 15632
rect 5908 15512 5960 15564
rect 7564 15555 7616 15564
rect 7564 15521 7573 15555
rect 7573 15521 7607 15555
rect 7607 15521 7616 15555
rect 7564 15512 7616 15521
rect 4804 15308 4856 15360
rect 5356 15308 5408 15360
rect 7932 15555 7984 15564
rect 7932 15521 7941 15555
rect 7941 15521 7975 15555
rect 7975 15521 7984 15555
rect 7932 15512 7984 15521
rect 11796 15555 11848 15564
rect 11796 15521 11805 15555
rect 11805 15521 11839 15555
rect 11839 15521 11848 15555
rect 11796 15512 11848 15521
rect 11980 15512 12032 15564
rect 12808 15512 12860 15564
rect 9588 15487 9640 15496
rect 9588 15453 9597 15487
rect 9597 15453 9631 15487
rect 9631 15453 9640 15487
rect 9588 15444 9640 15453
rect 11244 15444 11296 15496
rect 12164 15444 12216 15496
rect 10968 15376 11020 15428
rect 14096 15444 14148 15496
rect 14924 15444 14976 15496
rect 15660 15555 15712 15564
rect 15660 15521 15669 15555
rect 15669 15521 15703 15555
rect 15703 15521 15712 15555
rect 15660 15512 15712 15521
rect 16212 15512 16264 15564
rect 16764 15555 16816 15564
rect 16764 15521 16773 15555
rect 16773 15521 16807 15555
rect 16807 15521 16816 15555
rect 16764 15512 16816 15521
rect 17776 15555 17828 15564
rect 17776 15521 17785 15555
rect 17785 15521 17819 15555
rect 17819 15521 17828 15555
rect 17776 15512 17828 15521
rect 18604 15555 18656 15564
rect 18604 15521 18613 15555
rect 18613 15521 18647 15555
rect 18647 15521 18656 15555
rect 18604 15512 18656 15521
rect 23112 15648 23164 15700
rect 23204 15691 23256 15700
rect 23204 15657 23213 15691
rect 23213 15657 23247 15691
rect 23247 15657 23256 15691
rect 23204 15648 23256 15657
rect 21088 15512 21140 15564
rect 22100 15555 22152 15564
rect 22100 15521 22134 15555
rect 22134 15521 22152 15555
rect 22100 15512 22152 15521
rect 23204 15512 23256 15564
rect 25228 15580 25280 15632
rect 24768 15512 24820 15564
rect 18236 15444 18288 15496
rect 19524 15444 19576 15496
rect 17040 15376 17092 15428
rect 19064 15376 19116 15428
rect 22836 15376 22888 15428
rect 8760 15308 8812 15360
rect 11152 15308 11204 15360
rect 16396 15308 16448 15360
rect 19892 15308 19944 15360
rect 20444 15308 20496 15360
rect 21088 15351 21140 15360
rect 21088 15317 21097 15351
rect 21097 15317 21131 15351
rect 21131 15317 21140 15351
rect 21088 15308 21140 15317
rect 25044 15308 25096 15360
rect 3756 15206 3808 15258
rect 3820 15206 3872 15258
rect 3884 15206 3936 15258
rect 3948 15206 4000 15258
rect 4012 15206 4064 15258
rect 10472 15206 10524 15258
rect 10536 15206 10588 15258
rect 10600 15206 10652 15258
rect 10664 15206 10716 15258
rect 10728 15206 10780 15258
rect 17188 15206 17240 15258
rect 17252 15206 17304 15258
rect 17316 15206 17368 15258
rect 17380 15206 17432 15258
rect 17444 15206 17496 15258
rect 23904 15206 23956 15258
rect 23968 15206 24020 15258
rect 24032 15206 24084 15258
rect 24096 15206 24148 15258
rect 24160 15206 24212 15258
rect 6000 15104 6052 15156
rect 8300 15104 8352 15156
rect 10324 15104 10376 15156
rect 12716 15104 12768 15156
rect 12992 15104 13044 15156
rect 18604 15104 18656 15156
rect 18696 15104 18748 15156
rect 23756 15104 23808 15156
rect 24768 15147 24820 15156
rect 24768 15113 24777 15147
rect 24777 15113 24811 15147
rect 24811 15113 24820 15147
rect 24768 15104 24820 15113
rect 4068 14900 4120 14952
rect 4804 14943 4856 14952
rect 4804 14909 4813 14943
rect 4813 14909 4847 14943
rect 4847 14909 4856 14943
rect 4804 14900 4856 14909
rect 5448 14943 5500 14952
rect 5448 14909 5457 14943
rect 5457 14909 5491 14943
rect 5491 14909 5500 14943
rect 5448 14900 5500 14909
rect 5080 14875 5132 14884
rect 5080 14841 5089 14875
rect 5089 14841 5123 14875
rect 5123 14841 5132 14875
rect 5080 14832 5132 14841
rect 5632 14900 5684 14952
rect 6460 15036 6512 15088
rect 7932 15036 7984 15088
rect 9036 15036 9088 15088
rect 11704 15036 11756 15088
rect 13728 15036 13780 15088
rect 15568 15036 15620 15088
rect 16304 15036 16356 15088
rect 16396 15036 16448 15088
rect 13176 15011 13228 15020
rect 13176 14977 13185 15011
rect 13185 14977 13219 15011
rect 13219 14977 13228 15011
rect 13176 14968 13228 14977
rect 13820 14968 13872 15020
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 6368 14943 6420 14952
rect 6368 14909 6377 14943
rect 6377 14909 6411 14943
rect 6411 14909 6420 14943
rect 6368 14900 6420 14909
rect 8944 14900 8996 14952
rect 9588 14943 9640 14952
rect 9588 14909 9597 14943
rect 9597 14909 9631 14943
rect 9631 14909 9640 14943
rect 9588 14900 9640 14909
rect 10048 14943 10100 14952
rect 10048 14909 10057 14943
rect 10057 14909 10091 14943
rect 10091 14909 10100 14943
rect 10048 14900 10100 14909
rect 10968 14943 11020 14952
rect 10968 14909 10977 14943
rect 10977 14909 11011 14943
rect 11011 14909 11020 14943
rect 10968 14900 11020 14909
rect 8576 14764 8628 14816
rect 8668 14807 8720 14816
rect 8668 14773 8677 14807
rect 8677 14773 8711 14807
rect 8711 14773 8720 14807
rect 8668 14764 8720 14773
rect 8760 14764 8812 14816
rect 11152 14943 11204 14952
rect 11152 14909 11161 14943
rect 11161 14909 11195 14943
rect 11195 14909 11204 14943
rect 11152 14900 11204 14909
rect 11704 14900 11756 14952
rect 12072 14943 12124 14952
rect 12072 14909 12081 14943
rect 12081 14909 12115 14943
rect 12115 14909 12124 14943
rect 12072 14900 12124 14909
rect 12256 14943 12308 14952
rect 12256 14909 12265 14943
rect 12265 14909 12299 14943
rect 12299 14909 12308 14943
rect 12256 14900 12308 14909
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 12808 14900 12860 14952
rect 14464 14968 14516 15020
rect 17224 14968 17276 15020
rect 18144 15079 18196 15088
rect 18144 15045 18153 15079
rect 18153 15045 18187 15079
rect 18187 15045 18196 15079
rect 18144 15036 18196 15045
rect 19708 15036 19760 15088
rect 25412 15036 25464 15088
rect 11428 14832 11480 14884
rect 15660 14900 15712 14952
rect 15936 14900 15988 14952
rect 16304 14943 16356 14952
rect 16304 14909 16313 14943
rect 16313 14909 16347 14943
rect 16347 14909 16356 14943
rect 16304 14900 16356 14909
rect 16396 14943 16448 14952
rect 16396 14909 16405 14943
rect 16405 14909 16439 14943
rect 16439 14909 16448 14943
rect 16396 14900 16448 14909
rect 17040 14900 17092 14952
rect 17592 14968 17644 15020
rect 18328 14943 18380 14952
rect 18328 14909 18337 14943
rect 18337 14909 18371 14943
rect 18371 14909 18380 14943
rect 18328 14900 18380 14909
rect 19524 14900 19576 14952
rect 24032 14943 24084 14952
rect 24032 14909 24041 14943
rect 24041 14909 24075 14943
rect 24075 14909 24084 14943
rect 24032 14900 24084 14909
rect 24492 14968 24544 15020
rect 13912 14875 13964 14884
rect 13912 14841 13921 14875
rect 13921 14841 13955 14875
rect 13955 14841 13964 14875
rect 13912 14832 13964 14841
rect 16948 14832 17000 14884
rect 16028 14764 16080 14816
rect 17132 14764 17184 14816
rect 17408 14875 17460 14884
rect 17408 14841 17417 14875
rect 17417 14841 17451 14875
rect 17451 14841 17460 14875
rect 17408 14832 17460 14841
rect 17776 14764 17828 14816
rect 24860 14900 24912 14952
rect 24952 14943 25004 14952
rect 24952 14909 24961 14943
rect 24961 14909 24995 14943
rect 24995 14909 25004 14943
rect 24952 14900 25004 14909
rect 19064 14764 19116 14816
rect 21088 14764 21140 14816
rect 21456 14764 21508 14816
rect 23940 14764 23992 14816
rect 24400 14764 24452 14816
rect 24676 14832 24728 14884
rect 25044 14764 25096 14816
rect 7114 14662 7166 14714
rect 7178 14662 7230 14714
rect 7242 14662 7294 14714
rect 7306 14662 7358 14714
rect 7370 14662 7422 14714
rect 13830 14662 13882 14714
rect 13894 14662 13946 14714
rect 13958 14662 14010 14714
rect 14022 14662 14074 14714
rect 14086 14662 14138 14714
rect 20546 14662 20598 14714
rect 20610 14662 20662 14714
rect 20674 14662 20726 14714
rect 20738 14662 20790 14714
rect 20802 14662 20854 14714
rect 27262 14662 27314 14714
rect 27326 14662 27378 14714
rect 27390 14662 27442 14714
rect 27454 14662 27506 14714
rect 27518 14662 27570 14714
rect 4528 14560 4580 14612
rect 6368 14560 6420 14612
rect 8944 14603 8996 14612
rect 8944 14569 8953 14603
rect 8953 14569 8987 14603
rect 8987 14569 8996 14603
rect 8944 14560 8996 14569
rect 9404 14560 9456 14612
rect 9956 14560 10008 14612
rect 10324 14560 10376 14612
rect 12348 14603 12400 14612
rect 12348 14569 12357 14603
rect 12357 14569 12391 14603
rect 12391 14569 12400 14603
rect 12348 14560 12400 14569
rect 14188 14560 14240 14612
rect 18328 14560 18380 14612
rect 4988 14492 5040 14544
rect 2596 14467 2648 14476
rect 2596 14433 2630 14467
rect 2630 14433 2648 14467
rect 2596 14424 2648 14433
rect 4068 14356 4120 14408
rect 3332 14288 3384 14340
rect 2504 14220 2556 14272
rect 3608 14220 3660 14272
rect 4436 14424 4488 14476
rect 4896 14467 4948 14476
rect 4896 14433 4905 14467
rect 4905 14433 4939 14467
rect 4939 14433 4948 14467
rect 4896 14424 4948 14433
rect 5264 14424 5316 14476
rect 6920 14492 6972 14544
rect 8024 14492 8076 14544
rect 8576 14492 8628 14544
rect 10140 14492 10192 14544
rect 17684 14492 17736 14544
rect 19432 14492 19484 14544
rect 22100 14560 22152 14612
rect 24952 14560 25004 14612
rect 5080 14356 5132 14408
rect 8392 14424 8444 14476
rect 9588 14356 9640 14408
rect 10232 14399 10284 14408
rect 10232 14365 10241 14399
rect 10241 14365 10275 14399
rect 10275 14365 10284 14399
rect 10232 14356 10284 14365
rect 11428 14356 11480 14408
rect 11796 14356 11848 14408
rect 13176 14356 13228 14408
rect 7840 14220 7892 14272
rect 8852 14220 8904 14272
rect 12440 14220 12492 14272
rect 15200 14424 15252 14476
rect 16120 14424 16172 14476
rect 17132 14467 17184 14476
rect 17132 14433 17141 14467
rect 17141 14433 17175 14467
rect 17175 14433 17184 14467
rect 17132 14424 17184 14433
rect 17224 14424 17276 14476
rect 17868 14424 17920 14476
rect 18236 14467 18288 14476
rect 18236 14433 18245 14467
rect 18245 14433 18279 14467
rect 18279 14433 18288 14467
rect 18236 14424 18288 14433
rect 18328 14467 18380 14476
rect 18328 14433 18337 14467
rect 18337 14433 18371 14467
rect 18371 14433 18380 14467
rect 18328 14424 18380 14433
rect 13544 14356 13596 14408
rect 13728 14399 13780 14408
rect 13728 14365 13737 14399
rect 13737 14365 13771 14399
rect 13771 14365 13780 14399
rect 13728 14356 13780 14365
rect 14740 14356 14792 14408
rect 15108 14399 15160 14408
rect 15108 14365 15117 14399
rect 15117 14365 15151 14399
rect 15151 14365 15160 14399
rect 15108 14356 15160 14365
rect 16856 14288 16908 14340
rect 21180 14424 21232 14476
rect 22192 14467 22244 14476
rect 22192 14433 22201 14467
rect 22201 14433 22235 14467
rect 22235 14433 22244 14467
rect 22192 14424 22244 14433
rect 23940 14535 23992 14544
rect 22376 14424 22428 14476
rect 22836 14424 22888 14476
rect 23940 14501 23949 14535
rect 23949 14501 23983 14535
rect 23983 14501 23992 14535
rect 23940 14492 23992 14501
rect 25228 14492 25280 14544
rect 19524 14399 19576 14408
rect 19524 14365 19533 14399
rect 19533 14365 19567 14399
rect 19567 14365 19576 14399
rect 19524 14356 19576 14365
rect 14648 14220 14700 14272
rect 15844 14220 15896 14272
rect 15936 14220 15988 14272
rect 19432 14220 19484 14272
rect 23296 14467 23348 14476
rect 23296 14433 23305 14467
rect 23305 14433 23339 14467
rect 23339 14433 23348 14467
rect 23296 14424 23348 14433
rect 24492 14424 24544 14476
rect 25504 14424 25556 14476
rect 24032 14356 24084 14408
rect 23296 14288 23348 14340
rect 19800 14220 19852 14272
rect 20904 14263 20956 14272
rect 20904 14229 20913 14263
rect 20913 14229 20947 14263
rect 20947 14229 20956 14263
rect 20904 14220 20956 14229
rect 23664 14220 23716 14272
rect 24676 14288 24728 14340
rect 25596 14220 25648 14272
rect 3756 14118 3808 14170
rect 3820 14118 3872 14170
rect 3884 14118 3936 14170
rect 3948 14118 4000 14170
rect 4012 14118 4064 14170
rect 10472 14118 10524 14170
rect 10536 14118 10588 14170
rect 10600 14118 10652 14170
rect 10664 14118 10716 14170
rect 10728 14118 10780 14170
rect 17188 14118 17240 14170
rect 17252 14118 17304 14170
rect 17316 14118 17368 14170
rect 17380 14118 17432 14170
rect 17444 14118 17496 14170
rect 23904 14118 23956 14170
rect 23968 14118 24020 14170
rect 24032 14118 24084 14170
rect 24096 14118 24148 14170
rect 24160 14118 24212 14170
rect 2596 14016 2648 14068
rect 4988 14016 5040 14068
rect 9496 14016 9548 14068
rect 4252 13948 4304 14000
rect 8392 13991 8444 14000
rect 8392 13957 8401 13991
rect 8401 13957 8435 13991
rect 8435 13957 8444 13991
rect 8392 13948 8444 13957
rect 9128 13991 9180 14000
rect 9128 13957 9137 13991
rect 9137 13957 9171 13991
rect 9171 13957 9180 13991
rect 9128 13948 9180 13957
rect 2504 13880 2556 13932
rect 3332 13812 3384 13864
rect 5264 13923 5316 13932
rect 5264 13889 5273 13923
rect 5273 13889 5307 13923
rect 5307 13889 5316 13923
rect 5264 13880 5316 13889
rect 5448 13880 5500 13932
rect 5632 13855 5684 13864
rect 5632 13821 5641 13855
rect 5641 13821 5675 13855
rect 5675 13821 5684 13855
rect 5632 13812 5684 13821
rect 5724 13855 5776 13864
rect 5724 13821 5733 13855
rect 5733 13821 5767 13855
rect 5767 13821 5776 13855
rect 5724 13812 5776 13821
rect 5816 13855 5868 13864
rect 5816 13821 5825 13855
rect 5825 13821 5859 13855
rect 5859 13821 5868 13855
rect 5816 13812 5868 13821
rect 6460 13812 6512 13864
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 7840 13812 7892 13821
rect 8024 13855 8076 13864
rect 8024 13821 8033 13855
rect 8033 13821 8067 13855
rect 8067 13821 8076 13855
rect 8024 13812 8076 13821
rect 8668 13855 8720 13864
rect 8668 13821 8677 13855
rect 8677 13821 8711 13855
rect 8711 13821 8720 13855
rect 8668 13812 8720 13821
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 8760 13812 8812 13821
rect 8852 13855 8904 13864
rect 8852 13821 8861 13855
rect 8861 13821 8895 13855
rect 8895 13821 8904 13855
rect 8852 13812 8904 13821
rect 9036 13855 9088 13864
rect 9036 13821 9045 13855
rect 9045 13821 9079 13855
rect 9079 13821 9088 13855
rect 9036 13812 9088 13821
rect 9956 13948 10008 14000
rect 11336 14016 11388 14068
rect 12624 14016 12676 14068
rect 14740 14059 14792 14068
rect 14740 14025 14749 14059
rect 14749 14025 14783 14059
rect 14783 14025 14792 14059
rect 14740 14016 14792 14025
rect 14924 14016 14976 14068
rect 11520 13948 11572 14000
rect 15200 13948 15252 14000
rect 9588 13880 9640 13932
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 10324 13880 10376 13932
rect 9404 13855 9456 13864
rect 9404 13821 9413 13855
rect 9413 13821 9447 13855
rect 9447 13821 9456 13855
rect 9404 13812 9456 13821
rect 9496 13855 9548 13864
rect 9496 13821 9505 13855
rect 9505 13821 9539 13855
rect 9539 13821 9548 13855
rect 9496 13812 9548 13821
rect 8208 13787 8260 13796
rect 8208 13753 8217 13787
rect 8217 13753 8251 13787
rect 8251 13753 8260 13787
rect 8208 13744 8260 13753
rect 10232 13812 10284 13864
rect 10140 13744 10192 13796
rect 4712 13676 4764 13728
rect 11796 13812 11848 13864
rect 12992 13880 13044 13932
rect 13268 13880 13320 13932
rect 15108 13880 15160 13932
rect 16304 14016 16356 14068
rect 17132 14016 17184 14068
rect 16396 13948 16448 14000
rect 17316 13948 17368 14000
rect 11428 13676 11480 13728
rect 16028 13880 16080 13932
rect 18328 14016 18380 14068
rect 20904 14016 20956 14068
rect 21180 14059 21232 14068
rect 21180 14025 21189 14059
rect 21189 14025 21223 14059
rect 21223 14025 21232 14059
rect 21180 14016 21232 14025
rect 22376 14016 22428 14068
rect 23480 14016 23532 14068
rect 24032 14016 24084 14068
rect 15844 13812 15896 13864
rect 16672 13744 16724 13796
rect 16856 13812 16908 13864
rect 17316 13855 17368 13864
rect 17316 13821 17325 13855
rect 17325 13821 17359 13855
rect 17359 13821 17368 13855
rect 17316 13812 17368 13821
rect 17132 13787 17184 13796
rect 17132 13753 17141 13787
rect 17141 13753 17175 13787
rect 17175 13753 17184 13787
rect 17132 13744 17184 13753
rect 18236 13812 18288 13864
rect 18696 13855 18748 13864
rect 18696 13821 18705 13855
rect 18705 13821 18739 13855
rect 18739 13821 18748 13855
rect 18696 13812 18748 13821
rect 19800 13855 19852 13864
rect 19800 13821 19809 13855
rect 19809 13821 19843 13855
rect 19843 13821 19852 13855
rect 19800 13812 19852 13821
rect 21364 13880 21416 13932
rect 21916 13923 21968 13932
rect 21916 13889 21925 13923
rect 21925 13889 21959 13923
rect 21959 13889 21968 13923
rect 21916 13880 21968 13889
rect 22376 13923 22428 13932
rect 22376 13889 22385 13923
rect 22385 13889 22419 13923
rect 22419 13889 22428 13923
rect 22376 13880 22428 13889
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 25412 14059 25464 14068
rect 25412 14025 25421 14059
rect 25421 14025 25455 14059
rect 25455 14025 25464 14059
rect 25412 14016 25464 14025
rect 25504 14059 25556 14068
rect 25504 14025 25513 14059
rect 25513 14025 25547 14059
rect 25547 14025 25556 14059
rect 25504 14016 25556 14025
rect 25596 14016 25648 14068
rect 25780 13880 25832 13932
rect 21272 13855 21324 13864
rect 21272 13821 21281 13855
rect 21281 13821 21315 13855
rect 21315 13821 21324 13855
rect 21272 13812 21324 13821
rect 21456 13855 21508 13864
rect 21456 13821 21465 13855
rect 21465 13821 21499 13855
rect 21499 13821 21508 13855
rect 21456 13812 21508 13821
rect 21548 13812 21600 13864
rect 23296 13812 23348 13864
rect 17776 13787 17828 13796
rect 17776 13753 17785 13787
rect 17785 13753 17819 13787
rect 17819 13753 17828 13787
rect 17776 13744 17828 13753
rect 17868 13787 17920 13796
rect 17868 13753 17877 13787
rect 17877 13753 17911 13787
rect 17911 13753 17920 13787
rect 17868 13744 17920 13753
rect 24860 13744 24912 13796
rect 25136 13812 25188 13864
rect 25412 13812 25464 13864
rect 25872 13855 25924 13864
rect 25872 13821 25881 13855
rect 25881 13821 25915 13855
rect 25915 13821 25924 13855
rect 25872 13812 25924 13821
rect 25596 13744 25648 13796
rect 12256 13676 12308 13728
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 14188 13719 14240 13728
rect 14188 13685 14197 13719
rect 14197 13685 14231 13719
rect 14231 13685 14240 13719
rect 14188 13676 14240 13685
rect 14372 13676 14424 13728
rect 16120 13676 16172 13728
rect 7114 13574 7166 13626
rect 7178 13574 7230 13626
rect 7242 13574 7294 13626
rect 7306 13574 7358 13626
rect 7370 13574 7422 13626
rect 13830 13574 13882 13626
rect 13894 13574 13946 13626
rect 13958 13574 14010 13626
rect 14022 13574 14074 13626
rect 14086 13574 14138 13626
rect 20546 13574 20598 13626
rect 20610 13574 20662 13626
rect 20674 13574 20726 13626
rect 20738 13574 20790 13626
rect 20802 13574 20854 13626
rect 27262 13574 27314 13626
rect 27326 13574 27378 13626
rect 27390 13574 27442 13626
rect 27454 13574 27506 13626
rect 27518 13574 27570 13626
rect 5632 13472 5684 13524
rect 9864 13472 9916 13524
rect 10140 13472 10192 13524
rect 12440 13472 12492 13524
rect 13452 13515 13504 13524
rect 13452 13481 13461 13515
rect 13461 13481 13495 13515
rect 13495 13481 13504 13515
rect 13452 13472 13504 13481
rect 14188 13472 14240 13524
rect 24860 13472 24912 13524
rect 25872 13472 25924 13524
rect 4252 13404 4304 13456
rect 4436 13268 4488 13320
rect 4712 13379 4764 13388
rect 4712 13345 4721 13379
rect 4721 13345 4755 13379
rect 4755 13345 4764 13379
rect 4712 13336 4764 13345
rect 9680 13404 9732 13456
rect 9956 13404 10008 13456
rect 11888 13404 11940 13456
rect 8392 13336 8444 13388
rect 10232 13336 10284 13388
rect 11060 13336 11112 13388
rect 12440 13379 12492 13388
rect 12440 13345 12449 13379
rect 12449 13345 12483 13379
rect 12483 13345 12492 13379
rect 12440 13336 12492 13345
rect 4896 13268 4948 13320
rect 4988 13268 5040 13320
rect 8760 13268 8812 13320
rect 4160 13175 4212 13184
rect 4160 13141 4169 13175
rect 4169 13141 4203 13175
rect 4203 13141 4212 13175
rect 4160 13132 4212 13141
rect 6092 13132 6144 13184
rect 7932 13132 7984 13184
rect 9404 13268 9456 13320
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 12624 13379 12676 13388
rect 12624 13345 12633 13379
rect 12633 13345 12667 13379
rect 12667 13345 12676 13379
rect 12624 13336 12676 13345
rect 12348 13243 12400 13252
rect 12348 13209 12357 13243
rect 12357 13209 12391 13243
rect 12391 13209 12400 13243
rect 13544 13404 13596 13456
rect 15200 13336 15252 13388
rect 16120 13379 16172 13388
rect 16120 13345 16129 13379
rect 16129 13345 16163 13379
rect 16163 13345 16172 13379
rect 16120 13336 16172 13345
rect 16304 13447 16356 13456
rect 16304 13413 16313 13447
rect 16313 13413 16347 13447
rect 16347 13413 16356 13447
rect 16304 13404 16356 13413
rect 16672 13404 16724 13456
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 21548 13404 21600 13456
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 14556 13268 14608 13320
rect 15108 13311 15160 13320
rect 15108 13277 15117 13311
rect 15117 13277 15151 13311
rect 15151 13277 15160 13311
rect 15108 13268 15160 13277
rect 12348 13200 12400 13209
rect 16580 13200 16632 13252
rect 20904 13336 20956 13388
rect 24032 13379 24084 13388
rect 24032 13345 24041 13379
rect 24041 13345 24075 13379
rect 24075 13345 24084 13379
rect 24032 13336 24084 13345
rect 25044 13379 25096 13388
rect 25044 13345 25053 13379
rect 25053 13345 25087 13379
rect 25087 13345 25096 13379
rect 25044 13336 25096 13345
rect 17868 13268 17920 13320
rect 21272 13268 21324 13320
rect 18696 13200 18748 13252
rect 21088 13200 21140 13252
rect 22284 13268 22336 13320
rect 22560 13268 22612 13320
rect 23756 13268 23808 13320
rect 24308 13268 24360 13320
rect 24952 13268 25004 13320
rect 25412 13379 25464 13388
rect 25412 13345 25421 13379
rect 25421 13345 25455 13379
rect 25455 13345 25464 13379
rect 25412 13336 25464 13345
rect 25780 13336 25832 13388
rect 25320 13268 25372 13320
rect 25872 13200 25924 13252
rect 11336 13132 11388 13184
rect 12716 13132 12768 13184
rect 15936 13132 15988 13184
rect 24768 13132 24820 13184
rect 24952 13175 25004 13184
rect 24952 13141 24961 13175
rect 24961 13141 24995 13175
rect 24995 13141 25004 13175
rect 24952 13132 25004 13141
rect 25780 13175 25832 13184
rect 25780 13141 25789 13175
rect 25789 13141 25823 13175
rect 25823 13141 25832 13175
rect 25780 13132 25832 13141
rect 3756 13030 3808 13082
rect 3820 13030 3872 13082
rect 3884 13030 3936 13082
rect 3948 13030 4000 13082
rect 4012 13030 4064 13082
rect 10472 13030 10524 13082
rect 10536 13030 10588 13082
rect 10600 13030 10652 13082
rect 10664 13030 10716 13082
rect 10728 13030 10780 13082
rect 17188 13030 17240 13082
rect 17252 13030 17304 13082
rect 17316 13030 17368 13082
rect 17380 13030 17432 13082
rect 17444 13030 17496 13082
rect 23904 13030 23956 13082
rect 23968 13030 24020 13082
rect 24032 13030 24084 13082
rect 24096 13030 24148 13082
rect 24160 13030 24212 13082
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 6920 12971 6972 12980
rect 6920 12937 6929 12971
rect 6929 12937 6963 12971
rect 6963 12937 6972 12971
rect 6920 12928 6972 12937
rect 8392 12971 8444 12980
rect 8392 12937 8401 12971
rect 8401 12937 8435 12971
rect 8435 12937 8444 12971
rect 8392 12928 8444 12937
rect 11060 12928 11112 12980
rect 12440 12928 12492 12980
rect 13452 12928 13504 12980
rect 16120 12928 16172 12980
rect 17684 12928 17736 12980
rect 3608 12767 3660 12776
rect 3608 12733 3617 12767
rect 3617 12733 3651 12767
rect 3651 12733 3660 12767
rect 3608 12724 3660 12733
rect 4160 12792 4212 12844
rect 3976 12767 4028 12776
rect 3976 12733 3985 12767
rect 3985 12733 4019 12767
rect 4019 12733 4028 12767
rect 3976 12724 4028 12733
rect 4436 12767 4488 12776
rect 4436 12733 4445 12767
rect 4445 12733 4479 12767
rect 4479 12733 4488 12767
rect 4436 12724 4488 12733
rect 5356 12724 5408 12776
rect 15200 12860 15252 12912
rect 17500 12860 17552 12912
rect 20444 12928 20496 12980
rect 23756 12928 23808 12980
rect 18604 12860 18656 12912
rect 8208 12792 8260 12844
rect 9404 12792 9456 12844
rect 2780 12588 2832 12640
rect 3240 12631 3292 12640
rect 3240 12597 3249 12631
rect 3249 12597 3283 12631
rect 3283 12597 3292 12631
rect 3240 12588 3292 12597
rect 4896 12656 4948 12708
rect 5816 12656 5868 12708
rect 8208 12699 8260 12708
rect 8208 12665 8217 12699
rect 8217 12665 8251 12699
rect 8251 12665 8260 12699
rect 8208 12656 8260 12665
rect 9588 12724 9640 12776
rect 9956 12724 10008 12776
rect 9956 12588 10008 12640
rect 10508 12767 10560 12776
rect 10508 12733 10517 12767
rect 10517 12733 10551 12767
rect 10551 12733 10560 12767
rect 10508 12724 10560 12733
rect 11336 12767 11388 12776
rect 11336 12733 11345 12767
rect 11345 12733 11379 12767
rect 11379 12733 11388 12767
rect 11336 12724 11388 12733
rect 11428 12767 11480 12776
rect 11428 12733 11437 12767
rect 11437 12733 11471 12767
rect 11471 12733 11480 12767
rect 11428 12724 11480 12733
rect 11704 12724 11756 12776
rect 12348 12835 12400 12844
rect 12348 12801 12357 12835
rect 12357 12801 12391 12835
rect 12391 12801 12400 12835
rect 12348 12792 12400 12801
rect 12532 12835 12584 12844
rect 12532 12801 12541 12835
rect 12541 12801 12575 12835
rect 12575 12801 12584 12835
rect 12532 12792 12584 12801
rect 23480 12860 23532 12912
rect 24952 12928 25004 12980
rect 25044 12860 25096 12912
rect 25412 12860 25464 12912
rect 12716 12767 12768 12776
rect 12716 12733 12725 12767
rect 12725 12733 12759 12767
rect 12759 12733 12768 12767
rect 12716 12724 12768 12733
rect 15108 12724 15160 12776
rect 15936 12767 15988 12776
rect 15936 12733 15945 12767
rect 15945 12733 15979 12767
rect 15979 12733 15988 12767
rect 15936 12724 15988 12733
rect 16304 12724 16356 12776
rect 14372 12656 14424 12708
rect 10140 12631 10192 12640
rect 10140 12597 10149 12631
rect 10149 12597 10183 12631
rect 10183 12597 10192 12631
rect 10140 12588 10192 12597
rect 10232 12588 10284 12640
rect 12992 12588 13044 12640
rect 13452 12588 13504 12640
rect 14188 12588 14240 12640
rect 16580 12656 16632 12708
rect 17500 12656 17552 12708
rect 17776 12724 17828 12776
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 18236 12724 18288 12776
rect 18696 12767 18748 12776
rect 18696 12733 18705 12767
rect 18705 12733 18739 12767
rect 18739 12733 18748 12767
rect 18696 12724 18748 12733
rect 18788 12724 18840 12776
rect 20996 12792 21048 12844
rect 21272 12835 21324 12844
rect 21272 12801 21281 12835
rect 21281 12801 21315 12835
rect 21315 12801 21324 12835
rect 21272 12792 21324 12801
rect 21456 12835 21508 12844
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 21456 12792 21508 12801
rect 22468 12792 22520 12844
rect 25136 12792 25188 12844
rect 25228 12792 25280 12844
rect 19800 12724 19852 12776
rect 19984 12724 20036 12776
rect 21180 12767 21232 12776
rect 21180 12733 21189 12767
rect 21189 12733 21223 12767
rect 21223 12733 21232 12767
rect 21180 12724 21232 12733
rect 21548 12767 21600 12776
rect 21548 12733 21557 12767
rect 21557 12733 21591 12767
rect 21591 12733 21600 12767
rect 21548 12724 21600 12733
rect 18144 12656 18196 12708
rect 16948 12588 17000 12640
rect 18972 12588 19024 12640
rect 19432 12699 19484 12708
rect 19432 12665 19466 12699
rect 19466 12665 19484 12699
rect 19432 12656 19484 12665
rect 23756 12724 23808 12776
rect 25412 12767 25464 12776
rect 25412 12733 25421 12767
rect 25421 12733 25455 12767
rect 25455 12733 25464 12767
rect 25412 12724 25464 12733
rect 25780 12767 25832 12776
rect 25780 12733 25814 12767
rect 25814 12733 25832 12767
rect 25780 12724 25832 12733
rect 23296 12656 23348 12708
rect 24400 12656 24452 12708
rect 25596 12656 25648 12708
rect 23664 12588 23716 12640
rect 25044 12631 25096 12640
rect 25044 12597 25053 12631
rect 25053 12597 25087 12631
rect 25087 12597 25096 12631
rect 25044 12588 25096 12597
rect 25320 12588 25372 12640
rect 25872 12588 25924 12640
rect 26884 12631 26936 12640
rect 26884 12597 26893 12631
rect 26893 12597 26927 12631
rect 26927 12597 26936 12631
rect 26884 12588 26936 12597
rect 7114 12486 7166 12538
rect 7178 12486 7230 12538
rect 7242 12486 7294 12538
rect 7306 12486 7358 12538
rect 7370 12486 7422 12538
rect 13830 12486 13882 12538
rect 13894 12486 13946 12538
rect 13958 12486 14010 12538
rect 14022 12486 14074 12538
rect 14086 12486 14138 12538
rect 20546 12486 20598 12538
rect 20610 12486 20662 12538
rect 20674 12486 20726 12538
rect 20738 12486 20790 12538
rect 20802 12486 20854 12538
rect 27262 12486 27314 12538
rect 27326 12486 27378 12538
rect 27390 12486 27442 12538
rect 27454 12486 27506 12538
rect 27518 12486 27570 12538
rect 5356 12427 5408 12436
rect 5356 12393 5365 12427
rect 5365 12393 5399 12427
rect 5399 12393 5408 12427
rect 5356 12384 5408 12393
rect 5816 12427 5868 12436
rect 5816 12393 5825 12427
rect 5825 12393 5859 12427
rect 5859 12393 5868 12427
rect 5816 12384 5868 12393
rect 2780 12291 2832 12300
rect 2780 12257 2814 12291
rect 2814 12257 2832 12291
rect 5724 12316 5776 12368
rect 2780 12248 2832 12257
rect 4252 12291 4304 12300
rect 4252 12257 4286 12291
rect 4286 12257 4304 12291
rect 4252 12248 4304 12257
rect 6092 12291 6144 12300
rect 6092 12257 6101 12291
rect 6101 12257 6135 12291
rect 6135 12257 6144 12291
rect 6092 12248 6144 12257
rect 7932 12316 7984 12368
rect 6460 12291 6512 12300
rect 6460 12257 6469 12291
rect 6469 12257 6503 12291
rect 6503 12257 6512 12291
rect 6460 12248 6512 12257
rect 7840 12291 7892 12300
rect 7840 12257 7849 12291
rect 7849 12257 7883 12291
rect 7883 12257 7892 12291
rect 7840 12248 7892 12257
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 8484 12248 8536 12300
rect 10968 12384 11020 12436
rect 8944 12316 8996 12368
rect 9680 12316 9732 12368
rect 14556 12384 14608 12436
rect 14924 12384 14976 12436
rect 15108 12384 15160 12436
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 6736 12180 6788 12232
rect 8300 12223 8352 12232
rect 8300 12189 8309 12223
rect 8309 12189 8343 12223
rect 8343 12189 8352 12223
rect 8300 12180 8352 12189
rect 7380 12112 7432 12164
rect 8208 12112 8260 12164
rect 4712 12044 4764 12096
rect 5172 12044 5224 12096
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 10876 12248 10928 12300
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 9956 12112 10008 12164
rect 11336 12248 11388 12300
rect 14188 12316 14240 12368
rect 14648 12316 14700 12368
rect 12532 12180 12584 12232
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 11980 12112 12032 12164
rect 12440 12112 12492 12164
rect 14280 12248 14332 12300
rect 15016 12316 15068 12368
rect 14832 12291 14884 12300
rect 14832 12257 14841 12291
rect 14841 12257 14875 12291
rect 14875 12257 14884 12291
rect 14832 12248 14884 12257
rect 14924 12291 14976 12300
rect 14924 12257 14933 12291
rect 14933 12257 14967 12291
rect 14967 12257 14976 12291
rect 14924 12248 14976 12257
rect 15200 12248 15252 12300
rect 18144 12384 18196 12436
rect 18328 12384 18380 12436
rect 18420 12427 18472 12436
rect 18420 12393 18429 12427
rect 18429 12393 18463 12427
rect 18463 12393 18472 12427
rect 18420 12384 18472 12393
rect 19432 12384 19484 12436
rect 20352 12384 20404 12436
rect 22744 12384 22796 12436
rect 23020 12384 23072 12436
rect 24952 12384 25004 12436
rect 25320 12384 25372 12436
rect 16856 12316 16908 12368
rect 17040 12248 17092 12300
rect 17592 12316 17644 12368
rect 17776 12316 17828 12368
rect 17868 12316 17920 12368
rect 17684 12291 17736 12300
rect 17684 12257 17693 12291
rect 17693 12257 17727 12291
rect 17727 12257 17736 12291
rect 17684 12248 17736 12257
rect 18512 12248 18564 12300
rect 18972 12291 19024 12300
rect 18972 12257 18981 12291
rect 18981 12257 19015 12291
rect 19015 12257 19024 12291
rect 18972 12248 19024 12257
rect 19616 12291 19668 12300
rect 19616 12257 19625 12291
rect 19625 12257 19659 12291
rect 19659 12257 19668 12291
rect 19616 12248 19668 12257
rect 21548 12316 21600 12368
rect 23664 12316 23716 12368
rect 25044 12316 25096 12368
rect 20352 12248 20404 12300
rect 20444 12248 20496 12300
rect 23756 12248 23808 12300
rect 24492 12248 24544 12300
rect 25136 12291 25188 12300
rect 25136 12257 25145 12291
rect 25145 12257 25179 12291
rect 25179 12257 25188 12291
rect 25136 12248 25188 12257
rect 15016 12112 15068 12164
rect 10140 12044 10192 12096
rect 13084 12087 13136 12096
rect 13084 12053 13093 12087
rect 13093 12053 13127 12087
rect 13127 12053 13136 12087
rect 13084 12044 13136 12053
rect 13268 12044 13320 12096
rect 16396 12087 16448 12096
rect 16396 12053 16405 12087
rect 16405 12053 16439 12087
rect 16439 12053 16448 12087
rect 16396 12044 16448 12053
rect 16580 12112 16632 12164
rect 20996 12180 21048 12232
rect 21640 12180 21692 12232
rect 23296 12180 23348 12232
rect 23480 12180 23532 12232
rect 17592 12112 17644 12164
rect 17684 12112 17736 12164
rect 20076 12044 20128 12096
rect 20260 12044 20312 12096
rect 23112 12044 23164 12096
rect 23572 12087 23624 12096
rect 23572 12053 23581 12087
rect 23581 12053 23615 12087
rect 23615 12053 23624 12087
rect 23572 12044 23624 12053
rect 23664 12044 23716 12096
rect 26884 12180 26936 12232
rect 25228 12044 25280 12096
rect 25412 12044 25464 12096
rect 3756 11942 3808 11994
rect 3820 11942 3872 11994
rect 3884 11942 3936 11994
rect 3948 11942 4000 11994
rect 4012 11942 4064 11994
rect 10472 11942 10524 11994
rect 10536 11942 10588 11994
rect 10600 11942 10652 11994
rect 10664 11942 10716 11994
rect 10728 11942 10780 11994
rect 17188 11942 17240 11994
rect 17252 11942 17304 11994
rect 17316 11942 17368 11994
rect 17380 11942 17432 11994
rect 17444 11942 17496 11994
rect 23904 11942 23956 11994
rect 23968 11942 24020 11994
rect 24032 11942 24084 11994
rect 24096 11942 24148 11994
rect 24160 11942 24212 11994
rect 4252 11840 4304 11892
rect 6276 11840 6328 11892
rect 8024 11840 8076 11892
rect 8300 11840 8352 11892
rect 10324 11840 10376 11892
rect 11428 11840 11480 11892
rect 11980 11883 12032 11892
rect 11980 11849 11989 11883
rect 11989 11849 12023 11883
rect 12023 11849 12032 11883
rect 11980 11840 12032 11849
rect 6368 11772 6420 11824
rect 7932 11772 7984 11824
rect 11888 11704 11940 11756
rect 3240 11636 3292 11688
rect 4988 11679 5040 11688
rect 4988 11645 4997 11679
rect 4997 11645 5031 11679
rect 5031 11645 5040 11679
rect 4988 11636 5040 11645
rect 5356 11679 5408 11688
rect 5356 11645 5365 11679
rect 5365 11645 5399 11679
rect 5399 11645 5408 11679
rect 5356 11636 5408 11645
rect 5540 11679 5592 11688
rect 5540 11645 5549 11679
rect 5549 11645 5583 11679
rect 5583 11645 5592 11679
rect 5540 11636 5592 11645
rect 6276 11679 6328 11688
rect 6276 11645 6285 11679
rect 6285 11645 6319 11679
rect 6319 11645 6328 11679
rect 6276 11636 6328 11645
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 6736 11679 6788 11688
rect 6736 11645 6745 11679
rect 6745 11645 6779 11679
rect 6779 11645 6788 11679
rect 6736 11636 6788 11645
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 7472 11679 7524 11688
rect 7472 11645 7481 11679
rect 7481 11645 7515 11679
rect 7515 11645 7524 11679
rect 7472 11636 7524 11645
rect 7564 11679 7616 11688
rect 7564 11645 7573 11679
rect 7573 11645 7607 11679
rect 7607 11645 7616 11679
rect 7564 11636 7616 11645
rect 4620 11543 4672 11552
rect 4620 11509 4629 11543
rect 4629 11509 4663 11543
rect 4663 11509 4672 11543
rect 4620 11500 4672 11509
rect 5724 11543 5776 11552
rect 5724 11509 5733 11543
rect 5733 11509 5767 11543
rect 5767 11509 5776 11543
rect 5724 11500 5776 11509
rect 6368 11568 6420 11620
rect 7748 11636 7800 11688
rect 8116 11636 8168 11688
rect 9680 11636 9732 11688
rect 8208 11568 8260 11620
rect 9864 11636 9916 11688
rect 10324 11679 10376 11688
rect 10324 11645 10333 11679
rect 10333 11645 10367 11679
rect 10367 11645 10376 11679
rect 10324 11636 10376 11645
rect 11060 11636 11112 11688
rect 11336 11679 11388 11688
rect 11336 11645 11345 11679
rect 11345 11645 11379 11679
rect 11379 11645 11388 11679
rect 11336 11636 11388 11645
rect 11612 11636 11664 11688
rect 7012 11500 7064 11552
rect 8024 11500 8076 11552
rect 11428 11568 11480 11620
rect 13360 11679 13412 11688
rect 13360 11645 13369 11679
rect 13369 11645 13403 11679
rect 13403 11645 13412 11679
rect 13360 11636 13412 11645
rect 14280 11636 14332 11688
rect 14556 11679 14608 11688
rect 14556 11645 14565 11679
rect 14565 11645 14599 11679
rect 14599 11645 14608 11679
rect 14556 11636 14608 11645
rect 14648 11636 14700 11688
rect 19156 11772 19208 11824
rect 20076 11840 20128 11892
rect 20352 11772 20404 11824
rect 21272 11883 21324 11892
rect 21272 11849 21281 11883
rect 21281 11849 21315 11883
rect 21315 11849 21324 11883
rect 21272 11840 21324 11849
rect 23480 11840 23532 11892
rect 23756 11840 23808 11892
rect 27068 11840 27120 11892
rect 21640 11772 21692 11824
rect 17684 11747 17736 11756
rect 17684 11713 17693 11747
rect 17693 11713 17727 11747
rect 17727 11713 17736 11747
rect 17684 11704 17736 11713
rect 18788 11704 18840 11756
rect 13452 11568 13504 11620
rect 14832 11568 14884 11620
rect 8392 11500 8444 11552
rect 9128 11500 9180 11552
rect 9496 11500 9548 11552
rect 11152 11500 11204 11552
rect 14188 11500 14240 11552
rect 18144 11636 18196 11688
rect 23020 11704 23072 11756
rect 22652 11679 22704 11688
rect 22652 11645 22661 11679
rect 22661 11645 22695 11679
rect 22695 11645 22704 11679
rect 22652 11636 22704 11645
rect 24216 11704 24268 11756
rect 24400 11704 24452 11756
rect 23296 11636 23348 11688
rect 18696 11611 18748 11620
rect 18696 11577 18705 11611
rect 18705 11577 18739 11611
rect 18739 11577 18748 11611
rect 18696 11568 18748 11577
rect 18788 11568 18840 11620
rect 15476 11543 15528 11552
rect 15476 11509 15485 11543
rect 15485 11509 15519 11543
rect 15519 11509 15528 11543
rect 15476 11500 15528 11509
rect 16672 11543 16724 11552
rect 16672 11509 16681 11543
rect 16681 11509 16715 11543
rect 16715 11509 16724 11543
rect 16672 11500 16724 11509
rect 16948 11500 17000 11552
rect 17684 11500 17736 11552
rect 18236 11543 18288 11552
rect 18236 11509 18245 11543
rect 18245 11509 18279 11543
rect 18279 11509 18288 11543
rect 18236 11500 18288 11509
rect 19984 11543 20036 11552
rect 19984 11509 19993 11543
rect 19993 11509 20027 11543
rect 20027 11509 20036 11543
rect 19984 11500 20036 11509
rect 22192 11568 22244 11620
rect 23112 11611 23164 11620
rect 23112 11577 23121 11611
rect 23121 11577 23155 11611
rect 23155 11577 23164 11611
rect 23112 11568 23164 11577
rect 25044 11636 25096 11688
rect 22744 11543 22796 11552
rect 22744 11509 22753 11543
rect 22753 11509 22787 11543
rect 22787 11509 22796 11543
rect 22744 11500 22796 11509
rect 24308 11500 24360 11552
rect 25320 11568 25372 11620
rect 26148 11500 26200 11552
rect 7114 11398 7166 11450
rect 7178 11398 7230 11450
rect 7242 11398 7294 11450
rect 7306 11398 7358 11450
rect 7370 11398 7422 11450
rect 13830 11398 13882 11450
rect 13894 11398 13946 11450
rect 13958 11398 14010 11450
rect 14022 11398 14074 11450
rect 14086 11398 14138 11450
rect 20546 11398 20598 11450
rect 20610 11398 20662 11450
rect 20674 11398 20726 11450
rect 20738 11398 20790 11450
rect 20802 11398 20854 11450
rect 27262 11398 27314 11450
rect 27326 11398 27378 11450
rect 27390 11398 27442 11450
rect 27454 11398 27506 11450
rect 27518 11398 27570 11450
rect 1400 11296 1452 11348
rect 3148 11203 3200 11212
rect 3148 11169 3157 11203
rect 3157 11169 3191 11203
rect 3191 11169 3200 11203
rect 3148 11160 3200 11169
rect 4252 11160 4304 11212
rect 4344 11092 4396 11144
rect 7564 11296 7616 11348
rect 8116 11339 8168 11348
rect 8116 11305 8125 11339
rect 8125 11305 8159 11339
rect 8159 11305 8168 11339
rect 8116 11296 8168 11305
rect 8208 11339 8260 11348
rect 8208 11305 8217 11339
rect 8217 11305 8251 11339
rect 8251 11305 8260 11339
rect 8208 11296 8260 11305
rect 4988 11160 5040 11212
rect 5172 11160 5224 11212
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 6828 11160 6880 11212
rect 7012 11271 7064 11280
rect 7012 11237 7046 11271
rect 7046 11237 7064 11271
rect 7012 11228 7064 11237
rect 8392 11271 8444 11280
rect 8392 11237 8401 11271
rect 8401 11237 8435 11271
rect 8435 11237 8444 11271
rect 8392 11228 8444 11237
rect 9404 11296 9456 11348
rect 12348 11296 12400 11348
rect 13544 11296 13596 11348
rect 13820 11296 13872 11348
rect 21456 11296 21508 11348
rect 23296 11296 23348 11348
rect 24492 11339 24544 11348
rect 24492 11305 24501 11339
rect 24501 11305 24535 11339
rect 24535 11305 24544 11339
rect 24492 11296 24544 11305
rect 25320 11339 25372 11348
rect 25320 11305 25329 11339
rect 25329 11305 25363 11339
rect 25363 11305 25372 11339
rect 25320 11296 25372 11305
rect 9128 11228 9180 11280
rect 11888 11228 11940 11280
rect 16580 11228 16632 11280
rect 19248 11271 19300 11280
rect 19248 11237 19257 11271
rect 19257 11237 19291 11271
rect 19291 11237 19300 11271
rect 19248 11228 19300 11237
rect 21548 11271 21600 11280
rect 21548 11237 21557 11271
rect 21557 11237 21591 11271
rect 21591 11237 21600 11271
rect 21548 11228 21600 11237
rect 23480 11271 23532 11280
rect 23480 11237 23489 11271
rect 23489 11237 23523 11271
rect 23523 11237 23532 11271
rect 23480 11228 23532 11237
rect 24216 11228 24268 11280
rect 24860 11228 24912 11280
rect 7472 11160 7524 11212
rect 5540 11092 5592 11144
rect 10048 11160 10100 11212
rect 11060 11160 11112 11212
rect 11244 11203 11296 11212
rect 11244 11169 11254 11203
rect 11254 11169 11288 11203
rect 11288 11169 11296 11203
rect 11244 11160 11296 11169
rect 11428 11203 11480 11212
rect 11428 11169 11437 11203
rect 11437 11169 11471 11203
rect 11471 11169 11480 11203
rect 11428 11160 11480 11169
rect 11704 11160 11756 11212
rect 12624 11203 12676 11212
rect 12624 11169 12658 11203
rect 12658 11169 12676 11203
rect 12624 11160 12676 11169
rect 16304 11160 16356 11212
rect 16488 11203 16540 11212
rect 16488 11169 16522 11203
rect 16522 11169 16540 11203
rect 16488 11160 16540 11169
rect 17592 11160 17644 11212
rect 18512 11203 18564 11212
rect 18512 11169 18521 11203
rect 18521 11169 18555 11203
rect 18555 11169 18564 11203
rect 18512 11160 18564 11169
rect 18880 11203 18932 11212
rect 18880 11169 18889 11203
rect 18889 11169 18923 11203
rect 18923 11169 18932 11203
rect 18880 11160 18932 11169
rect 19524 11203 19576 11212
rect 19524 11169 19533 11203
rect 19533 11169 19567 11203
rect 19567 11169 19576 11203
rect 19524 11160 19576 11169
rect 19616 11203 19668 11212
rect 19616 11169 19625 11203
rect 19625 11169 19659 11203
rect 19659 11169 19668 11203
rect 19616 11160 19668 11169
rect 19708 11203 19760 11212
rect 19708 11169 19717 11203
rect 19717 11169 19751 11203
rect 19751 11169 19760 11203
rect 19708 11160 19760 11169
rect 19892 11203 19944 11212
rect 19892 11169 19901 11203
rect 19901 11169 19935 11203
rect 19935 11169 19944 11203
rect 19892 11160 19944 11169
rect 22652 11160 22704 11212
rect 25044 11160 25096 11212
rect 25136 11160 25188 11212
rect 25688 11160 25740 11212
rect 5080 11024 5132 11076
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 10968 11092 11020 11144
rect 9404 11024 9456 11076
rect 9680 11024 9732 11076
rect 3332 10999 3384 11008
rect 3332 10965 3341 10999
rect 3341 10965 3375 10999
rect 3375 10965 3384 10999
rect 3332 10956 3384 10965
rect 8392 10956 8444 11008
rect 12164 10956 12216 11008
rect 18604 11135 18656 11144
rect 18604 11101 18613 11135
rect 18613 11101 18647 11135
rect 18647 11101 18656 11135
rect 18604 11092 18656 11101
rect 20536 11092 20588 11144
rect 23572 11092 23624 11144
rect 24124 11135 24176 11144
rect 24124 11101 24133 11135
rect 24133 11101 24167 11135
rect 24167 11101 24176 11135
rect 24124 11092 24176 11101
rect 24216 11135 24268 11144
rect 24216 11101 24225 11135
rect 24225 11101 24259 11135
rect 24259 11101 24268 11135
rect 24216 11092 24268 11101
rect 24308 11135 24360 11144
rect 24308 11101 24317 11135
rect 24317 11101 24351 11135
rect 24351 11101 24360 11135
rect 24308 11092 24360 11101
rect 17960 11024 18012 11076
rect 20076 11024 20128 11076
rect 25596 11092 25648 11144
rect 26148 11203 26200 11212
rect 26148 11169 26157 11203
rect 26157 11169 26191 11203
rect 26191 11169 26200 11203
rect 26148 11160 26200 11169
rect 13360 10956 13412 11008
rect 14280 10956 14332 11008
rect 16948 10956 17000 11008
rect 22560 10956 22612 11008
rect 23572 10956 23624 11008
rect 24216 10956 24268 11008
rect 25780 10956 25832 11008
rect 25872 10956 25924 11008
rect 26056 10999 26108 11008
rect 26056 10965 26065 10999
rect 26065 10965 26099 10999
rect 26099 10965 26108 10999
rect 26056 10956 26108 10965
rect 3756 10854 3808 10906
rect 3820 10854 3872 10906
rect 3884 10854 3936 10906
rect 3948 10854 4000 10906
rect 4012 10854 4064 10906
rect 10472 10854 10524 10906
rect 10536 10854 10588 10906
rect 10600 10854 10652 10906
rect 10664 10854 10716 10906
rect 10728 10854 10780 10906
rect 17188 10854 17240 10906
rect 17252 10854 17304 10906
rect 17316 10854 17368 10906
rect 17380 10854 17432 10906
rect 17444 10854 17496 10906
rect 23904 10854 23956 10906
rect 23968 10854 24020 10906
rect 24032 10854 24084 10906
rect 24096 10854 24148 10906
rect 24160 10854 24212 10906
rect 4896 10684 4948 10736
rect 2504 10548 2556 10600
rect 3332 10548 3384 10600
rect 6000 10548 6052 10600
rect 6368 10548 6420 10600
rect 7748 10752 7800 10804
rect 9864 10752 9916 10804
rect 11244 10752 11296 10804
rect 7932 10727 7984 10736
rect 7932 10693 7941 10727
rect 7941 10693 7975 10727
rect 7975 10693 7984 10727
rect 7932 10684 7984 10693
rect 8392 10684 8444 10736
rect 10140 10616 10192 10668
rect 12348 10684 12400 10736
rect 12624 10795 12676 10804
rect 12624 10761 12633 10795
rect 12633 10761 12667 10795
rect 12667 10761 12676 10795
rect 12624 10752 12676 10761
rect 15568 10795 15620 10804
rect 15568 10761 15577 10795
rect 15577 10761 15611 10795
rect 15611 10761 15620 10795
rect 15568 10752 15620 10761
rect 16488 10752 16540 10804
rect 18880 10752 18932 10804
rect 19708 10752 19760 10804
rect 21272 10795 21324 10804
rect 21272 10761 21281 10795
rect 21281 10761 21315 10795
rect 21315 10761 21324 10795
rect 21272 10752 21324 10761
rect 22100 10795 22152 10804
rect 22100 10761 22109 10795
rect 22109 10761 22143 10795
rect 22143 10761 22152 10795
rect 22100 10752 22152 10761
rect 22192 10795 22244 10804
rect 22192 10761 22201 10795
rect 22201 10761 22235 10795
rect 22235 10761 22244 10795
rect 22192 10752 22244 10761
rect 23756 10752 23808 10804
rect 2412 10480 2464 10532
rect 7840 10591 7892 10600
rect 7840 10557 7849 10591
rect 7849 10557 7883 10591
rect 7883 10557 7892 10591
rect 7840 10548 7892 10557
rect 8116 10548 8168 10600
rect 8300 10548 8352 10600
rect 8944 10548 8996 10600
rect 11060 10548 11112 10600
rect 11704 10591 11756 10600
rect 11704 10557 11718 10591
rect 11718 10557 11752 10591
rect 11752 10557 11756 10591
rect 11704 10548 11756 10557
rect 11980 10591 12032 10600
rect 11980 10557 11989 10591
rect 11989 10557 12023 10591
rect 12023 10557 12032 10591
rect 11980 10548 12032 10557
rect 12164 10591 12216 10600
rect 12164 10557 12173 10591
rect 12173 10557 12207 10591
rect 12207 10557 12216 10591
rect 12164 10548 12216 10557
rect 12256 10591 12308 10600
rect 12256 10557 12265 10591
rect 12265 10557 12299 10591
rect 12299 10557 12308 10591
rect 12256 10548 12308 10557
rect 12716 10591 12768 10600
rect 12716 10557 12725 10591
rect 12725 10557 12759 10591
rect 12759 10557 12768 10591
rect 12716 10548 12768 10557
rect 16580 10727 16632 10736
rect 16580 10693 16589 10727
rect 16589 10693 16623 10727
rect 16623 10693 16632 10727
rect 16580 10684 16632 10693
rect 16672 10684 16724 10736
rect 20076 10684 20128 10736
rect 7932 10480 7984 10532
rect 11520 10523 11572 10532
rect 11520 10489 11529 10523
rect 11529 10489 11563 10523
rect 11563 10489 11572 10523
rect 11520 10480 11572 10489
rect 14280 10548 14332 10600
rect 15660 10548 15712 10600
rect 17960 10659 18012 10668
rect 17960 10625 17969 10659
rect 17969 10625 18003 10659
rect 18003 10625 18012 10659
rect 17960 10616 18012 10625
rect 16672 10591 16724 10600
rect 16672 10557 16681 10591
rect 16681 10557 16715 10591
rect 16715 10557 16724 10591
rect 16672 10548 16724 10557
rect 16764 10591 16816 10600
rect 16764 10557 16773 10591
rect 16773 10557 16807 10591
rect 16807 10557 16816 10591
rect 16764 10548 16816 10557
rect 16948 10591 17000 10600
rect 16948 10557 16957 10591
rect 16957 10557 16991 10591
rect 16991 10557 17000 10591
rect 16948 10548 17000 10557
rect 20076 10591 20128 10600
rect 20076 10557 20085 10591
rect 20085 10557 20119 10591
rect 20119 10557 20128 10591
rect 20076 10548 20128 10557
rect 4160 10412 4212 10464
rect 4712 10455 4764 10464
rect 4712 10421 4721 10455
rect 4721 10421 4755 10455
rect 4755 10421 4764 10455
rect 4712 10412 4764 10421
rect 9128 10412 9180 10464
rect 9680 10412 9732 10464
rect 18144 10480 18196 10532
rect 18328 10480 18380 10532
rect 20352 10591 20404 10600
rect 12440 10412 12492 10464
rect 12900 10412 12952 10464
rect 17224 10412 17276 10464
rect 18052 10412 18104 10464
rect 20352 10557 20361 10591
rect 20361 10557 20395 10591
rect 20395 10557 20404 10591
rect 20352 10548 20404 10557
rect 20536 10591 20588 10600
rect 20536 10557 20545 10591
rect 20545 10557 20579 10591
rect 20579 10557 20588 10591
rect 20536 10548 20588 10557
rect 21088 10591 21140 10600
rect 21088 10557 21097 10591
rect 21097 10557 21131 10591
rect 21131 10557 21140 10591
rect 21088 10548 21140 10557
rect 21456 10659 21508 10668
rect 21456 10625 21465 10659
rect 21465 10625 21499 10659
rect 21499 10625 21508 10659
rect 21456 10616 21508 10625
rect 22560 10659 22612 10668
rect 22560 10625 22569 10659
rect 22569 10625 22603 10659
rect 22603 10625 22612 10659
rect 22560 10616 22612 10625
rect 22928 10727 22980 10736
rect 22928 10693 22937 10727
rect 22937 10693 22971 10727
rect 22971 10693 22980 10727
rect 22928 10684 22980 10693
rect 22376 10591 22428 10600
rect 22376 10557 22385 10591
rect 22385 10557 22419 10591
rect 22419 10557 22428 10591
rect 22376 10548 22428 10557
rect 22744 10548 22796 10600
rect 21456 10480 21508 10532
rect 24124 10727 24176 10736
rect 24124 10693 24133 10727
rect 24133 10693 24167 10727
rect 24167 10693 24176 10727
rect 24124 10684 24176 10693
rect 25780 10727 25832 10736
rect 25780 10693 25789 10727
rect 25789 10693 25823 10727
rect 25823 10693 25832 10727
rect 25780 10684 25832 10693
rect 20904 10455 20956 10464
rect 20904 10421 20913 10455
rect 20913 10421 20947 10455
rect 20947 10421 20956 10455
rect 20904 10412 20956 10421
rect 21272 10412 21324 10464
rect 21824 10412 21876 10464
rect 22836 10455 22888 10464
rect 22836 10421 22845 10455
rect 22845 10421 22879 10455
rect 22879 10421 22888 10455
rect 22836 10412 22888 10421
rect 23572 10480 23624 10532
rect 24032 10591 24084 10600
rect 24032 10557 24041 10591
rect 24041 10557 24075 10591
rect 24075 10557 24084 10591
rect 24032 10548 24084 10557
rect 24676 10591 24728 10600
rect 24676 10557 24685 10591
rect 24685 10557 24719 10591
rect 24719 10557 24728 10591
rect 24676 10548 24728 10557
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 25596 10591 25648 10600
rect 25596 10557 25605 10591
rect 25605 10557 25639 10591
rect 25639 10557 25648 10591
rect 25596 10548 25648 10557
rect 25872 10591 25924 10600
rect 25872 10557 25881 10591
rect 25881 10557 25915 10591
rect 25915 10557 25924 10591
rect 25872 10548 25924 10557
rect 25780 10412 25832 10464
rect 7114 10310 7166 10362
rect 7178 10310 7230 10362
rect 7242 10310 7294 10362
rect 7306 10310 7358 10362
rect 7370 10310 7422 10362
rect 13830 10310 13882 10362
rect 13894 10310 13946 10362
rect 13958 10310 14010 10362
rect 14022 10310 14074 10362
rect 14086 10310 14138 10362
rect 20546 10310 20598 10362
rect 20610 10310 20662 10362
rect 20674 10310 20726 10362
rect 20738 10310 20790 10362
rect 20802 10310 20854 10362
rect 27262 10310 27314 10362
rect 27326 10310 27378 10362
rect 27390 10310 27442 10362
rect 27454 10310 27506 10362
rect 27518 10310 27570 10362
rect 2412 10208 2464 10260
rect 4160 10208 4212 10260
rect 4252 10251 4304 10260
rect 4252 10217 4261 10251
rect 4261 10217 4295 10251
rect 4295 10217 4304 10251
rect 4252 10208 4304 10217
rect 7840 10208 7892 10260
rect 9128 10208 9180 10260
rect 16672 10208 16724 10260
rect 16764 10208 16816 10260
rect 17960 10208 18012 10260
rect 18512 10251 18564 10260
rect 18512 10217 18521 10251
rect 18521 10217 18555 10251
rect 18555 10217 18564 10251
rect 18512 10208 18564 10217
rect 18696 10208 18748 10260
rect 2044 10115 2096 10124
rect 2044 10081 2053 10115
rect 2053 10081 2087 10115
rect 2087 10081 2096 10115
rect 2044 10072 2096 10081
rect 3608 10140 3660 10192
rect 2872 10072 2924 10124
rect 3148 9936 3200 9988
rect 4712 10072 4764 10124
rect 4896 10115 4948 10124
rect 4896 10081 4905 10115
rect 4905 10081 4939 10115
rect 4939 10081 4948 10115
rect 4896 10072 4948 10081
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 5172 10072 5224 10124
rect 5908 10115 5960 10124
rect 5908 10081 5917 10115
rect 5917 10081 5951 10115
rect 5951 10081 5960 10115
rect 5908 10072 5960 10081
rect 6368 10072 6420 10124
rect 6920 10072 6972 10124
rect 8208 10072 8260 10124
rect 10048 10115 10100 10124
rect 10048 10081 10057 10115
rect 10057 10081 10091 10115
rect 10091 10081 10100 10115
rect 10048 10072 10100 10081
rect 11060 10115 11112 10124
rect 11060 10081 11069 10115
rect 11069 10081 11103 10115
rect 11103 10081 11112 10115
rect 11060 10072 11112 10081
rect 11244 10115 11296 10124
rect 11244 10081 11251 10115
rect 11251 10081 11296 10115
rect 11244 10072 11296 10081
rect 11336 10115 11388 10124
rect 11336 10081 11345 10115
rect 11345 10081 11379 10115
rect 11379 10081 11388 10115
rect 11336 10072 11388 10081
rect 4252 10047 4304 10056
rect 4252 10013 4261 10047
rect 4261 10013 4295 10047
rect 4295 10013 4304 10047
rect 4252 10004 4304 10013
rect 4436 10047 4488 10056
rect 4436 10013 4445 10047
rect 4445 10013 4479 10047
rect 4479 10013 4488 10047
rect 4436 10004 4488 10013
rect 11428 10004 11480 10056
rect 2228 9911 2280 9920
rect 2228 9877 2237 9911
rect 2237 9877 2271 9911
rect 2271 9877 2280 9911
rect 2228 9868 2280 9877
rect 4252 9868 4304 9920
rect 5080 9868 5132 9920
rect 8392 9868 8444 9920
rect 11704 10072 11756 10124
rect 11888 10072 11940 10124
rect 12440 10140 12492 10192
rect 14280 10140 14332 10192
rect 17224 10183 17276 10192
rect 17224 10149 17233 10183
rect 17233 10149 17267 10183
rect 17267 10149 17276 10183
rect 17224 10140 17276 10149
rect 17684 10140 17736 10192
rect 19248 10183 19300 10192
rect 19248 10149 19282 10183
rect 19282 10149 19300 10183
rect 19248 10140 19300 10149
rect 19708 10208 19760 10260
rect 22744 10208 22796 10260
rect 23296 10208 23348 10260
rect 24676 10208 24728 10260
rect 26056 10208 26108 10260
rect 20904 10140 20956 10192
rect 11796 9936 11848 9988
rect 14372 10072 14424 10124
rect 18052 10072 18104 10124
rect 19708 10072 19760 10124
rect 22652 10140 22704 10192
rect 23480 10183 23532 10192
rect 23480 10149 23489 10183
rect 23489 10149 23523 10183
rect 23523 10149 23532 10183
rect 23480 10140 23532 10149
rect 24308 10140 24360 10192
rect 21548 10115 21600 10124
rect 21548 10081 21582 10115
rect 21582 10081 21600 10115
rect 21548 10072 21600 10081
rect 23020 10115 23072 10124
rect 23020 10081 23029 10115
rect 23029 10081 23063 10115
rect 23063 10081 23072 10115
rect 23020 10072 23072 10081
rect 25504 10140 25556 10192
rect 18696 10004 18748 10056
rect 12256 9868 12308 9920
rect 14464 9936 14516 9988
rect 22560 10004 22612 10056
rect 22928 10004 22980 10056
rect 25228 10072 25280 10124
rect 25320 10115 25372 10124
rect 25320 10081 25329 10115
rect 25329 10081 25363 10115
rect 25363 10081 25372 10115
rect 25320 10072 25372 10081
rect 20352 9979 20404 9988
rect 20352 9945 20361 9979
rect 20361 9945 20395 9979
rect 20395 9945 20404 9979
rect 20352 9936 20404 9945
rect 19340 9868 19392 9920
rect 20076 9868 20128 9920
rect 21088 9868 21140 9920
rect 23664 9936 23716 9988
rect 22560 9868 22612 9920
rect 22744 9868 22796 9920
rect 22928 9868 22980 9920
rect 24032 9868 24084 9920
rect 24768 9911 24820 9920
rect 24768 9877 24777 9911
rect 24777 9877 24811 9911
rect 24811 9877 24820 9911
rect 24768 9868 24820 9877
rect 24860 9911 24912 9920
rect 24860 9877 24869 9911
rect 24869 9877 24903 9911
rect 24903 9877 24912 9911
rect 24860 9868 24912 9877
rect 3756 9766 3808 9818
rect 3820 9766 3872 9818
rect 3884 9766 3936 9818
rect 3948 9766 4000 9818
rect 4012 9766 4064 9818
rect 10472 9766 10524 9818
rect 10536 9766 10588 9818
rect 10600 9766 10652 9818
rect 10664 9766 10716 9818
rect 10728 9766 10780 9818
rect 17188 9766 17240 9818
rect 17252 9766 17304 9818
rect 17316 9766 17368 9818
rect 17380 9766 17432 9818
rect 17444 9766 17496 9818
rect 23904 9766 23956 9818
rect 23968 9766 24020 9818
rect 24032 9766 24084 9818
rect 24096 9766 24148 9818
rect 24160 9766 24212 9818
rect 2044 9664 2096 9716
rect 2872 9664 2924 9716
rect 4160 9664 4212 9716
rect 4804 9664 4856 9716
rect 8208 9707 8260 9716
rect 8208 9673 8217 9707
rect 8217 9673 8251 9707
rect 8251 9673 8260 9707
rect 8208 9664 8260 9673
rect 2136 9596 2188 9648
rect 3608 9596 3660 9648
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 2228 9528 2280 9580
rect 5080 9596 5132 9648
rect 7748 9596 7800 9648
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 2136 9392 2188 9444
rect 3056 9435 3108 9444
rect 3056 9401 3065 9435
rect 3065 9401 3099 9435
rect 3099 9401 3108 9435
rect 3056 9392 3108 9401
rect 2596 9324 2648 9376
rect 3792 9503 3844 9512
rect 3792 9469 3801 9503
rect 3801 9469 3835 9503
rect 3835 9469 3844 9503
rect 3792 9460 3844 9469
rect 4252 9503 4304 9512
rect 4252 9469 4261 9503
rect 4261 9469 4295 9503
rect 4295 9469 4304 9503
rect 4252 9460 4304 9469
rect 4436 9503 4488 9512
rect 4436 9469 4445 9503
rect 4445 9469 4479 9503
rect 4479 9469 4488 9503
rect 4436 9460 4488 9469
rect 5908 9528 5960 9580
rect 8116 9596 8168 9648
rect 8576 9596 8628 9648
rect 9772 9596 9824 9648
rect 12716 9596 12768 9648
rect 13544 9596 13596 9648
rect 15200 9596 15252 9648
rect 16580 9664 16632 9716
rect 16856 9664 16908 9716
rect 21548 9664 21600 9716
rect 22192 9664 22244 9716
rect 22560 9664 22612 9716
rect 23020 9664 23072 9716
rect 19248 9596 19300 9648
rect 19616 9596 19668 9648
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 5172 9503 5224 9512
rect 5172 9469 5181 9503
rect 5181 9469 5215 9503
rect 5215 9469 5224 9503
rect 5172 9460 5224 9469
rect 5632 9460 5684 9512
rect 6368 9503 6420 9512
rect 6368 9469 6377 9503
rect 6377 9469 6411 9503
rect 6411 9469 6420 9503
rect 6368 9460 6420 9469
rect 6920 9460 6972 9512
rect 8024 9528 8076 9580
rect 5908 9435 5960 9444
rect 5908 9401 5917 9435
rect 5917 9401 5951 9435
rect 5951 9401 5960 9435
rect 5908 9392 5960 9401
rect 8392 9460 8444 9512
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 9220 9460 9272 9512
rect 13452 9528 13504 9580
rect 14004 9571 14056 9580
rect 14004 9537 14013 9571
rect 14013 9537 14047 9571
rect 14047 9537 14056 9571
rect 14004 9528 14056 9537
rect 9588 9460 9640 9512
rect 11428 9460 11480 9512
rect 11704 9503 11756 9512
rect 11704 9469 11711 9503
rect 11711 9469 11756 9503
rect 11704 9460 11756 9469
rect 12256 9460 12308 9512
rect 12348 9503 12400 9512
rect 12348 9469 12357 9503
rect 12357 9469 12391 9503
rect 12391 9469 12400 9503
rect 12348 9460 12400 9469
rect 13360 9460 13412 9512
rect 4252 9324 4304 9376
rect 4988 9324 5040 9376
rect 5080 9324 5132 9376
rect 5816 9367 5868 9376
rect 5816 9333 5825 9367
rect 5825 9333 5859 9367
rect 5859 9333 5868 9367
rect 5816 9324 5868 9333
rect 8484 9324 8536 9376
rect 9128 9367 9180 9376
rect 9128 9333 9137 9367
rect 9137 9333 9171 9367
rect 9171 9333 9180 9367
rect 9128 9324 9180 9333
rect 10048 9392 10100 9444
rect 11336 9392 11388 9444
rect 11796 9435 11848 9444
rect 11796 9401 11805 9435
rect 11805 9401 11839 9435
rect 11839 9401 11848 9435
rect 11796 9392 11848 9401
rect 9680 9324 9732 9376
rect 9864 9324 9916 9376
rect 15660 9392 15712 9444
rect 15752 9435 15804 9444
rect 15752 9401 15761 9435
rect 15761 9401 15795 9435
rect 15795 9401 15804 9435
rect 15752 9392 15804 9401
rect 18328 9528 18380 9580
rect 22836 9596 22888 9648
rect 16488 9460 16540 9512
rect 18788 9460 18840 9512
rect 16764 9392 16816 9444
rect 16856 9392 16908 9444
rect 11980 9324 12032 9376
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 12808 9324 12860 9376
rect 16120 9324 16172 9376
rect 17868 9324 17920 9376
rect 19248 9324 19300 9376
rect 19524 9324 19576 9376
rect 19708 9435 19760 9444
rect 19708 9401 19717 9435
rect 19717 9401 19751 9435
rect 19751 9401 19760 9435
rect 19708 9392 19760 9401
rect 19892 9503 19944 9512
rect 19892 9469 19900 9503
rect 19900 9469 19934 9503
rect 19934 9469 19944 9503
rect 19892 9460 19944 9469
rect 20904 9460 20956 9512
rect 21180 9460 21232 9512
rect 21456 9460 21508 9512
rect 22192 9503 22244 9512
rect 22192 9469 22201 9503
rect 22201 9469 22235 9503
rect 22235 9469 22244 9503
rect 22192 9460 22244 9469
rect 20168 9392 20220 9444
rect 22468 9503 22520 9512
rect 22468 9469 22477 9503
rect 22477 9469 22511 9503
rect 22511 9469 22520 9503
rect 22468 9460 22520 9469
rect 24032 9503 24084 9512
rect 24032 9469 24049 9503
rect 24049 9469 24084 9503
rect 24032 9460 24084 9469
rect 24400 9528 24452 9580
rect 24216 9435 24268 9444
rect 24216 9401 24225 9435
rect 24225 9401 24259 9435
rect 24259 9401 24268 9435
rect 24216 9392 24268 9401
rect 24492 9503 24544 9512
rect 24492 9469 24501 9503
rect 24501 9469 24535 9503
rect 24535 9469 24544 9503
rect 24492 9460 24544 9469
rect 24952 9528 25004 9580
rect 25780 9664 25832 9716
rect 24860 9460 24912 9512
rect 25320 9503 25372 9512
rect 25320 9469 25329 9503
rect 25329 9469 25363 9503
rect 25363 9469 25372 9503
rect 25320 9460 25372 9469
rect 26792 9528 26844 9580
rect 25780 9503 25832 9512
rect 25780 9469 25789 9503
rect 25789 9469 25823 9503
rect 25823 9469 25832 9503
rect 25780 9460 25832 9469
rect 21088 9324 21140 9376
rect 24032 9324 24084 9376
rect 25320 9324 25372 9376
rect 25412 9324 25464 9376
rect 7114 9222 7166 9274
rect 7178 9222 7230 9274
rect 7242 9222 7294 9274
rect 7306 9222 7358 9274
rect 7370 9222 7422 9274
rect 13830 9222 13882 9274
rect 13894 9222 13946 9274
rect 13958 9222 14010 9274
rect 14022 9222 14074 9274
rect 14086 9222 14138 9274
rect 20546 9222 20598 9274
rect 20610 9222 20662 9274
rect 20674 9222 20726 9274
rect 20738 9222 20790 9274
rect 20802 9222 20854 9274
rect 27262 9222 27314 9274
rect 27326 9222 27378 9274
rect 27390 9222 27442 9274
rect 27454 9222 27506 9274
rect 27518 9222 27570 9274
rect 3792 9120 3844 9172
rect 5632 9163 5684 9172
rect 5632 9129 5641 9163
rect 5641 9129 5675 9163
rect 5675 9129 5684 9163
rect 5632 9120 5684 9129
rect 8760 9120 8812 9172
rect 9588 9163 9640 9172
rect 9588 9129 9597 9163
rect 9597 9129 9631 9163
rect 9631 9129 9640 9163
rect 9588 9120 9640 9129
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 1952 9052 2004 9104
rect 3056 9052 3108 9104
rect 4436 9052 4488 9104
rect 5172 9052 5224 9104
rect 5816 9052 5868 9104
rect 5264 8984 5316 9036
rect 6368 9027 6420 9036
rect 6368 8993 6377 9027
rect 6377 8993 6411 9027
rect 6411 8993 6420 9027
rect 6368 8984 6420 8993
rect 6920 8984 6972 9036
rect 9128 9052 9180 9104
rect 9220 9052 9272 9104
rect 11980 9120 12032 9172
rect 12348 9163 12400 9172
rect 12348 9129 12357 9163
rect 12357 9129 12391 9163
rect 12391 9129 12400 9163
rect 12348 9120 12400 9129
rect 12992 9120 13044 9172
rect 13452 9163 13504 9172
rect 13452 9129 13461 9163
rect 13461 9129 13495 9163
rect 13495 9129 13504 9163
rect 13452 9120 13504 9129
rect 9864 9095 9916 9104
rect 9864 9061 9873 9095
rect 9873 9061 9907 9095
rect 9907 9061 9916 9095
rect 9864 9052 9916 9061
rect 10048 9095 10100 9104
rect 10048 9061 10057 9095
rect 10057 9061 10091 9095
rect 10091 9061 10100 9095
rect 10048 9052 10100 9061
rect 1492 8959 1544 8968
rect 1492 8925 1501 8959
rect 1501 8925 1535 8959
rect 1535 8925 1544 8959
rect 1492 8916 1544 8925
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 6092 8916 6144 8968
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 8116 8984 8168 9036
rect 8300 8984 8352 9036
rect 8484 9027 8536 9036
rect 8484 8993 8518 9027
rect 8518 8993 8536 9027
rect 8484 8984 8536 8993
rect 8024 8916 8076 8968
rect 7012 8848 7064 8900
rect 4436 8780 4488 8832
rect 6276 8780 6328 8832
rect 8116 8823 8168 8832
rect 8116 8789 8125 8823
rect 8125 8789 8159 8823
rect 8159 8789 8168 8823
rect 8116 8780 8168 8789
rect 8208 8780 8260 8832
rect 11244 9027 11296 9036
rect 11244 8993 11278 9027
rect 11278 8993 11296 9027
rect 11244 8984 11296 8993
rect 11520 9052 11572 9104
rect 11888 9052 11940 9104
rect 12164 9052 12216 9104
rect 13176 8984 13228 9036
rect 13544 9027 13596 9036
rect 13544 8993 13553 9027
rect 13553 8993 13587 9027
rect 13587 8993 13596 9027
rect 13544 8984 13596 8993
rect 14004 9052 14056 9104
rect 14740 9052 14792 9104
rect 16856 9163 16908 9172
rect 16856 9129 16865 9163
rect 16865 9129 16899 9163
rect 16899 9129 16908 9163
rect 16856 9120 16908 9129
rect 16764 9052 16816 9104
rect 19064 9120 19116 9172
rect 9680 8916 9732 8968
rect 12164 8916 12216 8968
rect 12900 8916 12952 8968
rect 13268 8916 13320 8968
rect 14280 9027 14332 9036
rect 14280 8993 14289 9027
rect 14289 8993 14323 9027
rect 14323 8993 14332 9027
rect 14280 8984 14332 8993
rect 9312 8848 9364 8900
rect 10140 8848 10192 8900
rect 10508 8848 10560 8900
rect 11980 8848 12032 8900
rect 16120 9027 16172 9036
rect 16120 8993 16129 9027
rect 16129 8993 16163 9027
rect 16163 8993 16172 9027
rect 16120 8984 16172 8993
rect 16304 8984 16356 9036
rect 16856 8984 16908 9036
rect 17132 9027 17184 9036
rect 17132 8993 17141 9027
rect 17141 8993 17175 9027
rect 17175 8993 17184 9027
rect 17132 8984 17184 8993
rect 18420 9052 18472 9104
rect 17684 8984 17736 9036
rect 17868 8984 17920 9036
rect 18328 9027 18380 9036
rect 18328 8993 18337 9027
rect 18337 8993 18371 9027
rect 18371 8993 18380 9027
rect 18328 8984 18380 8993
rect 19156 8984 19208 9036
rect 19248 8984 19300 9036
rect 24492 9120 24544 9172
rect 24584 9120 24636 9172
rect 21548 9052 21600 9104
rect 21824 9052 21876 9104
rect 18052 8916 18104 8968
rect 22468 8984 22520 9036
rect 24952 9052 25004 9104
rect 24308 8916 24360 8968
rect 24860 8984 24912 9036
rect 25136 9027 25188 9036
rect 25136 8993 25145 9027
rect 25145 8993 25179 9027
rect 25179 8993 25188 9027
rect 25136 8984 25188 8993
rect 25320 9027 25372 9036
rect 25320 8993 25329 9027
rect 25329 8993 25363 9027
rect 25363 8993 25372 9027
rect 25320 8984 25372 8993
rect 25412 9027 25464 9036
rect 25412 8993 25421 9027
rect 25421 8993 25455 9027
rect 25455 8993 25464 9027
rect 25412 8984 25464 8993
rect 25596 8984 25648 9036
rect 25780 8984 25832 9036
rect 25964 8984 26016 9036
rect 11612 8780 11664 8832
rect 12532 8780 12584 8832
rect 17960 8848 18012 8900
rect 19524 8848 19576 8900
rect 16948 8780 17000 8832
rect 20628 8823 20680 8832
rect 20628 8789 20637 8823
rect 20637 8789 20671 8823
rect 20671 8789 20680 8823
rect 20628 8780 20680 8789
rect 24492 8848 24544 8900
rect 26792 8916 26844 8968
rect 25964 8848 26016 8900
rect 24032 8780 24084 8832
rect 24676 8823 24728 8832
rect 24676 8789 24685 8823
rect 24685 8789 24719 8823
rect 24719 8789 24728 8823
rect 24676 8780 24728 8789
rect 24768 8823 24820 8832
rect 24768 8789 24777 8823
rect 24777 8789 24811 8823
rect 24811 8789 24820 8823
rect 24768 8780 24820 8789
rect 25780 8823 25832 8832
rect 25780 8789 25789 8823
rect 25789 8789 25823 8823
rect 25823 8789 25832 8823
rect 25780 8780 25832 8789
rect 25872 8823 25924 8832
rect 25872 8789 25881 8823
rect 25881 8789 25915 8823
rect 25915 8789 25924 8823
rect 25872 8780 25924 8789
rect 3756 8678 3808 8730
rect 3820 8678 3872 8730
rect 3884 8678 3936 8730
rect 3948 8678 4000 8730
rect 4012 8678 4064 8730
rect 10472 8678 10524 8730
rect 10536 8678 10588 8730
rect 10600 8678 10652 8730
rect 10664 8678 10716 8730
rect 10728 8678 10780 8730
rect 17188 8678 17240 8730
rect 17252 8678 17304 8730
rect 17316 8678 17368 8730
rect 17380 8678 17432 8730
rect 17444 8678 17496 8730
rect 23904 8678 23956 8730
rect 23968 8678 24020 8730
rect 24032 8678 24084 8730
rect 24096 8678 24148 8730
rect 24160 8678 24212 8730
rect 4804 8576 4856 8628
rect 4160 8508 4212 8560
rect 5080 8508 5132 8560
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 4068 8440 4120 8492
rect 4528 8415 4580 8424
rect 4528 8381 4537 8415
rect 4537 8381 4571 8415
rect 4571 8381 4580 8415
rect 4528 8372 4580 8381
rect 4712 8304 4764 8356
rect 4988 8347 5040 8356
rect 4988 8313 4997 8347
rect 4997 8313 5031 8347
rect 5031 8313 5040 8347
rect 4988 8304 5040 8313
rect 6644 8508 6696 8560
rect 11244 8619 11296 8628
rect 11244 8585 11253 8619
rect 11253 8585 11287 8619
rect 11287 8585 11296 8619
rect 11244 8576 11296 8585
rect 6368 8440 6420 8492
rect 5908 8415 5960 8424
rect 5908 8381 5917 8415
rect 5917 8381 5951 8415
rect 5951 8381 5960 8415
rect 5908 8372 5960 8381
rect 7472 8415 7524 8424
rect 7472 8381 7481 8415
rect 7481 8381 7515 8415
rect 7515 8381 7524 8415
rect 7472 8372 7524 8381
rect 9588 8440 9640 8492
rect 8208 8372 8260 8424
rect 9680 8372 9732 8424
rect 11428 8415 11480 8424
rect 11428 8381 11437 8415
rect 11437 8381 11471 8415
rect 11471 8381 11480 8415
rect 11428 8372 11480 8381
rect 11612 8372 11664 8424
rect 13636 8576 13688 8628
rect 12716 8508 12768 8560
rect 17592 8576 17644 8628
rect 6092 8304 6144 8356
rect 8116 8304 8168 8356
rect 12164 8440 12216 8492
rect 12256 8440 12308 8492
rect 11888 8415 11940 8424
rect 11888 8381 11897 8415
rect 11897 8381 11931 8415
rect 11931 8381 11940 8415
rect 11888 8372 11940 8381
rect 12072 8415 12124 8424
rect 12072 8381 12082 8415
rect 12082 8381 12116 8415
rect 12116 8381 12124 8415
rect 12072 8372 12124 8381
rect 3424 8236 3476 8288
rect 4436 8279 4488 8288
rect 4436 8245 4445 8279
rect 4445 8245 4479 8279
rect 4479 8245 4488 8279
rect 4436 8236 4488 8245
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 5264 8236 5316 8245
rect 11336 8236 11388 8288
rect 12164 8304 12216 8356
rect 12256 8347 12308 8356
rect 12256 8313 12265 8347
rect 12265 8313 12299 8347
rect 12299 8313 12308 8347
rect 12256 8304 12308 8313
rect 12348 8347 12400 8356
rect 12348 8313 12357 8347
rect 12357 8313 12391 8347
rect 12391 8313 12400 8347
rect 12348 8304 12400 8313
rect 12532 8236 12584 8288
rect 13452 8372 13504 8424
rect 18144 8508 18196 8560
rect 16488 8440 16540 8492
rect 19340 8576 19392 8628
rect 19892 8576 19944 8628
rect 21180 8576 21232 8628
rect 22468 8576 22520 8628
rect 25136 8508 25188 8560
rect 17040 8372 17092 8424
rect 17776 8415 17828 8424
rect 17776 8381 17785 8415
rect 17785 8381 17819 8415
rect 17819 8381 17828 8415
rect 17776 8372 17828 8381
rect 17960 8415 18012 8424
rect 17960 8381 17969 8415
rect 17969 8381 18003 8415
rect 18003 8381 18012 8415
rect 17960 8372 18012 8381
rect 13820 8304 13872 8356
rect 13912 8347 13964 8356
rect 13912 8313 13921 8347
rect 13921 8313 13955 8347
rect 13955 8313 13964 8347
rect 13912 8304 13964 8313
rect 14004 8304 14056 8356
rect 18144 8415 18196 8424
rect 18144 8381 18153 8415
rect 18153 8381 18187 8415
rect 18187 8381 18196 8415
rect 18144 8372 18196 8381
rect 22652 8440 22704 8492
rect 13268 8236 13320 8288
rect 13544 8236 13596 8288
rect 14372 8236 14424 8288
rect 14556 8236 14608 8288
rect 16764 8236 16816 8288
rect 16948 8236 17000 8288
rect 20628 8304 20680 8356
rect 20904 8304 20956 8356
rect 23020 8415 23072 8424
rect 23020 8381 23029 8415
rect 23029 8381 23063 8415
rect 23063 8381 23072 8415
rect 23020 8372 23072 8381
rect 25780 8415 25832 8424
rect 25780 8381 25814 8415
rect 25814 8381 25832 8415
rect 25780 8372 25832 8381
rect 21272 8236 21324 8288
rect 23664 8304 23716 8356
rect 24492 8304 24544 8356
rect 24952 8304 25004 8356
rect 22376 8236 22428 8288
rect 26792 8236 26844 8288
rect 7114 8134 7166 8186
rect 7178 8134 7230 8186
rect 7242 8134 7294 8186
rect 7306 8134 7358 8186
rect 7370 8134 7422 8186
rect 13830 8134 13882 8186
rect 13894 8134 13946 8186
rect 13958 8134 14010 8186
rect 14022 8134 14074 8186
rect 14086 8134 14138 8186
rect 20546 8134 20598 8186
rect 20610 8134 20662 8186
rect 20674 8134 20726 8186
rect 20738 8134 20790 8186
rect 20802 8134 20854 8186
rect 27262 8134 27314 8186
rect 27326 8134 27378 8186
rect 27390 8134 27442 8186
rect 27454 8134 27506 8186
rect 27518 8134 27570 8186
rect 4712 8032 4764 8084
rect 5356 8032 5408 8084
rect 5908 8032 5960 8084
rect 6920 8032 6972 8084
rect 7472 8032 7524 8084
rect 8576 8032 8628 8084
rect 1492 7896 1544 7948
rect 1952 7939 2004 7948
rect 1952 7905 1961 7939
rect 1961 7905 1995 7939
rect 1995 7905 2004 7939
rect 1952 7896 2004 7905
rect 3424 7939 3476 7948
rect 3424 7905 3433 7939
rect 3433 7905 3467 7939
rect 3467 7905 3476 7939
rect 3424 7896 3476 7905
rect 4160 7964 4212 8016
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 4068 7896 4120 7905
rect 4896 7896 4948 7948
rect 6092 8007 6144 8016
rect 6092 7973 6101 8007
rect 6101 7973 6135 8007
rect 6135 7973 6144 8007
rect 6092 7964 6144 7973
rect 8300 7964 8352 8016
rect 5080 7828 5132 7880
rect 8852 7939 8904 7948
rect 8852 7905 8861 7939
rect 8861 7905 8895 7939
rect 8895 7905 8904 7939
rect 8852 7896 8904 7905
rect 9588 8032 9640 8084
rect 9404 7939 9456 7948
rect 9404 7905 9413 7939
rect 9413 7905 9447 7939
rect 9447 7905 9456 7939
rect 9404 7896 9456 7905
rect 12532 8032 12584 8084
rect 12624 8032 12676 8084
rect 10876 7964 10928 8016
rect 16304 8032 16356 8084
rect 18144 8032 18196 8084
rect 7196 7828 7248 7880
rect 8760 7828 8812 7880
rect 11336 7939 11388 7948
rect 11336 7905 11345 7939
rect 11345 7905 11379 7939
rect 11379 7905 11388 7939
rect 11336 7896 11388 7905
rect 11520 7939 11572 7948
rect 11520 7905 11527 7939
rect 11527 7905 11572 7939
rect 11520 7896 11572 7905
rect 12164 7896 12216 7948
rect 12348 7939 12400 7948
rect 12348 7905 12382 7939
rect 12382 7905 12400 7939
rect 12348 7896 12400 7905
rect 12716 7896 12768 7948
rect 13728 7939 13780 7948
rect 13728 7905 13735 7939
rect 13735 7905 13780 7939
rect 11704 7828 11756 7880
rect 13728 7896 13780 7905
rect 14372 7964 14424 8016
rect 13912 7939 13964 7948
rect 13912 7905 13921 7939
rect 13921 7905 13955 7939
rect 13955 7905 13964 7939
rect 13912 7896 13964 7905
rect 14004 7939 14056 7948
rect 14004 7905 14018 7939
rect 14018 7905 14052 7939
rect 14052 7905 14056 7939
rect 14004 7896 14056 7905
rect 14556 7939 14608 7948
rect 14556 7905 14565 7939
rect 14565 7905 14599 7939
rect 14599 7905 14608 7939
rect 14556 7896 14608 7905
rect 5172 7760 5224 7812
rect 11612 7760 11664 7812
rect 4068 7692 4120 7744
rect 5264 7692 5316 7744
rect 6000 7692 6052 7744
rect 10048 7735 10100 7744
rect 10048 7701 10057 7735
rect 10057 7701 10091 7735
rect 10091 7701 10100 7735
rect 10048 7692 10100 7701
rect 12716 7692 12768 7744
rect 13544 7692 13596 7744
rect 15936 7828 15988 7880
rect 16120 7760 16172 7812
rect 17776 7964 17828 8016
rect 20352 8032 20404 8084
rect 20444 8032 20496 8084
rect 23020 8032 23072 8084
rect 23664 8075 23716 8084
rect 23664 8041 23673 8075
rect 23673 8041 23707 8075
rect 23707 8041 23716 8075
rect 23664 8032 23716 8041
rect 25136 8032 25188 8084
rect 17040 7896 17092 7948
rect 17868 7896 17920 7948
rect 19800 7939 19852 7948
rect 19800 7905 19809 7939
rect 19809 7905 19843 7939
rect 19843 7905 19852 7939
rect 19800 7896 19852 7905
rect 20352 7896 20404 7948
rect 20628 7939 20680 7948
rect 20628 7905 20637 7939
rect 20637 7905 20671 7939
rect 20671 7905 20680 7939
rect 20628 7896 20680 7905
rect 22100 7964 22152 8016
rect 20904 7896 20956 7948
rect 22376 7939 22428 7948
rect 22376 7905 22394 7939
rect 22394 7905 22428 7939
rect 22376 7896 22428 7905
rect 22652 7939 22704 7948
rect 22652 7905 22661 7939
rect 22661 7905 22695 7939
rect 22695 7905 22704 7939
rect 22652 7896 22704 7905
rect 23020 7939 23072 7948
rect 23020 7905 23029 7939
rect 23029 7905 23063 7939
rect 23063 7905 23072 7939
rect 23020 7896 23072 7905
rect 23204 7939 23256 7948
rect 23204 7905 23213 7939
rect 23213 7905 23247 7939
rect 23247 7905 23256 7939
rect 23204 7896 23256 7905
rect 16856 7828 16908 7880
rect 18420 7760 18472 7812
rect 19984 7760 20036 7812
rect 21088 7760 21140 7812
rect 21272 7803 21324 7812
rect 21272 7769 21281 7803
rect 21281 7769 21315 7803
rect 21315 7769 21324 7803
rect 21272 7760 21324 7769
rect 14832 7692 14884 7744
rect 19064 7692 19116 7744
rect 24860 7896 24912 7948
rect 24952 7939 25004 7948
rect 24952 7905 24961 7939
rect 24961 7905 24995 7939
rect 24995 7905 25004 7939
rect 24952 7896 25004 7905
rect 25596 7939 25648 7948
rect 25596 7905 25605 7939
rect 25605 7905 25639 7939
rect 25639 7905 25648 7939
rect 25596 7896 25648 7905
rect 26976 7964 27028 8016
rect 26792 7939 26844 7948
rect 26792 7905 26801 7939
rect 26801 7905 26835 7939
rect 26835 7905 26844 7939
rect 26792 7896 26844 7905
rect 25228 7828 25280 7880
rect 26056 7828 26108 7880
rect 24768 7760 24820 7812
rect 22468 7692 22520 7744
rect 25044 7692 25096 7744
rect 25964 7760 26016 7812
rect 25688 7735 25740 7744
rect 25688 7701 25697 7735
rect 25697 7701 25731 7735
rect 25731 7701 25740 7735
rect 25688 7692 25740 7701
rect 25872 7692 25924 7744
rect 3756 7590 3808 7642
rect 3820 7590 3872 7642
rect 3884 7590 3936 7642
rect 3948 7590 4000 7642
rect 4012 7590 4064 7642
rect 10472 7590 10524 7642
rect 10536 7590 10588 7642
rect 10600 7590 10652 7642
rect 10664 7590 10716 7642
rect 10728 7590 10780 7642
rect 17188 7590 17240 7642
rect 17252 7590 17304 7642
rect 17316 7590 17368 7642
rect 17380 7590 17432 7642
rect 17444 7590 17496 7642
rect 23904 7590 23956 7642
rect 23968 7590 24020 7642
rect 24032 7590 24084 7642
rect 24096 7590 24148 7642
rect 24160 7590 24212 7642
rect 4528 7488 4580 7540
rect 5172 7531 5224 7540
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 5356 7488 5408 7540
rect 4896 7463 4948 7472
rect 4896 7429 4905 7463
rect 4905 7429 4939 7463
rect 4939 7429 4948 7463
rect 4896 7420 4948 7429
rect 1952 7352 2004 7404
rect 4804 7352 4856 7404
rect 5540 7352 5592 7404
rect 4252 7284 4304 7336
rect 4436 7216 4488 7268
rect 5264 7327 5316 7336
rect 5264 7293 5273 7327
rect 5273 7293 5307 7327
rect 5307 7293 5316 7327
rect 5264 7284 5316 7293
rect 6920 7488 6972 7540
rect 7196 7531 7248 7540
rect 7196 7497 7205 7531
rect 7205 7497 7239 7531
rect 7239 7497 7248 7531
rect 7196 7488 7248 7497
rect 12348 7531 12400 7540
rect 12348 7497 12357 7531
rect 12357 7497 12391 7531
rect 12391 7497 12400 7531
rect 12348 7488 12400 7497
rect 15936 7531 15988 7540
rect 15936 7497 15945 7531
rect 15945 7497 15979 7531
rect 15979 7497 15988 7531
rect 15936 7488 15988 7497
rect 20628 7488 20680 7540
rect 21088 7488 21140 7540
rect 23020 7488 23072 7540
rect 23204 7488 23256 7540
rect 25596 7488 25648 7540
rect 26056 7531 26108 7540
rect 26056 7497 26065 7531
rect 26065 7497 26099 7531
rect 26099 7497 26108 7531
rect 26056 7488 26108 7497
rect 6828 7284 6880 7336
rect 9404 7352 9456 7404
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 5908 7216 5960 7268
rect 5816 7148 5868 7200
rect 9680 7284 9732 7336
rect 13912 7420 13964 7472
rect 13544 7395 13596 7404
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 18696 7420 18748 7472
rect 11704 7284 11756 7336
rect 12256 7284 12308 7336
rect 12624 7284 12676 7336
rect 12808 7284 12860 7336
rect 13176 7284 13228 7336
rect 13636 7216 13688 7268
rect 12624 7148 12676 7200
rect 13176 7148 13228 7200
rect 14372 7148 14424 7200
rect 14556 7327 14608 7336
rect 14556 7293 14565 7327
rect 14565 7293 14599 7327
rect 14599 7293 14608 7327
rect 14556 7284 14608 7293
rect 14832 7327 14884 7336
rect 14832 7293 14866 7327
rect 14866 7293 14884 7327
rect 14832 7284 14884 7293
rect 16028 7327 16080 7336
rect 16028 7293 16037 7327
rect 16037 7293 16071 7327
rect 16071 7293 16080 7327
rect 16028 7284 16080 7293
rect 16856 7352 16908 7404
rect 20996 7420 21048 7472
rect 17040 7284 17092 7336
rect 17592 7284 17644 7336
rect 16304 7259 16356 7268
rect 16304 7225 16313 7259
rect 16313 7225 16347 7259
rect 16347 7225 16356 7259
rect 16304 7216 16356 7225
rect 16396 7259 16448 7268
rect 16396 7225 16405 7259
rect 16405 7225 16439 7259
rect 16439 7225 16448 7259
rect 16396 7216 16448 7225
rect 16856 7216 16908 7268
rect 17960 7327 18012 7336
rect 17960 7293 17969 7327
rect 17969 7293 18003 7327
rect 18003 7293 18012 7327
rect 17960 7284 18012 7293
rect 22468 7463 22520 7472
rect 22468 7429 22477 7463
rect 22477 7429 22511 7463
rect 22511 7429 22520 7463
rect 22468 7420 22520 7429
rect 25872 7420 25924 7472
rect 19340 7216 19392 7268
rect 15568 7148 15620 7200
rect 17592 7148 17644 7200
rect 17776 7148 17828 7200
rect 17960 7148 18012 7200
rect 19892 7148 19944 7200
rect 21548 7327 21600 7336
rect 21548 7293 21557 7327
rect 21557 7293 21591 7327
rect 21591 7293 21600 7327
rect 21548 7284 21600 7293
rect 21640 7327 21692 7336
rect 21640 7293 21649 7327
rect 21649 7293 21683 7327
rect 21683 7293 21692 7327
rect 21640 7284 21692 7293
rect 24768 7352 24820 7404
rect 22376 7216 22428 7268
rect 24584 7284 24636 7336
rect 25044 7327 25096 7336
rect 25044 7293 25053 7327
rect 25053 7293 25087 7327
rect 25087 7293 25096 7327
rect 25044 7284 25096 7293
rect 25136 7284 25188 7336
rect 25872 7327 25924 7336
rect 25872 7293 25881 7327
rect 25881 7293 25915 7327
rect 25915 7293 25924 7327
rect 25872 7284 25924 7293
rect 26608 7327 26660 7336
rect 26608 7293 26617 7327
rect 26617 7293 26651 7327
rect 26651 7293 26660 7327
rect 26608 7284 26660 7293
rect 23020 7148 23072 7200
rect 24308 7148 24360 7200
rect 24584 7191 24636 7200
rect 24584 7157 24593 7191
rect 24593 7157 24627 7191
rect 24627 7157 24636 7191
rect 24584 7148 24636 7157
rect 7114 7046 7166 7098
rect 7178 7046 7230 7098
rect 7242 7046 7294 7098
rect 7306 7046 7358 7098
rect 7370 7046 7422 7098
rect 13830 7046 13882 7098
rect 13894 7046 13946 7098
rect 13958 7046 14010 7098
rect 14022 7046 14074 7098
rect 14086 7046 14138 7098
rect 20546 7046 20598 7098
rect 20610 7046 20662 7098
rect 20674 7046 20726 7098
rect 20738 7046 20790 7098
rect 20802 7046 20854 7098
rect 27262 7046 27314 7098
rect 27326 7046 27378 7098
rect 27390 7046 27442 7098
rect 27454 7046 27506 7098
rect 27518 7046 27570 7098
rect 5632 6944 5684 6996
rect 5908 6987 5960 6996
rect 5908 6953 5917 6987
rect 5917 6953 5951 6987
rect 5951 6953 5960 6987
rect 5908 6944 5960 6953
rect 8668 6987 8720 6996
rect 8668 6953 8677 6987
rect 8677 6953 8711 6987
rect 8711 6953 8720 6987
rect 8668 6944 8720 6953
rect 8852 6944 8904 6996
rect 9680 6944 9732 6996
rect 10876 6944 10928 6996
rect 12532 6944 12584 6996
rect 15292 6944 15344 6996
rect 16396 6944 16448 6996
rect 21640 6944 21692 6996
rect 24860 6944 24912 6996
rect 25872 6944 25924 6996
rect 26608 6944 26660 6996
rect 7932 6876 7984 6928
rect 5540 6808 5592 6860
rect 5816 6851 5868 6860
rect 5816 6817 5825 6851
rect 5825 6817 5859 6851
rect 5859 6817 5868 6851
rect 5816 6808 5868 6817
rect 6000 6851 6052 6860
rect 6000 6817 6009 6851
rect 6009 6817 6043 6851
rect 6043 6817 6052 6851
rect 6000 6808 6052 6817
rect 8116 6851 8168 6860
rect 8116 6817 8125 6851
rect 8125 6817 8159 6851
rect 8159 6817 8168 6851
rect 8116 6808 8168 6817
rect 8576 6808 8628 6860
rect 9036 6851 9088 6860
rect 9036 6817 9045 6851
rect 9045 6817 9079 6851
rect 9079 6817 9088 6851
rect 9036 6808 9088 6817
rect 10048 6808 10100 6860
rect 11888 6851 11940 6860
rect 11888 6817 11897 6851
rect 11897 6817 11931 6851
rect 11931 6817 11940 6851
rect 11888 6808 11940 6817
rect 11980 6851 12032 6860
rect 11980 6817 11989 6851
rect 11989 6817 12023 6851
rect 12023 6817 12032 6851
rect 11980 6808 12032 6817
rect 12164 6851 12216 6860
rect 12164 6817 12173 6851
rect 12173 6817 12207 6851
rect 12207 6817 12216 6851
rect 12164 6808 12216 6817
rect 13636 6876 13688 6928
rect 12624 6851 12676 6860
rect 12624 6817 12633 6851
rect 12633 6817 12667 6851
rect 12667 6817 12676 6851
rect 12624 6808 12676 6817
rect 12716 6851 12768 6860
rect 12716 6817 12725 6851
rect 12725 6817 12759 6851
rect 12759 6817 12768 6851
rect 12716 6808 12768 6817
rect 12900 6851 12952 6860
rect 12900 6817 12909 6851
rect 12909 6817 12943 6851
rect 12943 6817 12952 6851
rect 12900 6808 12952 6817
rect 12992 6808 13044 6860
rect 7104 6740 7156 6792
rect 11244 6740 11296 6792
rect 12808 6740 12860 6792
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 14096 6808 14148 6860
rect 14832 6851 14884 6860
rect 14832 6817 14866 6851
rect 14866 6817 14884 6851
rect 14832 6808 14884 6817
rect 24584 6919 24636 6928
rect 13544 6740 13596 6749
rect 14556 6783 14608 6792
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 17960 6808 18012 6860
rect 24584 6885 24618 6919
rect 24618 6885 24636 6919
rect 24584 6876 24636 6885
rect 19340 6851 19392 6860
rect 19340 6817 19349 6851
rect 19349 6817 19383 6851
rect 19383 6817 19392 6851
rect 19340 6808 19392 6817
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 16856 6740 16908 6792
rect 17684 6740 17736 6792
rect 19156 6740 19208 6792
rect 12440 6672 12492 6724
rect 5356 6604 5408 6656
rect 6828 6647 6880 6656
rect 6828 6613 6837 6647
rect 6837 6613 6871 6647
rect 6871 6613 6880 6647
rect 6828 6604 6880 6613
rect 10968 6604 11020 6656
rect 12256 6604 12308 6656
rect 15200 6604 15252 6656
rect 16304 6604 16356 6656
rect 20996 6808 21048 6860
rect 21456 6808 21508 6860
rect 25596 6808 25648 6860
rect 23296 6783 23348 6792
rect 23296 6749 23305 6783
rect 23305 6749 23339 6783
rect 23339 6749 23348 6783
rect 23296 6740 23348 6749
rect 24308 6783 24360 6792
rect 24308 6749 24317 6783
rect 24317 6749 24351 6783
rect 24351 6749 24360 6783
rect 24308 6740 24360 6749
rect 26792 6740 26844 6792
rect 26976 6783 27028 6792
rect 26976 6749 26985 6783
rect 26985 6749 27019 6783
rect 27019 6749 27028 6783
rect 26976 6740 27028 6749
rect 18972 6604 19024 6656
rect 21732 6604 21784 6656
rect 3756 6502 3808 6554
rect 3820 6502 3872 6554
rect 3884 6502 3936 6554
rect 3948 6502 4000 6554
rect 4012 6502 4064 6554
rect 10472 6502 10524 6554
rect 10536 6502 10588 6554
rect 10600 6502 10652 6554
rect 10664 6502 10716 6554
rect 10728 6502 10780 6554
rect 17188 6502 17240 6554
rect 17252 6502 17304 6554
rect 17316 6502 17368 6554
rect 17380 6502 17432 6554
rect 17444 6502 17496 6554
rect 23904 6502 23956 6554
rect 23968 6502 24020 6554
rect 24032 6502 24084 6554
rect 24096 6502 24148 6554
rect 24160 6502 24212 6554
rect 5540 6443 5592 6452
rect 5540 6409 5549 6443
rect 5549 6409 5583 6443
rect 5583 6409 5592 6443
rect 5540 6400 5592 6409
rect 6092 6400 6144 6452
rect 6644 6443 6696 6452
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 7104 6443 7156 6452
rect 7104 6409 7113 6443
rect 7113 6409 7147 6443
rect 7147 6409 7156 6443
rect 7104 6400 7156 6409
rect 7564 6400 7616 6452
rect 7932 6400 7984 6452
rect 13360 6400 13412 6452
rect 14832 6400 14884 6452
rect 17684 6400 17736 6452
rect 6000 6332 6052 6384
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 6276 6332 6328 6384
rect 11980 6332 12032 6384
rect 17592 6332 17644 6384
rect 21272 6400 21324 6452
rect 4252 6128 4304 6180
rect 5908 6239 5960 6248
rect 5908 6205 5917 6239
rect 5917 6205 5951 6239
rect 5951 6205 5960 6239
rect 5908 6196 5960 6205
rect 6920 6196 6972 6248
rect 8300 6264 8352 6316
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 11796 6264 11848 6316
rect 6184 6060 6236 6112
rect 6736 6128 6788 6180
rect 7564 6239 7616 6248
rect 7564 6205 7573 6239
rect 7573 6205 7607 6239
rect 7607 6205 7616 6239
rect 7564 6196 7616 6205
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 8668 6196 8720 6205
rect 9864 6239 9916 6248
rect 9864 6205 9873 6239
rect 9873 6205 9907 6239
rect 9907 6205 9916 6239
rect 9864 6196 9916 6205
rect 11520 6196 11572 6248
rect 11888 6239 11940 6248
rect 11888 6205 11897 6239
rect 11897 6205 11931 6239
rect 11931 6205 11940 6239
rect 11888 6196 11940 6205
rect 11980 6239 12032 6248
rect 11980 6205 11989 6239
rect 11989 6205 12023 6239
rect 12023 6205 12032 6239
rect 11980 6196 12032 6205
rect 12256 6264 12308 6316
rect 17040 6264 17092 6316
rect 9036 6128 9088 6180
rect 11336 6128 11388 6180
rect 12348 6196 12400 6248
rect 14372 6239 14424 6248
rect 14372 6205 14381 6239
rect 14381 6205 14415 6239
rect 14415 6205 14424 6239
rect 14372 6196 14424 6205
rect 14648 6239 14700 6248
rect 14648 6205 14657 6239
rect 14657 6205 14691 6239
rect 14691 6205 14700 6239
rect 14648 6196 14700 6205
rect 14924 6196 14976 6248
rect 12256 6128 12308 6180
rect 7748 6103 7800 6112
rect 7748 6069 7757 6103
rect 7757 6069 7791 6103
rect 7791 6069 7800 6103
rect 7748 6060 7800 6069
rect 8392 6060 8444 6112
rect 8576 6060 8628 6112
rect 9588 6103 9640 6112
rect 9588 6069 9597 6103
rect 9597 6069 9631 6103
rect 9631 6069 9640 6103
rect 9588 6060 9640 6069
rect 9680 6060 9732 6112
rect 11612 6060 11664 6112
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 11796 6060 11848 6112
rect 14556 6128 14608 6180
rect 16580 6196 16632 6248
rect 18696 6264 18748 6316
rect 16120 6128 16172 6180
rect 15384 6060 15436 6112
rect 18972 6239 19024 6248
rect 18972 6205 18981 6239
rect 18981 6205 19015 6239
rect 19015 6205 19024 6239
rect 18972 6196 19024 6205
rect 19064 6239 19116 6248
rect 19064 6205 19073 6239
rect 19073 6205 19107 6239
rect 19107 6205 19116 6239
rect 19064 6196 19116 6205
rect 21732 6264 21784 6316
rect 19248 6128 19300 6180
rect 21640 6239 21692 6248
rect 21640 6205 21649 6239
rect 21649 6205 21683 6239
rect 21683 6205 21692 6239
rect 21640 6196 21692 6205
rect 23296 6400 23348 6452
rect 26976 6400 27028 6452
rect 21916 6332 21968 6384
rect 22100 6332 22152 6384
rect 22376 6264 22428 6316
rect 22100 6239 22152 6248
rect 22100 6205 22112 6239
rect 22112 6205 22146 6239
rect 22146 6205 22152 6239
rect 22100 6196 22152 6205
rect 24308 6264 24360 6316
rect 22376 6128 22428 6180
rect 24400 6239 24452 6248
rect 24400 6205 24409 6239
rect 24409 6205 24443 6239
rect 24443 6205 24452 6239
rect 24400 6196 24452 6205
rect 25688 6196 25740 6248
rect 17224 6103 17276 6112
rect 17224 6069 17233 6103
rect 17233 6069 17267 6103
rect 17267 6069 17276 6103
rect 17224 6060 17276 6069
rect 19340 6060 19392 6112
rect 20352 6060 20404 6112
rect 20444 6060 20496 6112
rect 22192 6060 22244 6112
rect 23204 6060 23256 6112
rect 23480 6060 23532 6112
rect 7114 5958 7166 6010
rect 7178 5958 7230 6010
rect 7242 5958 7294 6010
rect 7306 5958 7358 6010
rect 7370 5958 7422 6010
rect 13830 5958 13882 6010
rect 13894 5958 13946 6010
rect 13958 5958 14010 6010
rect 14022 5958 14074 6010
rect 14086 5958 14138 6010
rect 20546 5958 20598 6010
rect 20610 5958 20662 6010
rect 20674 5958 20726 6010
rect 20738 5958 20790 6010
rect 20802 5958 20854 6010
rect 27262 5958 27314 6010
rect 27326 5958 27378 6010
rect 27390 5958 27442 6010
rect 27454 5958 27506 6010
rect 27518 5958 27570 6010
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 6000 5856 6052 5908
rect 6184 5788 6236 5840
rect 6736 5856 6788 5908
rect 8852 5856 8904 5908
rect 10140 5899 10192 5908
rect 10140 5865 10149 5899
rect 10149 5865 10183 5899
rect 10183 5865 10192 5899
rect 10140 5856 10192 5865
rect 11980 5856 12032 5908
rect 13360 5856 13412 5908
rect 5356 5763 5408 5772
rect 5356 5729 5374 5763
rect 5374 5729 5408 5763
rect 5356 5720 5408 5729
rect 6092 5720 6144 5772
rect 6920 5788 6972 5840
rect 8024 5788 8076 5840
rect 7380 5720 7432 5772
rect 9680 5788 9732 5840
rect 8576 5763 8628 5772
rect 8576 5729 8610 5763
rect 8610 5729 8628 5763
rect 8576 5720 8628 5729
rect 8944 5720 8996 5772
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 6644 5627 6696 5636
rect 6644 5593 6653 5627
rect 6653 5593 6687 5627
rect 6687 5593 6696 5627
rect 6644 5584 6696 5593
rect 10968 5763 11020 5772
rect 10968 5729 10977 5763
rect 10977 5729 11011 5763
rect 11011 5729 11020 5763
rect 10968 5720 11020 5729
rect 11704 5788 11756 5840
rect 12072 5788 12124 5840
rect 12164 5788 12216 5840
rect 11336 5720 11388 5772
rect 11428 5763 11480 5772
rect 11428 5729 11437 5763
rect 11437 5729 11471 5763
rect 11471 5729 11480 5763
rect 11428 5720 11480 5729
rect 11520 5763 11572 5772
rect 11520 5729 11529 5763
rect 11529 5729 11563 5763
rect 11563 5729 11572 5763
rect 11520 5720 11572 5729
rect 11612 5763 11664 5772
rect 11612 5729 11621 5763
rect 11621 5729 11655 5763
rect 11655 5729 11664 5763
rect 11612 5720 11664 5729
rect 13636 5695 13688 5704
rect 13636 5661 13645 5695
rect 13645 5661 13679 5695
rect 13679 5661 13688 5695
rect 13636 5652 13688 5661
rect 14924 5899 14976 5908
rect 14924 5865 14933 5899
rect 14933 5865 14967 5899
rect 14967 5865 14976 5899
rect 14924 5856 14976 5865
rect 16120 5899 16172 5908
rect 16120 5865 16129 5899
rect 16129 5865 16163 5899
rect 16163 5865 16172 5899
rect 16120 5856 16172 5865
rect 17224 5856 17276 5908
rect 19708 5856 19760 5908
rect 20444 5856 20496 5908
rect 16948 5788 17000 5840
rect 14372 5763 14424 5772
rect 14372 5729 14381 5763
rect 14381 5729 14415 5763
rect 14415 5729 14424 5763
rect 14372 5720 14424 5729
rect 14464 5763 14516 5772
rect 14464 5729 14473 5763
rect 14473 5729 14507 5763
rect 14507 5729 14516 5763
rect 14464 5720 14516 5729
rect 14648 5763 14700 5772
rect 14648 5729 14657 5763
rect 14657 5729 14691 5763
rect 14691 5729 14700 5763
rect 14648 5720 14700 5729
rect 15200 5763 15252 5772
rect 15200 5729 15209 5763
rect 15209 5729 15243 5763
rect 15243 5729 15252 5763
rect 15200 5720 15252 5729
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 15384 5763 15436 5772
rect 15384 5729 15393 5763
rect 15393 5729 15427 5763
rect 15427 5729 15436 5763
rect 15384 5720 15436 5729
rect 15568 5763 15620 5772
rect 15568 5729 15577 5763
rect 15577 5729 15611 5763
rect 15611 5729 15620 5763
rect 15568 5720 15620 5729
rect 5816 5559 5868 5568
rect 5816 5525 5825 5559
rect 5825 5525 5859 5559
rect 5859 5525 5868 5559
rect 5816 5516 5868 5525
rect 6276 5516 6328 5568
rect 6736 5516 6788 5568
rect 8944 5516 8996 5568
rect 9036 5516 9088 5568
rect 11244 5627 11296 5636
rect 11244 5593 11253 5627
rect 11253 5593 11287 5627
rect 11287 5593 11296 5627
rect 11244 5584 11296 5593
rect 11336 5516 11388 5568
rect 11520 5516 11572 5568
rect 17500 5763 17552 5772
rect 17500 5729 17509 5763
rect 17509 5729 17543 5763
rect 17543 5729 17552 5763
rect 17500 5720 17552 5729
rect 17592 5720 17644 5772
rect 18052 5763 18104 5772
rect 18052 5729 18061 5763
rect 18061 5729 18095 5763
rect 18095 5729 18104 5763
rect 18052 5720 18104 5729
rect 18144 5763 18196 5772
rect 18144 5729 18153 5763
rect 18153 5729 18187 5763
rect 18187 5729 18196 5763
rect 18144 5720 18196 5729
rect 18972 5763 19024 5772
rect 18972 5729 18982 5763
rect 18982 5729 19016 5763
rect 19016 5729 19024 5763
rect 18972 5720 19024 5729
rect 19156 5763 19208 5772
rect 19156 5729 19165 5763
rect 19165 5729 19199 5763
rect 19199 5729 19208 5763
rect 19156 5720 19208 5729
rect 19248 5763 19300 5772
rect 19248 5729 19257 5763
rect 19257 5729 19291 5763
rect 19291 5729 19300 5763
rect 19248 5720 19300 5729
rect 20904 5788 20956 5840
rect 20352 5763 20404 5772
rect 20352 5729 20361 5763
rect 20361 5729 20395 5763
rect 20395 5729 20404 5763
rect 20352 5720 20404 5729
rect 21548 5856 21600 5908
rect 21916 5899 21968 5908
rect 21916 5865 21925 5899
rect 21925 5865 21959 5899
rect 21959 5865 21968 5899
rect 21916 5856 21968 5865
rect 24400 5856 24452 5908
rect 21548 5763 21600 5772
rect 21548 5729 21557 5763
rect 21557 5729 21591 5763
rect 21591 5729 21600 5763
rect 21548 5720 21600 5729
rect 19708 5652 19760 5704
rect 20076 5652 20128 5704
rect 21824 5720 21876 5772
rect 20260 5584 20312 5636
rect 13544 5516 13596 5568
rect 18972 5516 19024 5568
rect 19984 5516 20036 5568
rect 20996 5559 21048 5568
rect 20996 5525 21005 5559
rect 21005 5525 21039 5559
rect 21039 5525 21048 5559
rect 20996 5516 21048 5525
rect 21548 5584 21600 5636
rect 22376 5763 22428 5772
rect 22376 5729 22385 5763
rect 22385 5729 22419 5763
rect 22419 5729 22428 5763
rect 22376 5720 22428 5729
rect 23756 5788 23808 5840
rect 24308 5788 24360 5840
rect 24676 5788 24728 5840
rect 22652 5763 22704 5772
rect 22652 5729 22661 5763
rect 22661 5729 22695 5763
rect 22695 5729 22704 5763
rect 22652 5720 22704 5729
rect 22744 5763 22796 5772
rect 22744 5729 22753 5763
rect 22753 5729 22787 5763
rect 22787 5729 22796 5763
rect 22744 5720 22796 5729
rect 22100 5652 22152 5704
rect 23020 5720 23072 5772
rect 25412 5695 25464 5704
rect 25412 5661 25421 5695
rect 25421 5661 25455 5695
rect 25455 5661 25464 5695
rect 25412 5652 25464 5661
rect 22744 5584 22796 5636
rect 22652 5516 22704 5568
rect 23112 5516 23164 5568
rect 3756 5414 3808 5466
rect 3820 5414 3872 5466
rect 3884 5414 3936 5466
rect 3948 5414 4000 5466
rect 4012 5414 4064 5466
rect 10472 5414 10524 5466
rect 10536 5414 10588 5466
rect 10600 5414 10652 5466
rect 10664 5414 10716 5466
rect 10728 5414 10780 5466
rect 17188 5414 17240 5466
rect 17252 5414 17304 5466
rect 17316 5414 17368 5466
rect 17380 5414 17432 5466
rect 17444 5414 17496 5466
rect 23904 5414 23956 5466
rect 23968 5414 24020 5466
rect 24032 5414 24084 5466
rect 24096 5414 24148 5466
rect 24160 5414 24212 5466
rect 5908 5312 5960 5364
rect 6644 5312 6696 5364
rect 7380 5355 7432 5364
rect 7380 5321 7389 5355
rect 7389 5321 7423 5355
rect 7423 5321 7432 5355
rect 7380 5312 7432 5321
rect 8392 5312 8444 5364
rect 8668 5312 8720 5364
rect 11428 5312 11480 5364
rect 12348 5312 12400 5364
rect 6368 5244 6420 5296
rect 8852 5176 8904 5228
rect 4620 5151 4672 5160
rect 4620 5117 4629 5151
rect 4629 5117 4663 5151
rect 4663 5117 4672 5151
rect 4620 5108 4672 5117
rect 5816 5108 5868 5160
rect 7564 5108 7616 5160
rect 8024 5108 8076 5160
rect 8392 5083 8444 5092
rect 8392 5049 8401 5083
rect 8401 5049 8435 5083
rect 8435 5049 8444 5083
rect 8392 5040 8444 5049
rect 9036 5151 9088 5160
rect 9036 5117 9045 5151
rect 9045 5117 9079 5151
rect 9079 5117 9088 5151
rect 9036 5108 9088 5117
rect 11152 5244 11204 5296
rect 11704 5244 11756 5296
rect 13636 5312 13688 5364
rect 18052 5312 18104 5364
rect 19064 5312 19116 5364
rect 20076 5355 20128 5364
rect 20076 5321 20085 5355
rect 20085 5321 20119 5355
rect 20119 5321 20128 5355
rect 20076 5312 20128 5321
rect 21640 5312 21692 5364
rect 25412 5312 25464 5364
rect 13636 5176 13688 5228
rect 14096 5176 14148 5228
rect 11612 5108 11664 5160
rect 12992 5108 13044 5160
rect 16580 5176 16632 5228
rect 12256 5040 12308 5092
rect 12440 5083 12492 5092
rect 12440 5049 12458 5083
rect 12458 5049 12492 5083
rect 12440 5040 12492 5049
rect 16856 5108 16908 5160
rect 17960 5108 18012 5160
rect 18512 5108 18564 5160
rect 19892 5108 19944 5160
rect 7748 4972 7800 5024
rect 11336 4972 11388 5024
rect 16948 5040 17000 5092
rect 18972 5083 19024 5092
rect 18972 5049 19006 5083
rect 19006 5049 19024 5083
rect 18972 5040 19024 5049
rect 19340 5040 19392 5092
rect 20260 5108 20312 5160
rect 21732 5244 21784 5296
rect 23756 5244 23808 5296
rect 20996 5108 21048 5160
rect 21088 5151 21140 5160
rect 21088 5117 21097 5151
rect 21097 5117 21131 5151
rect 21131 5117 21140 5151
rect 21088 5108 21140 5117
rect 21272 5108 21324 5160
rect 22928 5151 22980 5160
rect 22928 5117 22937 5151
rect 22937 5117 22971 5151
rect 22971 5117 22980 5151
rect 22928 5108 22980 5117
rect 23112 5151 23164 5160
rect 23112 5117 23121 5151
rect 23121 5117 23155 5151
rect 23155 5117 23164 5151
rect 23112 5108 23164 5117
rect 23204 5151 23256 5160
rect 23204 5117 23213 5151
rect 23213 5117 23247 5151
rect 23247 5117 23256 5151
rect 23204 5108 23256 5117
rect 23480 5108 23532 5160
rect 24676 5108 24728 5160
rect 25872 5151 25924 5160
rect 25872 5117 25881 5151
rect 25881 5117 25915 5151
rect 25915 5117 25924 5151
rect 25872 5108 25924 5117
rect 21364 5040 21416 5092
rect 22376 5040 22428 5092
rect 23572 5040 23624 5092
rect 14464 4972 14516 5024
rect 14648 4972 14700 5024
rect 15568 4972 15620 5024
rect 17500 4972 17552 5024
rect 19984 4972 20036 5024
rect 20260 4972 20312 5024
rect 20536 4972 20588 5024
rect 20904 4972 20956 5024
rect 22836 4972 22888 5024
rect 7114 4870 7166 4922
rect 7178 4870 7230 4922
rect 7242 4870 7294 4922
rect 7306 4870 7358 4922
rect 7370 4870 7422 4922
rect 13830 4870 13882 4922
rect 13894 4870 13946 4922
rect 13958 4870 14010 4922
rect 14022 4870 14074 4922
rect 14086 4870 14138 4922
rect 20546 4870 20598 4922
rect 20610 4870 20662 4922
rect 20674 4870 20726 4922
rect 20738 4870 20790 4922
rect 20802 4870 20854 4922
rect 27262 4870 27314 4922
rect 27326 4870 27378 4922
rect 27390 4870 27442 4922
rect 27454 4870 27506 4922
rect 27518 4870 27570 4922
rect 7564 4811 7616 4820
rect 7564 4777 7573 4811
rect 7573 4777 7607 4811
rect 7607 4777 7616 4811
rect 7564 4768 7616 4777
rect 8300 4768 8352 4820
rect 5264 4675 5316 4684
rect 5264 4641 5273 4675
rect 5273 4641 5307 4675
rect 5307 4641 5316 4675
rect 5264 4632 5316 4641
rect 18604 4768 18656 4820
rect 6276 4675 6328 4684
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 6368 4632 6420 4684
rect 7472 4675 7524 4684
rect 7472 4641 7481 4675
rect 7481 4641 7515 4675
rect 7515 4641 7524 4675
rect 7472 4632 7524 4641
rect 6552 4564 6604 4616
rect 7840 4675 7892 4684
rect 7840 4641 7849 4675
rect 7849 4641 7883 4675
rect 7883 4641 7892 4675
rect 7840 4632 7892 4641
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 9956 4700 10008 4752
rect 12440 4700 12492 4752
rect 9036 4675 9088 4684
rect 9036 4641 9045 4675
rect 9045 4641 9079 4675
rect 9079 4641 9088 4675
rect 9036 4632 9088 4641
rect 12900 4700 12952 4752
rect 12716 4632 12768 4684
rect 12808 4675 12860 4684
rect 12808 4641 12817 4675
rect 12817 4641 12851 4675
rect 12851 4641 12860 4675
rect 12808 4632 12860 4641
rect 13176 4675 13228 4684
rect 13176 4641 13185 4675
rect 13185 4641 13219 4675
rect 13219 4641 13228 4675
rect 13176 4632 13228 4641
rect 13636 4632 13688 4684
rect 14004 4675 14056 4684
rect 14004 4641 14013 4675
rect 14013 4641 14047 4675
rect 14047 4641 14056 4675
rect 14004 4632 14056 4641
rect 9588 4564 9640 4616
rect 14464 4632 14516 4684
rect 14832 4675 14884 4684
rect 14832 4641 14866 4675
rect 14866 4641 14884 4675
rect 14832 4632 14884 4641
rect 15200 4632 15252 4684
rect 8024 4496 8076 4548
rect 9128 4496 9180 4548
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 11520 4496 11572 4548
rect 11796 4496 11848 4548
rect 12808 4496 12860 4548
rect 13636 4496 13688 4548
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 17224 4675 17276 4684
rect 17224 4641 17233 4675
rect 17233 4641 17267 4675
rect 17267 4641 17276 4675
rect 17224 4632 17276 4641
rect 19432 4743 19484 4752
rect 19432 4709 19441 4743
rect 19441 4709 19475 4743
rect 19475 4709 19484 4743
rect 19432 4700 19484 4709
rect 22652 4768 22704 4820
rect 22928 4768 22980 4820
rect 17500 4675 17552 4684
rect 17500 4641 17509 4675
rect 17509 4641 17543 4675
rect 17543 4641 17552 4675
rect 17500 4632 17552 4641
rect 19984 4632 20036 4684
rect 20260 4675 20312 4684
rect 20260 4641 20269 4675
rect 20269 4641 20303 4675
rect 20303 4641 20312 4675
rect 20260 4632 20312 4641
rect 20352 4675 20404 4684
rect 20352 4641 20362 4675
rect 20362 4641 20396 4675
rect 20396 4641 20404 4675
rect 20352 4632 20404 4641
rect 20904 4632 20956 4684
rect 22376 4675 22428 4684
rect 22376 4641 22385 4675
rect 22385 4641 22419 4675
rect 22419 4641 22428 4675
rect 22376 4632 22428 4641
rect 4896 4428 4948 4480
rect 8576 4428 8628 4480
rect 8668 4471 8720 4480
rect 8668 4437 8677 4471
rect 8677 4437 8711 4471
rect 8711 4437 8720 4471
rect 8668 4428 8720 4437
rect 9312 4428 9364 4480
rect 10876 4428 10928 4480
rect 11336 4471 11388 4480
rect 11336 4437 11345 4471
rect 11345 4437 11379 4471
rect 11379 4437 11388 4471
rect 11336 4428 11388 4437
rect 15292 4428 15344 4480
rect 18512 4428 18564 4480
rect 21088 4428 21140 4480
rect 21364 4428 21416 4480
rect 21916 4428 21968 4480
rect 22744 4607 22796 4616
rect 22744 4573 22753 4607
rect 22753 4573 22787 4607
rect 22787 4573 22796 4607
rect 22744 4564 22796 4573
rect 23756 4768 23808 4820
rect 25872 4768 25924 4820
rect 23664 4675 23716 4684
rect 23664 4641 23673 4675
rect 23673 4641 23707 4675
rect 23707 4641 23716 4675
rect 23664 4632 23716 4641
rect 23572 4564 23624 4616
rect 24308 4428 24360 4480
rect 3756 4326 3808 4378
rect 3820 4326 3872 4378
rect 3884 4326 3936 4378
rect 3948 4326 4000 4378
rect 4012 4326 4064 4378
rect 10472 4326 10524 4378
rect 10536 4326 10588 4378
rect 10600 4326 10652 4378
rect 10664 4326 10716 4378
rect 10728 4326 10780 4378
rect 17188 4326 17240 4378
rect 17252 4326 17304 4378
rect 17316 4326 17368 4378
rect 17380 4326 17432 4378
rect 17444 4326 17496 4378
rect 23904 4326 23956 4378
rect 23968 4326 24020 4378
rect 24032 4326 24084 4378
rect 24096 4326 24148 4378
rect 24160 4326 24212 4378
rect 8576 4267 8628 4276
rect 8576 4233 8585 4267
rect 8585 4233 8619 4267
rect 8619 4233 8628 4267
rect 8576 4224 8628 4233
rect 9036 4224 9088 4276
rect 9956 4224 10008 4276
rect 8116 4199 8168 4208
rect 8116 4165 8125 4199
rect 8125 4165 8159 4199
rect 8159 4165 8168 4199
rect 8116 4156 8168 4165
rect 6552 4088 6604 4140
rect 4620 4063 4672 4072
rect 4620 4029 4629 4063
rect 4629 4029 4663 4063
rect 4663 4029 4672 4063
rect 4620 4020 4672 4029
rect 4896 3995 4948 4004
rect 4896 3961 4930 3995
rect 4930 3961 4948 3995
rect 4896 3952 4948 3961
rect 6368 4020 6420 4072
rect 7472 4020 7524 4072
rect 7932 4131 7984 4140
rect 7932 4097 7941 4131
rect 7941 4097 7975 4131
rect 7975 4097 7984 4131
rect 7932 4088 7984 4097
rect 12532 4224 12584 4276
rect 13176 4224 13228 4276
rect 14832 4267 14884 4276
rect 14832 4233 14841 4267
rect 14841 4233 14875 4267
rect 14875 4233 14884 4267
rect 14832 4224 14884 4233
rect 12256 4156 12308 4208
rect 13544 4156 13596 4208
rect 8300 4020 8352 4072
rect 6828 3952 6880 4004
rect 7012 3884 7064 3936
rect 7748 3952 7800 4004
rect 8392 3995 8444 4004
rect 8392 3961 8401 3995
rect 8401 3961 8435 3995
rect 8435 3961 8444 3995
rect 8392 3952 8444 3961
rect 7564 3927 7616 3936
rect 7564 3893 7573 3927
rect 7573 3893 7607 3927
rect 7607 3893 7616 3927
rect 7564 3884 7616 3893
rect 7932 3927 7984 3936
rect 7932 3893 7941 3927
rect 7941 3893 7975 3927
rect 7975 3893 7984 3927
rect 7932 3884 7984 3893
rect 8208 3884 8260 3936
rect 8576 3927 8628 3936
rect 8576 3893 8601 3927
rect 8601 3893 8628 3927
rect 9128 4020 9180 4072
rect 9312 4063 9364 4072
rect 9312 4029 9346 4063
rect 9346 4029 9364 4063
rect 9312 4020 9364 4029
rect 10876 4020 10928 4072
rect 11612 4020 11664 4072
rect 8576 3884 8628 3893
rect 12716 4063 12768 4072
rect 12716 4029 12725 4063
rect 12725 4029 12759 4063
rect 12759 4029 12768 4063
rect 12716 4020 12768 4029
rect 13636 4020 13688 4072
rect 14188 4020 14240 4072
rect 14464 4020 14516 4072
rect 15016 4020 15068 4072
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 15384 4088 15436 4140
rect 15292 4063 15344 4072
rect 15292 4029 15301 4063
rect 15301 4029 15335 4063
rect 15335 4029 15344 4063
rect 15292 4020 15344 4029
rect 15660 4088 15712 4140
rect 15568 4020 15620 4072
rect 19984 4088 20036 4140
rect 21732 4224 21784 4276
rect 22744 4224 22796 4276
rect 22836 4224 22888 4276
rect 23296 4267 23348 4276
rect 23296 4233 23305 4267
rect 23305 4233 23339 4267
rect 23339 4233 23348 4267
rect 23296 4224 23348 4233
rect 22652 4156 22704 4208
rect 23204 4088 23256 4140
rect 23664 4088 23716 4140
rect 16488 4020 16540 4072
rect 18512 4020 18564 4072
rect 21088 4063 21140 4072
rect 21088 4029 21122 4063
rect 21122 4029 21140 4063
rect 21088 4020 21140 4029
rect 22192 4020 22244 4072
rect 22560 4063 22612 4072
rect 22560 4029 22567 4063
rect 22567 4029 22612 4063
rect 22560 4020 22612 4029
rect 22836 4063 22888 4072
rect 22836 4029 22850 4063
rect 22850 4029 22884 4063
rect 22884 4029 22888 4063
rect 22836 4020 22888 4029
rect 23020 4020 23072 4072
rect 23296 4020 23348 4072
rect 24124 4063 24176 4072
rect 24124 4029 24133 4063
rect 24133 4029 24167 4063
rect 24167 4029 24176 4063
rect 24124 4020 24176 4029
rect 24308 4063 24360 4072
rect 24308 4029 24353 4063
rect 24353 4029 24360 4063
rect 24308 4020 24360 4029
rect 16764 3952 16816 4004
rect 17592 3952 17644 4004
rect 19064 3952 19116 4004
rect 22652 3995 22704 4004
rect 22652 3961 22661 3995
rect 22661 3961 22695 3995
rect 22695 3961 22704 3995
rect 22652 3952 22704 3961
rect 13176 3884 13228 3936
rect 14924 3884 14976 3936
rect 15476 3884 15528 3936
rect 17960 3884 18012 3936
rect 18144 3884 18196 3936
rect 20076 3884 20128 3936
rect 20260 3884 20312 3936
rect 23204 3884 23256 3936
rect 23388 3884 23440 3936
rect 24400 3884 24452 3936
rect 25136 4063 25188 4072
rect 25136 4029 25145 4063
rect 25145 4029 25179 4063
rect 25179 4029 25188 4063
rect 25136 4020 25188 4029
rect 24676 3884 24728 3936
rect 7114 3782 7166 3834
rect 7178 3782 7230 3834
rect 7242 3782 7294 3834
rect 7306 3782 7358 3834
rect 7370 3782 7422 3834
rect 13830 3782 13882 3834
rect 13894 3782 13946 3834
rect 13958 3782 14010 3834
rect 14022 3782 14074 3834
rect 14086 3782 14138 3834
rect 20546 3782 20598 3834
rect 20610 3782 20662 3834
rect 20674 3782 20726 3834
rect 20738 3782 20790 3834
rect 20802 3782 20854 3834
rect 27262 3782 27314 3834
rect 27326 3782 27378 3834
rect 27390 3782 27442 3834
rect 27454 3782 27506 3834
rect 27518 3782 27570 3834
rect 5264 3680 5316 3732
rect 6276 3680 6328 3732
rect 8300 3723 8352 3732
rect 8300 3689 8309 3723
rect 8309 3689 8343 3723
rect 8343 3689 8352 3723
rect 8300 3680 8352 3689
rect 12256 3680 12308 3732
rect 7104 3655 7156 3664
rect 7104 3621 7138 3655
rect 7138 3621 7156 3655
rect 7104 3612 7156 3621
rect 7564 3612 7616 3664
rect 8668 3612 8720 3664
rect 6552 3544 6604 3596
rect 8208 3544 8260 3596
rect 12992 3612 13044 3664
rect 13176 3655 13228 3664
rect 13176 3621 13185 3655
rect 13185 3621 13219 3655
rect 13219 3621 13228 3655
rect 13176 3612 13228 3621
rect 15384 3680 15436 3732
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 9956 3544 10008 3553
rect 11612 3544 11664 3596
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 13452 3587 13504 3596
rect 13452 3553 13461 3587
rect 13461 3553 13495 3587
rect 13495 3553 13504 3587
rect 13452 3544 13504 3553
rect 13544 3587 13596 3596
rect 13544 3553 13553 3587
rect 13553 3553 13587 3587
rect 13587 3553 13596 3587
rect 13544 3544 13596 3553
rect 14188 3544 14240 3596
rect 14740 3587 14792 3596
rect 14740 3553 14749 3587
rect 14749 3553 14783 3587
rect 14783 3553 14792 3587
rect 14740 3544 14792 3553
rect 5632 3408 5684 3460
rect 13268 3476 13320 3528
rect 9680 3451 9732 3460
rect 9680 3417 9689 3451
rect 9689 3417 9723 3451
rect 9723 3417 9732 3451
rect 15016 3587 15068 3596
rect 15016 3553 15025 3587
rect 15025 3553 15059 3587
rect 15059 3553 15068 3587
rect 15016 3544 15068 3553
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 17592 3723 17644 3732
rect 17592 3689 17601 3723
rect 17601 3689 17635 3723
rect 17635 3689 17644 3723
rect 17592 3680 17644 3689
rect 18420 3680 18472 3732
rect 19064 3723 19116 3732
rect 19064 3689 19073 3723
rect 19073 3689 19107 3723
rect 19107 3689 19116 3723
rect 19064 3680 19116 3689
rect 25136 3680 25188 3732
rect 25596 3723 25648 3732
rect 25596 3689 25605 3723
rect 25605 3689 25639 3723
rect 25639 3689 25648 3723
rect 25596 3680 25648 3689
rect 15660 3587 15712 3596
rect 15660 3553 15669 3587
rect 15669 3553 15703 3587
rect 15703 3553 15712 3587
rect 15660 3544 15712 3553
rect 16028 3544 16080 3596
rect 16488 3612 16540 3664
rect 18052 3612 18104 3664
rect 17960 3544 18012 3596
rect 17868 3476 17920 3528
rect 18604 3587 18656 3596
rect 18604 3553 18613 3587
rect 18613 3553 18647 3587
rect 18647 3553 18656 3587
rect 18604 3544 18656 3553
rect 20260 3587 20312 3596
rect 20260 3553 20269 3587
rect 20269 3553 20303 3587
rect 20303 3553 20312 3587
rect 20260 3544 20312 3553
rect 21548 3587 21600 3596
rect 21548 3553 21557 3587
rect 21557 3553 21591 3587
rect 21591 3553 21600 3587
rect 21548 3544 21600 3553
rect 21732 3587 21784 3596
rect 21732 3553 21741 3587
rect 21741 3553 21775 3587
rect 21775 3553 21784 3587
rect 21732 3544 21784 3553
rect 21916 3587 21968 3596
rect 21916 3553 21925 3587
rect 21925 3553 21959 3587
rect 21959 3553 21968 3587
rect 23388 3612 23440 3664
rect 24676 3612 24728 3664
rect 21916 3544 21968 3553
rect 22376 3587 22428 3596
rect 22376 3553 22385 3587
rect 22385 3553 22419 3587
rect 22419 3553 22428 3587
rect 22376 3544 22428 3553
rect 24492 3587 24544 3596
rect 24492 3553 24526 3587
rect 24526 3553 24544 3587
rect 24492 3544 24544 3553
rect 22468 3476 22520 3528
rect 23112 3476 23164 3528
rect 9680 3408 9732 3417
rect 7748 3340 7800 3392
rect 21824 3408 21876 3460
rect 12900 3383 12952 3392
rect 12900 3349 12909 3383
rect 12909 3349 12943 3383
rect 12943 3349 12952 3383
rect 12900 3340 12952 3349
rect 13636 3340 13688 3392
rect 18052 3340 18104 3392
rect 20352 3383 20404 3392
rect 20352 3349 20361 3383
rect 20361 3349 20395 3383
rect 20395 3349 20404 3383
rect 20352 3340 20404 3349
rect 21916 3340 21968 3392
rect 22284 3340 22336 3392
rect 23756 3340 23808 3392
rect 3756 3238 3808 3290
rect 3820 3238 3872 3290
rect 3884 3238 3936 3290
rect 3948 3238 4000 3290
rect 4012 3238 4064 3290
rect 10472 3238 10524 3290
rect 10536 3238 10588 3290
rect 10600 3238 10652 3290
rect 10664 3238 10716 3290
rect 10728 3238 10780 3290
rect 17188 3238 17240 3290
rect 17252 3238 17304 3290
rect 17316 3238 17368 3290
rect 17380 3238 17432 3290
rect 17444 3238 17496 3290
rect 23904 3238 23956 3290
rect 23968 3238 24020 3290
rect 24032 3238 24084 3290
rect 24096 3238 24148 3290
rect 24160 3238 24212 3290
rect 6368 3179 6420 3188
rect 6368 3145 6377 3179
rect 6377 3145 6411 3179
rect 6411 3145 6420 3179
rect 6368 3136 6420 3145
rect 6460 3068 6512 3120
rect 2596 3000 2648 3052
rect 4528 3000 4580 3052
rect 8576 3136 8628 3188
rect 8668 3136 8720 3188
rect 11796 3179 11848 3188
rect 11796 3145 11805 3179
rect 11805 3145 11839 3179
rect 11839 3145 11848 3179
rect 11796 3136 11848 3145
rect 12440 3179 12492 3188
rect 12440 3145 12449 3179
rect 12449 3145 12483 3179
rect 12483 3145 12492 3179
rect 12440 3136 12492 3145
rect 12992 3136 13044 3188
rect 14188 3136 14240 3188
rect 15660 3136 15712 3188
rect 16764 3136 16816 3188
rect 21548 3136 21600 3188
rect 21640 3136 21692 3188
rect 22376 3136 22428 3188
rect 23296 3136 23348 3188
rect 8208 3111 8260 3120
rect 8208 3077 8217 3111
rect 8217 3077 8251 3111
rect 8251 3077 8260 3111
rect 8208 3068 8260 3077
rect 13452 3068 13504 3120
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 12532 3000 12584 3052
rect 13360 3043 13412 3052
rect 13360 3009 13369 3043
rect 13369 3009 13403 3043
rect 13403 3009 13412 3043
rect 13360 3000 13412 3009
rect 18052 3000 18104 3052
rect 22008 3068 22060 3120
rect 24492 3136 24544 3188
rect 22468 3000 22520 3052
rect 9680 2932 9732 2984
rect 7564 2864 7616 2916
rect 7748 2864 7800 2916
rect 9128 2907 9180 2916
rect 9128 2873 9137 2907
rect 9137 2873 9171 2907
rect 9171 2873 9180 2907
rect 9128 2864 9180 2873
rect 11428 2975 11480 2984
rect 11428 2941 11437 2975
rect 11437 2941 11471 2975
rect 11471 2941 11480 2975
rect 11428 2932 11480 2941
rect 12256 2932 12308 2984
rect 12992 2932 13044 2984
rect 15292 2932 15344 2984
rect 17868 2932 17920 2984
rect 18144 2932 18196 2984
rect 18420 2975 18472 2984
rect 18420 2941 18429 2975
rect 18429 2941 18463 2975
rect 18463 2941 18472 2975
rect 18420 2932 18472 2941
rect 18696 2975 18748 2984
rect 18696 2941 18705 2975
rect 18705 2941 18739 2975
rect 18739 2941 18748 2975
rect 18696 2932 18748 2941
rect 19984 2932 20036 2984
rect 21824 2932 21876 2984
rect 8116 2796 8168 2848
rect 10048 2796 10100 2848
rect 11336 2796 11388 2848
rect 20352 2864 20404 2916
rect 24032 2975 24084 2984
rect 24032 2941 24041 2975
rect 24041 2941 24075 2975
rect 24075 2941 24084 2975
rect 24032 2932 24084 2941
rect 25596 3068 25648 3120
rect 25688 3000 25740 3052
rect 25228 2864 25280 2916
rect 13176 2796 13228 2848
rect 13728 2796 13780 2848
rect 15200 2796 15252 2848
rect 16120 2796 16172 2848
rect 17224 2796 17276 2848
rect 19340 2839 19392 2848
rect 19340 2805 19349 2839
rect 19349 2805 19383 2839
rect 19383 2805 19392 2839
rect 19340 2796 19392 2805
rect 21456 2796 21508 2848
rect 22192 2796 22244 2848
rect 22836 2796 22888 2848
rect 23204 2796 23256 2848
rect 23388 2796 23440 2848
rect 24492 2796 24544 2848
rect 7114 2694 7166 2746
rect 7178 2694 7230 2746
rect 7242 2694 7294 2746
rect 7306 2694 7358 2746
rect 7370 2694 7422 2746
rect 13830 2694 13882 2746
rect 13894 2694 13946 2746
rect 13958 2694 14010 2746
rect 14022 2694 14074 2746
rect 14086 2694 14138 2746
rect 20546 2694 20598 2746
rect 20610 2694 20662 2746
rect 20674 2694 20726 2746
rect 20738 2694 20790 2746
rect 20802 2694 20854 2746
rect 27262 2694 27314 2746
rect 27326 2694 27378 2746
rect 27390 2694 27442 2746
rect 27454 2694 27506 2746
rect 27518 2694 27570 2746
rect 7564 2635 7616 2644
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 11244 2592 11296 2644
rect 11520 2592 11572 2644
rect 12256 2592 12308 2644
rect 13360 2592 13412 2644
rect 7472 2499 7524 2508
rect 7472 2465 7481 2499
rect 7481 2465 7515 2499
rect 7515 2465 7524 2499
rect 7472 2456 7524 2465
rect 7932 2456 7984 2508
rect 10048 2499 10100 2508
rect 10048 2465 10057 2499
rect 10057 2465 10091 2499
rect 10091 2465 10100 2499
rect 10048 2456 10100 2465
rect 11060 2499 11112 2508
rect 11060 2465 11069 2499
rect 11069 2465 11103 2499
rect 11103 2465 11112 2499
rect 11060 2456 11112 2465
rect 10324 2320 10376 2372
rect 10968 2388 11020 2440
rect 11428 2456 11480 2508
rect 12532 2567 12584 2576
rect 12532 2533 12541 2567
rect 12541 2533 12575 2567
rect 12575 2533 12584 2567
rect 12532 2524 12584 2533
rect 13268 2524 13320 2576
rect 14188 2592 14240 2644
rect 16120 2592 16172 2644
rect 17224 2592 17276 2644
rect 13912 2524 13964 2576
rect 14280 2524 14332 2576
rect 11336 2388 11388 2440
rect 11980 2388 12032 2440
rect 12256 2499 12308 2508
rect 12256 2465 12265 2499
rect 12265 2465 12299 2499
rect 12299 2465 12308 2499
rect 12256 2456 12308 2465
rect 12716 2456 12768 2508
rect 12992 2456 13044 2508
rect 14096 2499 14148 2508
rect 14096 2465 14105 2499
rect 14105 2465 14139 2499
rect 14139 2465 14148 2499
rect 14096 2456 14148 2465
rect 14740 2499 14792 2508
rect 14740 2465 14749 2499
rect 14749 2465 14783 2499
rect 14783 2465 14792 2499
rect 14740 2456 14792 2465
rect 15016 2499 15068 2508
rect 15016 2465 15025 2499
rect 15025 2465 15059 2499
rect 15059 2465 15068 2499
rect 15016 2456 15068 2465
rect 12992 2320 13044 2372
rect 9680 2252 9732 2304
rect 10140 2295 10192 2304
rect 10140 2261 10149 2295
rect 10149 2261 10183 2295
rect 10183 2261 10192 2295
rect 10140 2252 10192 2261
rect 13268 2252 13320 2304
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13360 2252 13412 2261
rect 13544 2295 13596 2304
rect 13544 2261 13553 2295
rect 13553 2261 13587 2295
rect 13587 2261 13596 2295
rect 13544 2252 13596 2261
rect 13636 2252 13688 2304
rect 14372 2388 14424 2440
rect 15384 2499 15436 2508
rect 15384 2465 15393 2499
rect 15393 2465 15427 2499
rect 15427 2465 15436 2499
rect 15384 2456 15436 2465
rect 14648 2320 14700 2372
rect 15016 2320 15068 2372
rect 16672 2431 16724 2440
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 17224 2499 17276 2508
rect 17224 2465 17233 2499
rect 17233 2465 17267 2499
rect 17267 2465 17276 2499
rect 17224 2456 17276 2465
rect 17868 2592 17920 2644
rect 19432 2592 19484 2644
rect 19340 2524 19392 2576
rect 21732 2592 21784 2644
rect 22376 2592 22428 2644
rect 22652 2592 22704 2644
rect 23020 2592 23072 2644
rect 24032 2592 24084 2644
rect 18052 2456 18104 2508
rect 18052 2320 18104 2372
rect 14464 2252 14516 2304
rect 15108 2252 15160 2304
rect 15936 2252 15988 2304
rect 16856 2295 16908 2304
rect 16856 2261 16865 2295
rect 16865 2261 16899 2295
rect 16899 2261 16908 2295
rect 16856 2252 16908 2261
rect 17592 2252 17644 2304
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 21456 2499 21508 2508
rect 21456 2465 21460 2499
rect 21460 2465 21494 2499
rect 21494 2465 21508 2499
rect 21456 2456 21508 2465
rect 21824 2499 21876 2508
rect 21824 2465 21832 2499
rect 21832 2465 21866 2499
rect 21866 2465 21876 2499
rect 21824 2456 21876 2465
rect 22008 2456 22060 2508
rect 22192 2499 22244 2508
rect 22192 2465 22196 2499
rect 22196 2465 22230 2499
rect 22230 2465 22244 2499
rect 22192 2456 22244 2465
rect 22284 2499 22336 2508
rect 22284 2465 22293 2499
rect 22293 2465 22327 2499
rect 22327 2465 22336 2499
rect 22284 2456 22336 2465
rect 22376 2499 22428 2508
rect 22376 2465 22385 2499
rect 22385 2465 22419 2499
rect 22419 2465 22428 2499
rect 22376 2456 22428 2465
rect 22468 2499 22520 2508
rect 22468 2465 22513 2499
rect 22513 2465 22520 2499
rect 22468 2456 22520 2465
rect 22652 2320 22704 2372
rect 23020 2499 23072 2508
rect 23020 2465 23029 2499
rect 23029 2465 23063 2499
rect 23063 2465 23072 2499
rect 23020 2456 23072 2465
rect 23204 2499 23256 2508
rect 23204 2465 23218 2499
rect 23218 2465 23252 2499
rect 23252 2465 23256 2499
rect 23204 2456 23256 2465
rect 25688 2524 25740 2576
rect 23756 2388 23808 2440
rect 19984 2295 20036 2304
rect 19984 2261 19993 2295
rect 19993 2261 20027 2295
rect 20027 2261 20036 2295
rect 19984 2252 20036 2261
rect 21732 2252 21784 2304
rect 22100 2252 22152 2304
rect 23388 2320 23440 2372
rect 25964 2388 26016 2440
rect 23020 2252 23072 2304
rect 24308 2252 24360 2304
rect 25228 2252 25280 2304
rect 25872 2252 25924 2304
rect 3756 2150 3808 2202
rect 3820 2150 3872 2202
rect 3884 2150 3936 2202
rect 3948 2150 4000 2202
rect 4012 2150 4064 2202
rect 10472 2150 10524 2202
rect 10536 2150 10588 2202
rect 10600 2150 10652 2202
rect 10664 2150 10716 2202
rect 10728 2150 10780 2202
rect 17188 2150 17240 2202
rect 17252 2150 17304 2202
rect 17316 2150 17368 2202
rect 17380 2150 17432 2202
rect 17444 2150 17496 2202
rect 23904 2150 23956 2202
rect 23968 2150 24020 2202
rect 24032 2150 24084 2202
rect 24096 2150 24148 2202
rect 24160 2150 24212 2202
rect 9680 2091 9732 2100
rect 9680 2057 9689 2091
rect 9689 2057 9723 2091
rect 9723 2057 9732 2091
rect 9680 2048 9732 2057
rect 10140 1865 10192 1896
rect 9220 1751 9272 1760
rect 9220 1717 9229 1751
rect 9229 1717 9263 1751
rect 9263 1717 9272 1751
rect 9220 1708 9272 1717
rect 10140 1844 10150 1865
rect 10150 1844 10184 1865
rect 10184 1844 10192 1865
rect 9864 1819 9916 1828
rect 9864 1785 9873 1819
rect 9873 1785 9907 1819
rect 9907 1785 9916 1819
rect 9864 1776 9916 1785
rect 10968 2048 11020 2100
rect 11060 2048 11112 2100
rect 13544 2048 13596 2100
rect 14280 2091 14332 2100
rect 14280 2057 14289 2091
rect 14289 2057 14323 2091
rect 14323 2057 14332 2091
rect 14280 2048 14332 2057
rect 16672 2048 16724 2100
rect 18696 2048 18748 2100
rect 10600 1912 10652 1964
rect 10508 1887 10560 1896
rect 10508 1853 10517 1887
rect 10517 1853 10551 1887
rect 10551 1853 10560 1887
rect 10508 1844 10560 1853
rect 11520 1912 11572 1964
rect 15660 1955 15712 1964
rect 15660 1921 15669 1955
rect 15669 1921 15703 1955
rect 15703 1921 15712 1955
rect 15660 1912 15712 1921
rect 18144 1980 18196 2032
rect 18420 1980 18472 2032
rect 22284 2048 22336 2100
rect 22376 2048 22428 2100
rect 12348 1844 12400 1896
rect 13636 1844 13688 1896
rect 11152 1751 11204 1760
rect 11152 1717 11161 1751
rect 11161 1717 11195 1751
rect 11195 1717 11204 1751
rect 11152 1708 11204 1717
rect 11980 1751 12032 1760
rect 11980 1717 11989 1751
rect 11989 1717 12023 1751
rect 12023 1717 12032 1751
rect 11980 1708 12032 1717
rect 13176 1708 13228 1760
rect 14372 1887 14424 1896
rect 14372 1853 14381 1887
rect 14381 1853 14415 1887
rect 14415 1853 14424 1887
rect 14372 1844 14424 1853
rect 14464 1887 14516 1896
rect 14464 1853 14473 1887
rect 14473 1853 14507 1887
rect 14507 1853 14516 1887
rect 14464 1844 14516 1853
rect 14648 1887 14700 1896
rect 14648 1853 14657 1887
rect 14657 1853 14691 1887
rect 14691 1853 14700 1887
rect 14648 1844 14700 1853
rect 14372 1708 14424 1760
rect 14832 1751 14884 1760
rect 14832 1717 14841 1751
rect 14841 1717 14875 1751
rect 14875 1717 14884 1751
rect 14832 1708 14884 1717
rect 15108 1887 15160 1896
rect 15108 1853 15117 1887
rect 15117 1853 15151 1887
rect 15151 1853 15160 1887
rect 15108 1844 15160 1853
rect 15200 1887 15252 1896
rect 15200 1853 15209 1887
rect 15209 1853 15243 1887
rect 15243 1853 15252 1887
rect 15200 1844 15252 1853
rect 15936 1887 15988 1896
rect 15936 1853 15970 1887
rect 15970 1853 15988 1887
rect 15936 1844 15988 1853
rect 17868 1887 17920 1896
rect 17868 1853 17877 1887
rect 17877 1853 17911 1887
rect 17911 1853 17920 1887
rect 17868 1844 17920 1853
rect 18052 1887 18104 1896
rect 18052 1853 18061 1887
rect 18061 1853 18095 1887
rect 18095 1853 18104 1887
rect 18052 1844 18104 1853
rect 18144 1887 18196 1896
rect 18144 1853 18153 1887
rect 18153 1853 18187 1887
rect 18187 1853 18196 1887
rect 18144 1844 18196 1853
rect 19984 1980 20036 2032
rect 19892 1912 19944 1964
rect 22192 1955 22244 1964
rect 22192 1921 22201 1955
rect 22201 1921 22235 1955
rect 22235 1921 22244 1955
rect 22192 1912 22244 1921
rect 22376 1912 22428 1964
rect 18972 1887 19024 1896
rect 18972 1853 18981 1887
rect 18981 1853 19015 1887
rect 19015 1853 19024 1887
rect 18972 1844 19024 1853
rect 19064 1887 19116 1896
rect 19064 1853 19073 1887
rect 19073 1853 19107 1887
rect 19107 1853 19116 1887
rect 19064 1844 19116 1853
rect 17960 1776 18012 1828
rect 19432 1844 19484 1896
rect 20904 1844 20956 1896
rect 22836 1887 22888 1896
rect 22836 1853 22845 1887
rect 22845 1853 22879 1887
rect 22879 1853 22888 1887
rect 22836 1844 22888 1853
rect 23388 1844 23440 1896
rect 24308 1980 24360 2032
rect 23480 1776 23532 1828
rect 24216 1819 24268 1828
rect 24216 1785 24225 1819
rect 24225 1785 24259 1819
rect 24259 1785 24268 1819
rect 24216 1776 24268 1785
rect 24492 1844 24544 1896
rect 24768 1887 24820 1896
rect 24768 1853 24775 1887
rect 24775 1853 24820 1887
rect 24768 1844 24820 1853
rect 25964 2091 26016 2100
rect 25964 2057 25973 2091
rect 25973 2057 26007 2091
rect 26007 2057 26016 2091
rect 25964 2048 26016 2057
rect 25228 1844 25280 1896
rect 15292 1708 15344 1760
rect 18696 1751 18748 1760
rect 18696 1717 18705 1751
rect 18705 1717 18739 1751
rect 18739 1717 18748 1751
rect 18696 1708 18748 1717
rect 22468 1708 22520 1760
rect 23112 1708 23164 1760
rect 25596 1887 25648 1896
rect 25596 1853 25605 1887
rect 25605 1853 25639 1887
rect 25639 1853 25648 1887
rect 25596 1844 25648 1853
rect 25688 1887 25740 1896
rect 25688 1853 25697 1887
rect 25697 1853 25731 1887
rect 25731 1853 25740 1887
rect 25688 1844 25740 1853
rect 25872 1844 25924 1896
rect 25780 1708 25832 1760
rect 26700 1751 26752 1760
rect 26700 1717 26709 1751
rect 26709 1717 26743 1751
rect 26743 1717 26752 1751
rect 26700 1708 26752 1717
rect 7114 1606 7166 1658
rect 7178 1606 7230 1658
rect 7242 1606 7294 1658
rect 7306 1606 7358 1658
rect 7370 1606 7422 1658
rect 13830 1606 13882 1658
rect 13894 1606 13946 1658
rect 13958 1606 14010 1658
rect 14022 1606 14074 1658
rect 14086 1606 14138 1658
rect 20546 1606 20598 1658
rect 20610 1606 20662 1658
rect 20674 1606 20726 1658
rect 20738 1606 20790 1658
rect 20802 1606 20854 1658
rect 27262 1606 27314 1658
rect 27326 1606 27378 1658
rect 27390 1606 27442 1658
rect 27454 1606 27506 1658
rect 27518 1606 27570 1658
rect 8392 1504 8444 1556
rect 9864 1504 9916 1556
rect 10048 1504 10100 1556
rect 10600 1504 10652 1556
rect 9220 1436 9272 1488
rect 11152 1436 11204 1488
rect 12716 1436 12768 1488
rect 14832 1504 14884 1556
rect 19616 1504 19668 1556
rect 22192 1504 22244 1556
rect 15384 1436 15436 1488
rect 16856 1436 16908 1488
rect 18512 1436 18564 1488
rect 12808 1368 12860 1420
rect 14372 1368 14424 1420
rect 11612 1164 11664 1216
rect 12348 1207 12400 1216
rect 12348 1173 12357 1207
rect 12357 1173 12391 1207
rect 12391 1173 12400 1207
rect 15016 1368 15068 1420
rect 15660 1368 15712 1420
rect 16028 1368 16080 1420
rect 19800 1368 19852 1420
rect 19892 1368 19944 1420
rect 23204 1368 23256 1420
rect 24768 1504 24820 1556
rect 26700 1368 26752 1420
rect 12348 1164 12400 1173
rect 17960 1232 18012 1284
rect 17592 1164 17644 1216
rect 17684 1207 17736 1216
rect 17684 1173 17693 1207
rect 17693 1173 17727 1207
rect 17727 1173 17736 1207
rect 17684 1164 17736 1173
rect 19340 1164 19392 1216
rect 23756 1232 23808 1284
rect 23480 1164 23532 1216
rect 3756 1062 3808 1114
rect 3820 1062 3872 1114
rect 3884 1062 3936 1114
rect 3948 1062 4000 1114
rect 4012 1062 4064 1114
rect 10472 1062 10524 1114
rect 10536 1062 10588 1114
rect 10600 1062 10652 1114
rect 10664 1062 10716 1114
rect 10728 1062 10780 1114
rect 17188 1062 17240 1114
rect 17252 1062 17304 1114
rect 17316 1062 17368 1114
rect 17380 1062 17432 1114
rect 17444 1062 17496 1114
rect 23904 1062 23956 1114
rect 23968 1062 24020 1114
rect 24032 1062 24084 1114
rect 24096 1062 24148 1114
rect 24160 1062 24212 1114
rect 12808 960 12860 1012
rect 18972 960 19024 1012
rect 19340 1003 19392 1012
rect 19340 969 19349 1003
rect 19349 969 19383 1003
rect 19383 969 19392 1003
rect 19340 960 19392 969
rect 19800 960 19852 1012
rect 22836 960 22888 1012
rect 23204 960 23256 1012
rect 25780 960 25832 1012
rect 22744 892 22796 944
rect 23296 892 23348 944
rect 17684 824 17736 876
rect 18696 867 18748 876
rect 18696 833 18705 867
rect 18705 833 18739 867
rect 18739 833 18748 867
rect 18696 824 18748 833
rect 19064 824 19116 876
rect 13360 756 13412 808
rect 19432 799 19484 808
rect 19432 765 19441 799
rect 19441 765 19475 799
rect 19475 765 19484 799
rect 19432 756 19484 765
rect 19616 799 19668 808
rect 19616 765 19625 799
rect 19625 765 19659 799
rect 19659 765 19668 799
rect 19616 756 19668 765
rect 20904 756 20956 808
rect 21640 756 21692 808
rect 21732 799 21784 808
rect 21732 765 21741 799
rect 21741 765 21775 799
rect 21775 765 21784 799
rect 21732 756 21784 765
rect 22100 756 22152 808
rect 22468 799 22520 808
rect 22468 765 22475 799
rect 22475 765 22520 799
rect 22468 756 22520 765
rect 22560 799 22612 808
rect 22560 765 22569 799
rect 22569 765 22603 799
rect 22603 765 22612 799
rect 22560 756 22612 765
rect 22652 799 22704 808
rect 22652 765 22661 799
rect 22661 765 22695 799
rect 22695 765 22704 799
rect 22652 756 22704 765
rect 22928 756 22980 808
rect 23296 799 23348 808
rect 23296 765 23305 799
rect 23305 765 23339 799
rect 23339 765 23348 799
rect 23296 756 23348 765
rect 24768 892 24820 944
rect 23480 756 23532 808
rect 22744 620 22796 672
rect 7114 518 7166 570
rect 7178 518 7230 570
rect 7242 518 7294 570
rect 7306 518 7358 570
rect 7370 518 7422 570
rect 13830 518 13882 570
rect 13894 518 13946 570
rect 13958 518 14010 570
rect 14022 518 14074 570
rect 14086 518 14138 570
rect 20546 518 20598 570
rect 20610 518 20662 570
rect 20674 518 20726 570
rect 20738 518 20790 570
rect 20802 518 20854 570
rect 27262 518 27314 570
rect 27326 518 27378 570
rect 27390 518 27442 570
rect 27454 518 27506 570
rect 27518 518 27570 570
<< metal2 >>
rect 754 17600 810 18000
rect 1398 17600 1454 18000
rect 2042 17762 2098 18000
rect 2042 17734 2176 17762
rect 2042 17600 2098 17734
rect 768 16794 796 17600
rect 756 16788 808 16794
rect 756 16730 808 16736
rect 1412 11354 1440 17600
rect 2148 17338 2176 17734
rect 2686 17600 2742 18000
rect 3330 17762 3386 18000
rect 3330 17734 3464 17762
rect 3330 17600 3386 17734
rect 2700 17338 2728 17600
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 3436 17202 3464 17734
rect 3974 17600 4030 18000
rect 4618 17600 4674 18000
rect 5262 17600 5318 18000
rect 5906 17600 5962 18000
rect 6550 17600 6606 18000
rect 7194 17762 7250 18000
rect 7194 17734 7328 17762
rect 7194 17600 7250 17734
rect 3988 17542 4016 17600
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3620 17338 3648 17478
rect 3756 17436 4064 17445
rect 3756 17434 3762 17436
rect 3818 17434 3842 17436
rect 3898 17434 3922 17436
rect 3978 17434 4002 17436
rect 4058 17434 4064 17436
rect 3818 17382 3820 17434
rect 4000 17382 4002 17434
rect 3756 17380 3762 17382
rect 3818 17380 3842 17382
rect 3898 17380 3922 17382
rect 3978 17380 4002 17382
rect 4058 17380 4064 17382
rect 3756 17371 4064 17380
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 4632 17202 4660 17600
rect 5276 17202 5304 17600
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4172 16726 4200 16934
rect 5644 16794 5672 17478
rect 5920 16794 5948 17600
rect 6564 17134 6592 17600
rect 7300 17338 7328 17734
rect 7838 17600 7894 18000
rect 8482 17600 8538 18000
rect 9126 17600 9182 18000
rect 9770 17600 9826 18000
rect 10414 17762 10470 18000
rect 10414 17734 10732 17762
rect 9956 17604 10008 17610
rect 7852 17338 7880 17600
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 6736 17264 6788 17270
rect 6736 17206 6788 17212
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6748 16998 6776 17206
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5908 16788 5960 16794
rect 5908 16730 5960 16736
rect 4160 16720 4212 16726
rect 4160 16662 4212 16668
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3252 16114 3280 16526
rect 5644 16402 5672 16730
rect 6748 16658 6776 16934
rect 7114 16892 7422 16901
rect 7114 16890 7120 16892
rect 7176 16890 7200 16892
rect 7256 16890 7280 16892
rect 7336 16890 7360 16892
rect 7416 16890 7422 16892
rect 7176 16838 7178 16890
rect 7358 16838 7360 16890
rect 7114 16836 7120 16838
rect 7176 16836 7200 16838
rect 7256 16836 7280 16838
rect 7336 16836 7360 16838
rect 7416 16836 7422 16838
rect 7114 16827 7422 16836
rect 7484 16658 7512 17138
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 5460 16374 5672 16402
rect 3756 16348 4064 16357
rect 3756 16346 3762 16348
rect 3818 16346 3842 16348
rect 3898 16346 3922 16348
rect 3978 16346 4002 16348
rect 4058 16346 4064 16348
rect 3818 16294 3820 16346
rect 4000 16294 4002 16346
rect 3756 16292 3762 16294
rect 3818 16292 3842 16294
rect 3898 16292 3922 16294
rect 3978 16292 4002 16294
rect 4058 16292 4064 16294
rect 3756 16283 4064 16292
rect 4804 16176 4856 16182
rect 5460 16130 5488 16374
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 4804 16118 4856 16124
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3344 15706 3372 15982
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 4816 15570 4844 16118
rect 5276 16102 5488 16130
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 3608 15496 3660 15502
rect 3608 15438 3660 15444
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2516 13938 2544 14214
rect 2608 14074 2636 14418
rect 3332 14340 3384 14346
rect 3332 14282 3384 14288
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2516 12238 2544 13874
rect 3344 13870 3372 14282
rect 3620 14278 3648 15438
rect 3756 15260 4064 15269
rect 3756 15258 3762 15260
rect 3818 15258 3842 15260
rect 3898 15258 3922 15260
rect 3978 15258 4002 15260
rect 4058 15258 4064 15260
rect 3818 15206 3820 15258
rect 4000 15206 4002 15258
rect 3756 15204 3762 15206
rect 3818 15204 3842 15206
rect 3898 15204 3922 15206
rect 3978 15204 4002 15206
rect 4058 15204 4064 15206
rect 3756 15195 4064 15204
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4080 14414 4108 14894
rect 4448 14482 4476 15506
rect 5000 15434 5028 15574
rect 4988 15428 5040 15434
rect 4988 15370 5040 15376
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4816 14958 4844 15302
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4894 14920 4950 14929
rect 4894 14855 4950 14864
rect 4908 14634 4936 14855
rect 4540 14618 4936 14634
rect 4528 14612 4936 14618
rect 4580 14606 4936 14612
rect 4528 14554 4580 14560
rect 4908 14482 4936 14606
rect 5000 14550 5028 15370
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 4988 14544 5040 14550
rect 4988 14486 5040 14492
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3620 12782 3648 14214
rect 3756 14172 4064 14181
rect 3756 14170 3762 14172
rect 3818 14170 3842 14172
rect 3898 14170 3922 14172
rect 3978 14170 4002 14172
rect 4058 14170 4064 14172
rect 3818 14118 3820 14170
rect 4000 14118 4002 14170
rect 3756 14116 3762 14118
rect 3818 14116 3842 14118
rect 3898 14116 3922 14118
rect 3978 14116 4002 14118
rect 4058 14116 4064 14118
rect 3756 14107 4064 14116
rect 4252 14000 4304 14006
rect 4252 13942 4304 13948
rect 4264 13462 4292 13942
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 4448 13326 4476 14418
rect 5000 14074 5028 14486
rect 5092 14414 5120 14826
rect 5276 14634 5304 16102
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5368 15366 5396 15982
rect 5460 15570 5488 16102
rect 5552 15638 5580 16186
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5368 14940 5396 15302
rect 5644 14958 5672 15982
rect 5908 15904 5960 15910
rect 5908 15846 5960 15852
rect 5920 15570 5948 15846
rect 5908 15564 5960 15570
rect 5908 15506 5960 15512
rect 6012 15162 6040 16594
rect 6840 16250 6868 16594
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6644 16176 6696 16182
rect 6644 16118 6696 16124
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6288 15706 6316 15982
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6460 15088 6512 15094
rect 6460 15030 6512 15036
rect 5448 14952 5500 14958
rect 5368 14912 5448 14940
rect 5448 14894 5500 14900
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 5276 14606 5396 14634
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 4988 14068 5040 14074
rect 4908 14028 4988 14056
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4724 13394 4752 13670
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 3756 13084 4064 13093
rect 3756 13082 3762 13084
rect 3818 13082 3842 13084
rect 3898 13082 3922 13084
rect 3978 13082 4002 13084
rect 4058 13082 4064 13084
rect 3818 13030 3820 13082
rect 4000 13030 4002 13082
rect 3756 13028 3762 13030
rect 3818 13028 3842 13030
rect 3898 13028 3922 13030
rect 3978 13028 4002 13030
rect 4058 13028 4064 13030
rect 3756 13019 4064 13028
rect 4172 12850 4200 13126
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4448 12782 4476 13262
rect 3608 12776 3660 12782
rect 3976 12776 4028 12782
rect 3660 12736 3976 12764
rect 3608 12718 3660 12724
rect 3976 12718 4028 12724
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 2792 12306 2820 12582
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 2516 10606 2544 12174
rect 3252 11694 3280 12582
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 3756 11996 4064 12005
rect 3756 11994 3762 11996
rect 3818 11994 3842 11996
rect 3898 11994 3922 11996
rect 3978 11994 4002 11996
rect 4058 11994 4064 11996
rect 3818 11942 3820 11994
rect 4000 11942 4002 11994
rect 3756 11940 3762 11942
rect 3818 11940 3842 11942
rect 3898 11940 3922 11942
rect 3978 11940 4002 11942
rect 4058 11940 4064 11942
rect 3756 11931 4064 11940
rect 4264 11898 4292 12242
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2412 10532 2464 10538
rect 2412 10474 2464 10480
rect 2424 10266 2452 10474
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2056 9722 2084 10066
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1964 9110 1992 9522
rect 2148 9450 2176 9590
rect 2240 9586 2268 9862
rect 2884 9722 2912 10066
rect 3160 9994 3188 11154
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3344 10606 3372 10950
rect 3756 10908 4064 10917
rect 3756 10906 3762 10908
rect 3818 10906 3842 10908
rect 3898 10906 3922 10908
rect 3978 10906 4002 10908
rect 4058 10906 4064 10908
rect 3818 10854 3820 10906
rect 4000 10854 4002 10906
rect 3756 10852 3762 10854
rect 3818 10852 3842 10854
rect 3898 10852 3922 10854
rect 3978 10852 4002 10854
rect 4058 10852 4064 10854
rect 3756 10843 4064 10852
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4172 10266 4200 10406
rect 4264 10266 4292 11154
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 3620 9654 3648 10134
rect 4252 10056 4304 10062
rect 4172 10004 4252 10010
rect 4172 9998 4304 10004
rect 4172 9982 4292 9998
rect 3756 9820 4064 9829
rect 3756 9818 3762 9820
rect 3818 9818 3842 9820
rect 3898 9818 3922 9820
rect 3978 9818 4002 9820
rect 4058 9818 4064 9820
rect 3818 9766 3820 9818
rect 4000 9766 4002 9818
rect 3756 9764 3762 9766
rect 3818 9764 3842 9766
rect 3898 9764 3922 9766
rect 3978 9764 4002 9766
rect 4058 9764 4064 9766
rect 3756 9755 4064 9764
rect 4172 9722 4200 9982
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 3608 9648 3660 9654
rect 3608 9590 3660 9596
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 4264 9518 4292 9862
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 2136 9444 2188 9450
rect 2136 9386 2188 9392
rect 2596 9376 2648 9382
rect 2884 9364 2912 9454
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 2648 9336 2912 9364
rect 2596 9318 2648 9324
rect 3068 9110 3096 9386
rect 3804 9178 3832 9454
rect 4264 9382 4292 9454
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 1952 9104 2004 9110
rect 1952 9046 2004 9052
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 1504 7954 1532 8910
rect 3756 8732 4064 8741
rect 3756 8730 3762 8732
rect 3818 8730 3842 8732
rect 3898 8730 3922 8732
rect 3978 8730 4002 8732
rect 4058 8730 4064 8732
rect 3818 8678 3820 8730
rect 4000 8678 4002 8730
rect 3756 8676 3762 8678
rect 3818 8676 3842 8678
rect 3898 8676 3922 8678
rect 3978 8676 4002 8678
rect 4058 8676 4064 8678
rect 3756 8667 4064 8676
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7954 3464 8230
rect 4080 7954 4108 8434
rect 4172 8022 4200 8502
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 1964 7410 1992 7890
rect 4080 7750 4108 7890
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 3756 7644 4064 7653
rect 3756 7642 3762 7644
rect 3818 7642 3842 7644
rect 3898 7642 3922 7644
rect 3978 7642 4002 7644
rect 4058 7642 4064 7644
rect 3818 7590 3820 7642
rect 4000 7590 4002 7642
rect 3756 7588 3762 7590
rect 3818 7588 3842 7590
rect 3898 7588 3922 7590
rect 3978 7588 4002 7590
rect 4058 7588 4064 7590
rect 3756 7579 4064 7588
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 4264 7342 4292 8910
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 3756 6556 4064 6565
rect 3756 6554 3762 6556
rect 3818 6554 3842 6556
rect 3898 6554 3922 6556
rect 3978 6554 4002 6556
rect 4058 6554 4064 6556
rect 3818 6502 3820 6554
rect 4000 6502 4002 6554
rect 3756 6500 3762 6502
rect 3818 6500 3842 6502
rect 3898 6500 3922 6502
rect 3978 6500 4002 6502
rect 4058 6500 4064 6502
rect 3756 6491 4064 6500
rect 4252 6180 4304 6186
rect 4252 6122 4304 6128
rect 4264 5914 4292 6122
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 3756 5468 4064 5477
rect 3756 5466 3762 5468
rect 3818 5466 3842 5468
rect 3898 5466 3922 5468
rect 3978 5466 4002 5468
rect 4058 5466 4064 5468
rect 3818 5414 3820 5466
rect 4000 5414 4002 5466
rect 3756 5412 3762 5414
rect 3818 5412 3842 5414
rect 3898 5412 3922 5414
rect 3978 5412 4002 5414
rect 4058 5412 4064 5414
rect 3756 5403 4064 5412
rect 3756 4380 4064 4389
rect 3756 4378 3762 4380
rect 3818 4378 3842 4380
rect 3898 4378 3922 4380
rect 3978 4378 4002 4380
rect 4058 4378 4064 4380
rect 3818 4326 3820 4378
rect 4000 4326 4002 4378
rect 3756 4324 3762 4326
rect 3818 4324 3842 4326
rect 3898 4324 3922 4326
rect 3978 4324 4002 4326
rect 4058 4324 4064 4326
rect 3756 4315 4064 4324
rect 846 3496 902 3505
rect 846 3431 902 3440
rect 860 400 888 3431
rect 3756 3292 4064 3301
rect 3756 3290 3762 3292
rect 3818 3290 3842 3292
rect 3898 3290 3922 3292
rect 3978 3290 4002 3292
rect 4058 3290 4064 3292
rect 3818 3238 3820 3290
rect 4000 3238 4002 3290
rect 3756 3236 3762 3238
rect 3818 3236 3842 3238
rect 3898 3236 3922 3238
rect 3978 3236 4002 3238
rect 4058 3236 4064 3238
rect 3756 3227 4064 3236
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2608 400 2636 2994
rect 3756 2204 4064 2213
rect 3756 2202 3762 2204
rect 3818 2202 3842 2204
rect 3898 2202 3922 2204
rect 3978 2202 4002 2204
rect 4058 2202 4064 2204
rect 3818 2150 3820 2202
rect 4000 2150 4002 2202
rect 3756 2148 3762 2150
rect 3818 2148 3842 2150
rect 3898 2148 3922 2150
rect 3978 2148 4002 2150
rect 4058 2148 4064 2150
rect 3756 2139 4064 2148
rect 3756 1116 4064 1125
rect 3756 1114 3762 1116
rect 3818 1114 3842 1116
rect 3898 1114 3922 1116
rect 3978 1114 4002 1116
rect 4058 1114 4064 1116
rect 3818 1062 3820 1114
rect 4000 1062 4002 1114
rect 3756 1060 3762 1062
rect 3818 1060 3842 1062
rect 3898 1060 3922 1062
rect 3978 1060 4002 1062
rect 4058 1060 4064 1062
rect 3756 1051 4064 1060
rect 4356 400 4384 11086
rect 4448 10062 4476 12718
rect 4724 12102 4752 13330
rect 4908 13326 4936 14028
rect 4988 14010 5040 14016
rect 5276 13938 5304 14418
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5368 13818 5396 14606
rect 5460 13938 5488 14894
rect 6380 14618 6408 14894
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 5814 13968 5870 13977
rect 5448 13932 5500 13938
rect 5814 13903 5870 13912
rect 5448 13874 5500 13880
rect 5828 13870 5856 13903
rect 6472 13870 6500 15030
rect 5632 13864 5684 13870
rect 5368 13790 5488 13818
rect 5632 13806 5684 13812
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 4908 12714 4936 13262
rect 5000 12986 5028 13262
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 5368 12442 5396 12718
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 5172 12096 5224 12102
rect 5460 12050 5488 13790
rect 5644 13530 5672 13806
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5736 12374 5764 13806
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 5816 12708 5868 12714
rect 5816 12650 5868 12656
rect 5828 12442 5856 12650
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 6104 12306 6132 13126
rect 6472 12306 6500 13806
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 5172 12038 5224 12044
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4448 9110 4476 9454
rect 4436 9104 4488 9110
rect 4436 9046 4488 9052
rect 4448 8838 4476 9046
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4448 7274 4476 8230
rect 4540 7546 4568 8366
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4436 7268 4488 7274
rect 4436 7210 4488 7216
rect 4632 5250 4660 11494
rect 5000 11218 5028 11630
rect 5184 11218 5212 12038
rect 5368 12022 5488 12050
rect 5368 11694 5396 12022
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6288 11694 6316 11834
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5552 11150 5580 11630
rect 6380 11626 6408 11766
rect 6656 11694 6684 16118
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7114 15804 7422 15813
rect 7114 15802 7120 15804
rect 7176 15802 7200 15804
rect 7256 15802 7280 15804
rect 7336 15802 7360 15804
rect 7416 15802 7422 15804
rect 7176 15750 7178 15802
rect 7358 15750 7360 15802
rect 7114 15748 7120 15750
rect 7176 15748 7200 15750
rect 7256 15748 7280 15750
rect 7336 15748 7360 15750
rect 7416 15748 7422 15750
rect 7114 15739 7422 15748
rect 7484 15706 7512 15914
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7576 15570 7604 16390
rect 8036 16114 8064 16526
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 8036 15638 8064 16050
rect 8128 15638 8156 16186
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 8116 15632 8168 15638
rect 8116 15574 8168 15580
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7944 15094 7972 15506
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 7114 14716 7422 14725
rect 7114 14714 7120 14716
rect 7176 14714 7200 14716
rect 7256 14714 7280 14716
rect 7336 14714 7360 14716
rect 7416 14714 7422 14716
rect 7176 14662 7178 14714
rect 7358 14662 7360 14714
rect 7114 14660 7120 14662
rect 7176 14660 7200 14662
rect 7256 14660 7280 14662
rect 7336 14660 7360 14662
rect 7416 14660 7422 14662
rect 7114 14651 7422 14660
rect 8036 14550 8064 15574
rect 8312 15162 8340 15982
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8496 15065 8524 17600
rect 9140 17338 9168 17600
rect 9784 17338 9812 17600
rect 10414 17600 10470 17734
rect 10704 17678 10732 17734
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 11058 17600 11114 18000
rect 11702 17600 11758 18000
rect 12346 17600 12402 18000
rect 12990 17600 13046 18000
rect 13634 17600 13690 18000
rect 14278 17762 14334 18000
rect 14922 17762 14978 18000
rect 14200 17734 14334 17762
rect 9956 17546 10008 17552
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9968 17202 9996 17546
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8680 16250 8708 16594
rect 8956 16250 8984 16934
rect 9416 16794 9444 17002
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9876 16794 9904 16934
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9968 16454 9996 17138
rect 10336 17134 10364 17478
rect 10472 17436 10780 17445
rect 10472 17434 10478 17436
rect 10534 17434 10558 17436
rect 10614 17434 10638 17436
rect 10694 17434 10718 17436
rect 10774 17434 10780 17436
rect 10534 17382 10536 17434
rect 10716 17382 10718 17434
rect 10472 17380 10478 17382
rect 10534 17380 10558 17382
rect 10614 17380 10638 17382
rect 10694 17380 10718 17382
rect 10774 17380 10780 17382
rect 10472 17371 10780 17380
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 11072 16794 11100 17600
rect 11716 16794 11744 17600
rect 12360 17338 12388 17600
rect 13004 17338 13032 17600
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11900 16726 11928 16934
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 11888 16720 11940 16726
rect 11888 16662 11940 16668
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 8772 15366 8800 16050
rect 9312 15972 9364 15978
rect 9312 15914 9364 15920
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8482 15056 8538 15065
rect 8482 14991 8538 15000
rect 8482 14920 8538 14929
rect 8482 14855 8538 14864
rect 6920 14544 6972 14550
rect 6920 14486 6972 14492
rect 8024 14544 8076 14550
rect 8024 14486 8076 14492
rect 6932 12986 6960 14486
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7852 13870 7880 14214
rect 8404 14006 8432 14418
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 7840 13864 7892 13870
rect 8024 13864 8076 13870
rect 7840 13806 7892 13812
rect 8022 13832 8024 13841
rect 8076 13832 8078 13841
rect 8022 13767 8078 13776
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 7114 13628 7422 13637
rect 7114 13626 7120 13628
rect 7176 13626 7200 13628
rect 7256 13626 7280 13628
rect 7336 13626 7360 13628
rect 7416 13626 7422 13628
rect 7176 13574 7178 13626
rect 7358 13574 7360 13626
rect 7114 13572 7120 13574
rect 7176 13572 7200 13574
rect 7256 13572 7280 13574
rect 7336 13572 7360 13574
rect 7416 13572 7422 13574
rect 7114 13563 7422 13572
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6748 11694 6776 12174
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6368 11620 6420 11626
rect 6368 11562 6420 11568
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4724 10130 4752 10406
rect 4908 10130 4936 10678
rect 5092 10130 5120 11018
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4816 8634 4844 9658
rect 5092 9654 5120 9862
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5092 9518 5120 9590
rect 5184 9518 5212 10066
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4724 8090 4752 8298
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4816 7410 4844 8570
rect 5000 8362 5028 9318
rect 5092 8566 5120 9318
rect 5184 9110 5212 9454
rect 5644 9178 5672 9454
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 4988 8356 5040 8362
rect 4988 8298 5040 8304
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4908 7478 4936 7890
rect 5092 7886 5120 8502
rect 5276 8294 5304 8978
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 5172 7812 5224 7818
rect 5172 7754 5224 7760
rect 5184 7546 5212 7754
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 5276 7342 5304 7686
rect 5368 7546 5396 8026
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5552 6984 5580 7346
rect 5632 6996 5684 7002
rect 5552 6956 5632 6984
rect 5632 6938 5684 6944
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 5778 5396 6598
rect 5552 6458 5580 6802
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5644 6322 5672 6938
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 4540 5222 4660 5250
rect 4540 3058 4568 5222
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4632 4078 4660 5102
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4908 4010 4936 4422
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 5276 3738 5304 4626
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5644 3466 5672 6258
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 846 0 902 400
rect 2594 0 2650 400
rect 4342 0 4398 400
rect 5736 354 5764 11494
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6828 11212 6880 11218
rect 6932 11200 6960 12922
rect 7114 12540 7422 12549
rect 7114 12538 7120 12540
rect 7176 12538 7200 12540
rect 7256 12538 7280 12540
rect 7336 12538 7360 12540
rect 7416 12538 7422 12540
rect 7176 12486 7178 12538
rect 7358 12486 7360 12538
rect 7114 12484 7120 12486
rect 7176 12484 7200 12486
rect 7256 12484 7280 12486
rect 7336 12484 7360 12486
rect 7416 12484 7422 12486
rect 7114 12475 7422 12484
rect 7944 12374 7972 13126
rect 8220 12850 8248 13738
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8404 12986 8432 13330
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 8220 12481 8248 12650
rect 8206 12472 8262 12481
rect 8206 12407 8262 12416
rect 7932 12368 7984 12374
rect 7838 12336 7894 12345
rect 7932 12310 7984 12316
rect 8496 12306 8524 14855
rect 8772 14822 8800 15302
rect 9036 15088 9088 15094
rect 9036 15030 9088 15036
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8588 14550 8616 14758
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8680 13870 8708 14758
rect 8772 13870 8800 14758
rect 8956 14618 8984 14894
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8864 13870 8892 14214
rect 9048 13870 9076 15030
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 9036 13864 9088 13870
rect 9140 13841 9168 13942
rect 9036 13806 9088 13812
rect 9126 13832 9182 13841
rect 8772 13326 8800 13806
rect 9126 13767 9182 13776
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 7838 12271 7840 12280
rect 7892 12271 7894 12280
rect 8024 12300 8076 12306
rect 7840 12242 7892 12248
rect 8024 12242 8076 12248
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 7380 12164 7432 12170
rect 7380 12106 7432 12112
rect 7392 11694 7420 12106
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7380 11688 7432 11694
rect 7472 11688 7524 11694
rect 7380 11630 7432 11636
rect 7470 11656 7472 11665
rect 7564 11688 7616 11694
rect 7524 11656 7526 11665
rect 7564 11630 7616 11636
rect 7470 11591 7526 11600
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 7024 11286 7052 11494
rect 7114 11452 7422 11461
rect 7114 11450 7120 11452
rect 7176 11450 7200 11452
rect 7256 11450 7280 11452
rect 7336 11450 7360 11452
rect 7416 11450 7422 11452
rect 7176 11398 7178 11450
rect 7358 11398 7360 11450
rect 7114 11396 7120 11398
rect 7176 11396 7200 11398
rect 7256 11396 7280 11398
rect 7336 11396 7360 11398
rect 7416 11396 7422 11398
rect 7114 11387 7422 11396
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 7484 11218 7512 11591
rect 7576 11354 7604 11630
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 6880 11172 6960 11200
rect 6828 11154 6880 11160
rect 6012 10606 6040 11154
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6380 10130 6408 10542
rect 6932 10130 6960 11172
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7114 10364 7422 10373
rect 7114 10362 7120 10364
rect 7176 10362 7200 10364
rect 7256 10362 7280 10364
rect 7336 10362 7360 10364
rect 7416 10362 7422 10364
rect 7176 10310 7178 10362
rect 7358 10310 7360 10362
rect 7114 10308 7120 10310
rect 7176 10308 7200 10310
rect 7256 10308 7280 10310
rect 7336 10308 7360 10310
rect 7416 10308 7422 10310
rect 7114 10299 7422 10308
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 5920 9586 5948 10066
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5920 9450 5948 9522
rect 6380 9518 6408 10066
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 9110 5856 9318
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5828 8401 5856 9046
rect 6380 9042 6408 9454
rect 6932 9042 6960 9454
rect 7114 9276 7422 9285
rect 7114 9274 7120 9276
rect 7176 9274 7200 9276
rect 7256 9274 7280 9276
rect 7336 9274 7360 9276
rect 7416 9274 7422 9276
rect 7176 9222 7178 9274
rect 7358 9222 7360 9274
rect 7114 9220 7120 9222
rect 7176 9220 7200 9222
rect 7256 9220 7280 9222
rect 7336 9220 7360 9222
rect 7416 9220 7422 9222
rect 7114 9211 7422 9220
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 5908 8424 5960 8430
rect 5814 8392 5870 8401
rect 5908 8366 5960 8372
rect 5814 8327 5870 8336
rect 5920 8090 5948 8366
rect 6104 8362 6132 8910
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 6104 8022 6132 8298
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5828 6866 5856 7142
rect 5920 7002 5948 7210
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 6012 6866 6040 7686
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6012 6390 6040 6802
rect 6288 6474 6316 8774
rect 6380 8498 6408 8978
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 7024 8634 7052 8842
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6092 6452 6144 6458
rect 6288 6446 6408 6474
rect 6656 6458 6684 8502
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7114 8188 7422 8197
rect 7114 8186 7120 8188
rect 7176 8186 7200 8188
rect 7256 8186 7280 8188
rect 7336 8186 7360 8188
rect 7416 8186 7422 8188
rect 7176 8134 7178 8186
rect 7358 8134 7360 8186
rect 7114 8132 7120 8134
rect 7176 8132 7200 8134
rect 7256 8132 7280 8134
rect 7336 8132 7360 8134
rect 7416 8132 7422 8134
rect 7114 8123 7422 8132
rect 7484 8090 7512 8366
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 6932 7546 6960 8026
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7208 7546 7236 7822
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6840 6662 6868 7278
rect 7114 7100 7422 7109
rect 7114 7098 7120 7100
rect 7176 7098 7200 7100
rect 7256 7098 7280 7100
rect 7336 7098 7360 7100
rect 7416 7098 7422 7100
rect 7176 7046 7178 7098
rect 7358 7046 7360 7098
rect 7114 7044 7120 7046
rect 7176 7044 7200 7046
rect 7256 7044 7280 7046
rect 7336 7044 7360 7046
rect 7416 7044 7422 7046
rect 7114 7035 7422 7044
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6092 6394 6144 6400
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5828 5166 5856 5510
rect 5920 5370 5948 6190
rect 6012 5914 6040 6326
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6104 5778 6132 6394
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5846 6224 6054
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6288 5574 6316 6326
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 6288 4690 6316 5510
rect 6380 5302 6408 6446
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6656 5794 6684 6394
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6748 5914 6776 6122
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6656 5766 6776 5794
rect 6642 5672 6698 5681
rect 6642 5607 6644 5616
rect 6696 5607 6698 5616
rect 6644 5578 6696 5584
rect 6656 5370 6684 5578
rect 6748 5574 6776 5766
rect 6840 5710 6868 6598
rect 7116 6458 7144 6734
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7576 6254 7604 6394
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 6932 5846 6960 6190
rect 7576 6066 7604 6190
rect 7484 6038 7604 6066
rect 7114 6012 7422 6021
rect 7114 6010 7120 6012
rect 7176 6010 7200 6012
rect 7256 6010 7280 6012
rect 7336 6010 7360 6012
rect 7416 6010 7422 6012
rect 7176 5958 7178 6010
rect 7358 5958 7360 6010
rect 7114 5956 7120 5958
rect 7176 5956 7200 5958
rect 7256 5956 7280 5958
rect 7336 5956 7360 5958
rect 7416 5956 7422 5958
rect 7114 5947 7422 5956
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6380 4690 6408 5238
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6368 4684 6420 4690
rect 6420 4644 6500 4672
rect 6368 4626 6420 4632
rect 6288 3738 6316 4626
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6380 3194 6408 4014
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6472 3126 6500 4644
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6564 4146 6592 4558
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6564 3602 6592 4082
rect 6840 4010 6868 5646
rect 7392 5370 7420 5714
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7114 4924 7422 4933
rect 7114 4922 7120 4924
rect 7176 4922 7200 4924
rect 7256 4922 7280 4924
rect 7336 4922 7360 4924
rect 7416 4922 7422 4924
rect 7176 4870 7178 4922
rect 7358 4870 7360 4922
rect 7114 4868 7120 4870
rect 7176 4868 7200 4870
rect 7256 4868 7280 4870
rect 7336 4868 7360 4870
rect 7416 4868 7422 4870
rect 7114 4859 7422 4868
rect 7484 4690 7512 6038
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7576 4826 7604 5102
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6840 3534 6868 3946
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 7024 3652 7052 3878
rect 7114 3836 7422 3845
rect 7114 3834 7120 3836
rect 7176 3834 7200 3836
rect 7256 3834 7280 3836
rect 7336 3834 7360 3836
rect 7416 3834 7422 3836
rect 7176 3782 7178 3834
rect 7358 3782 7360 3834
rect 7114 3780 7120 3782
rect 7176 3780 7200 3782
rect 7256 3780 7280 3782
rect 7336 3780 7360 3782
rect 7416 3780 7422 3782
rect 7114 3771 7422 3780
rect 7104 3664 7156 3670
rect 7024 3624 7104 3652
rect 7104 3606 7156 3612
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6460 3120 6512 3126
rect 6460 3062 6512 3068
rect 6840 3058 6868 3470
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 7114 2748 7422 2757
rect 7114 2746 7120 2748
rect 7176 2746 7200 2748
rect 7256 2746 7280 2748
rect 7336 2746 7360 2748
rect 7416 2746 7422 2748
rect 7176 2694 7178 2746
rect 7358 2694 7360 2746
rect 7114 2692 7120 2694
rect 7176 2692 7200 2694
rect 7256 2692 7280 2694
rect 7336 2692 7360 2694
rect 7416 2692 7422 2694
rect 7114 2683 7422 2692
rect 7484 2514 7512 4014
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7576 3670 7604 3878
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7576 2650 7604 2858
rect 7668 2774 7696 12038
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7760 10810 7788 11630
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7852 10690 7880 12242
rect 8036 11898 8064 12242
rect 8956 12238 8984 12310
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7944 10742 7972 11766
rect 8036 11558 8064 11834
rect 8220 11778 8248 12106
rect 8312 11898 8340 12174
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8220 11750 8340 11778
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8128 11354 8156 11630
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 8220 11354 8248 11562
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8312 11234 8340 11750
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 11286 8432 11494
rect 8128 11206 8340 11234
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 7760 10662 7880 10690
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 7760 9654 7788 10662
rect 8128 10606 8156 11206
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10742 8432 10950
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8956 10606 8984 12174
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9140 11286 9168 11494
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 7852 10266 7880 10542
rect 7932 10532 7984 10538
rect 7984 10492 8064 10520
rect 7932 10474 7984 10480
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 8036 9586 8064 10492
rect 8128 9654 8156 10542
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8220 9722 8248 10066
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7838 9480 7894 9489
rect 7838 9415 7894 9424
rect 7852 9042 7880 9415
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 8036 8974 8064 9522
rect 8128 9042 8156 9590
rect 8312 9042 8340 10542
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 10266 9168 10406
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8404 9518 8432 9862
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8588 9518 8616 9590
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8496 9042 8524 9318
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8128 8362 8156 8774
rect 8220 8430 8248 8774
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8588 8090 8616 9454
rect 8772 9178 8800 9454
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 9140 9110 9168 9318
rect 9232 9110 9260 9454
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9220 9104 9272 9110
rect 9220 9046 9272 9052
rect 9324 8906 9352 15914
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9600 14958 9628 15438
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9416 13870 9444 14554
rect 9600 14414 9628 14894
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9508 13870 9536 14010
rect 9586 13968 9642 13977
rect 9586 13903 9588 13912
rect 9640 13903 9642 13912
rect 9588 13874 9640 13880
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9416 12850 9444 13262
rect 9508 12866 9536 13806
rect 9692 13462 9720 16050
rect 10060 15706 10088 16390
rect 10244 16114 10272 16662
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11242 16552 11298 16561
rect 11242 16487 11298 16496
rect 10472 16348 10780 16357
rect 10472 16346 10478 16348
rect 10534 16346 10558 16348
rect 10614 16346 10638 16348
rect 10694 16346 10718 16348
rect 10774 16346 10780 16348
rect 10534 16294 10536 16346
rect 10716 16294 10718 16346
rect 10472 16292 10478 16294
rect 10534 16292 10558 16294
rect 10614 16292 10638 16294
rect 10694 16292 10718 16294
rect 10774 16292 10780 16294
rect 10472 16283 10780 16292
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10324 15972 10376 15978
rect 10324 15914 10376 15920
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10060 14958 10088 15642
rect 10336 15162 10364 15914
rect 11256 15502 11284 16487
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10472 15260 10780 15269
rect 10472 15258 10478 15260
rect 10534 15258 10558 15260
rect 10614 15258 10638 15260
rect 10694 15258 10718 15260
rect 10774 15258 10780 15260
rect 10534 15206 10536 15258
rect 10716 15206 10718 15258
rect 10472 15204 10478 15206
rect 10534 15204 10558 15206
rect 10614 15204 10638 15206
rect 10694 15204 10718 15206
rect 10774 15204 10780 15206
rect 10472 15195 10780 15204
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10980 14958 11008 15370
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11164 14958 11192 15302
rect 10048 14952 10100 14958
rect 9968 14912 10048 14940
rect 9968 14618 9996 14912
rect 10048 14894 10100 14900
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 9404 12844 9456 12850
rect 9508 12838 9628 12866
rect 9404 12786 9456 12792
rect 9600 12782 9628 12838
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9692 12374 9720 13398
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9876 11694 9904 13466
rect 9968 13462 9996 13942
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9968 12782 9996 13398
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9968 12170 9996 12582
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9416 11082 9444 11290
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 7944 6458 7972 6870
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7760 5030 7788 6054
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 4672 7788 4966
rect 7840 4684 7892 4690
rect 7760 4644 7840 4672
rect 7840 4626 7892 4632
rect 7944 4146 7972 6394
rect 8128 6361 8156 6802
rect 8114 6352 8170 6361
rect 8312 6322 8340 7958
rect 8588 6866 8616 8026
rect 8850 7984 8906 7993
rect 8850 7919 8852 7928
rect 8904 7919 8906 7928
rect 9404 7948 9456 7954
rect 8852 7890 8904 7896
rect 9404 7890 9456 7896
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8772 7342 8800 7822
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8680 7002 8708 7278
rect 8864 7002 8892 7890
rect 9416 7410 9444 7890
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8114 6287 8170 6296
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 8036 5166 8064 5782
rect 8404 5370 8432 6054
rect 8588 5778 8616 6054
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8680 5370 8708 6190
rect 8864 5914 8892 6258
rect 9048 6186 9076 6802
rect 9036 6180 9088 6186
rect 9036 6122 9088 6128
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8864 5234 8892 5850
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8956 5574 8984 5714
rect 9048 5574 9076 6122
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 9048 5166 9076 5510
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 8036 4554 8064 5102
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8312 4690 8340 4762
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 7760 3398 7788 3946
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7760 2922 7788 3334
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7668 2746 7880 2774
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 7114 1660 7422 1669
rect 7114 1658 7120 1660
rect 7176 1658 7200 1660
rect 7256 1658 7280 1660
rect 7336 1658 7360 1660
rect 7416 1658 7422 1660
rect 7176 1606 7178 1658
rect 7358 1606 7360 1658
rect 7114 1604 7120 1606
rect 7176 1604 7200 1606
rect 7256 1604 7280 1606
rect 7336 1604 7360 1606
rect 7416 1604 7422 1606
rect 7114 1595 7422 1604
rect 7114 572 7422 581
rect 7114 570 7120 572
rect 7176 570 7200 572
rect 7256 570 7280 572
rect 7336 570 7360 572
rect 7416 570 7422 572
rect 7176 518 7178 570
rect 7358 518 7360 570
rect 7114 516 7120 518
rect 7176 516 7200 518
rect 7256 516 7280 518
rect 7336 516 7360 518
rect 7416 516 7422 518
rect 7114 507 7422 516
rect 6012 462 6132 490
rect 6012 354 6040 462
rect 6104 400 6132 462
rect 7852 400 7880 2746
rect 7944 2514 7972 3878
rect 8128 2854 8156 4150
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8220 3602 8248 3878
rect 8312 3738 8340 4014
rect 8404 4010 8432 5034
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8588 4282 8616 4422
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8680 4026 8708 4422
rect 9048 4282 9076 4626
rect 9128 4548 9180 4554
rect 9128 4490 9180 4496
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 9140 4078 9168 4490
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 4078 9352 4422
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8588 3998 8708 4026
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8220 3126 8248 3538
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8404 1562 8432 3946
rect 8588 3942 8616 3998
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8588 3194 8616 3878
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8680 3194 8708 3606
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 9140 2922 9168 4014
rect 9128 2916 9180 2922
rect 9128 2858 9180 2864
rect 9508 2774 9536 11494
rect 9692 11393 9720 11630
rect 9678 11384 9734 11393
rect 9734 11342 9812 11370
rect 9678 11319 9734 11328
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 10470 9720 11018
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9784 9654 9812 11342
rect 10060 11336 10088 13874
rect 10152 13802 10180 14486
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10244 13870 10272 14350
rect 10336 13938 10364 14554
rect 10472 14172 10780 14181
rect 10472 14170 10478 14172
rect 10534 14170 10558 14172
rect 10614 14170 10638 14172
rect 10694 14170 10718 14172
rect 10774 14170 10780 14172
rect 10534 14118 10536 14170
rect 10716 14118 10718 14170
rect 10472 14116 10478 14118
rect 10534 14116 10558 14118
rect 10614 14116 10638 14118
rect 10694 14116 10718 14118
rect 10774 14116 10780 14118
rect 10472 14107 10780 14116
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10152 13530 10180 13738
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10244 13394 10272 13806
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10244 12646 10272 13330
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10472 13084 10780 13093
rect 10472 13082 10478 13084
rect 10534 13082 10558 13084
rect 10614 13082 10638 13084
rect 10694 13082 10718 13084
rect 10774 13082 10780 13084
rect 10534 13030 10536 13082
rect 10716 13030 10718 13082
rect 10472 13028 10478 13030
rect 10534 13028 10558 13030
rect 10614 13028 10638 13030
rect 10694 13028 10718 13030
rect 10774 13028 10780 13030
rect 10472 13019 10780 13028
rect 10506 12880 10562 12889
rect 10506 12815 10562 12824
rect 10520 12782 10548 12815
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10152 12102 10180 12582
rect 10874 12472 10930 12481
rect 10980 12442 11008 13262
rect 11072 12986 11100 13330
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10874 12407 10930 12416
rect 10968 12436 11020 12442
rect 10888 12306 10916 12407
rect 10968 12378 11020 12384
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10888 12209 10916 12242
rect 10874 12200 10930 12209
rect 10874 12135 10930 12144
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10472 11996 10780 12005
rect 10472 11994 10478 11996
rect 10534 11994 10558 11996
rect 10614 11994 10638 11996
rect 10694 11994 10718 11996
rect 10774 11994 10780 11996
rect 10534 11942 10536 11994
rect 10716 11942 10718 11994
rect 10472 11940 10478 11942
rect 10534 11940 10558 11942
rect 10614 11940 10638 11942
rect 10694 11940 10718 11942
rect 10774 11940 10780 11942
rect 10472 11931 10780 11940
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10336 11694 10364 11834
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10060 11308 10180 11336
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9876 10810 9904 11086
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 10060 10130 10088 11154
rect 10152 10674 10180 11308
rect 10980 11150 11008 12378
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11072 11529 11100 11630
rect 11152 11552 11204 11558
rect 11058 11520 11114 11529
rect 11152 11494 11204 11500
rect 11058 11455 11114 11464
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10472 10908 10780 10917
rect 10472 10906 10478 10908
rect 10534 10906 10558 10908
rect 10614 10906 10638 10908
rect 10694 10906 10718 10908
rect 10774 10906 10780 10908
rect 10534 10854 10536 10906
rect 10716 10854 10718 10906
rect 10472 10852 10478 10854
rect 10534 10852 10558 10854
rect 10614 10852 10638 10854
rect 10694 10852 10718 10854
rect 10774 10852 10780 10854
rect 10472 10843 10780 10852
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 11072 10606 11100 11154
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 11072 10130 11100 10542
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9600 9178 9628 9454
rect 10060 9450 10088 10066
rect 10472 9820 10780 9829
rect 10472 9818 10478 9820
rect 10534 9818 10558 9820
rect 10614 9818 10638 9820
rect 10694 9818 10718 9820
rect 10774 9818 10780 9820
rect 10534 9766 10536 9818
rect 10716 9766 10718 9818
rect 10472 9764 10478 9766
rect 10534 9764 10558 9766
rect 10614 9764 10638 9766
rect 10694 9764 10718 9766
rect 10774 9764 10780 9766
rect 10472 9755 10780 9764
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9692 9178 9720 9318
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9876 9110 9904 9318
rect 10060 9110 10088 9386
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9600 8090 9628 8434
rect 9692 8430 9720 8910
rect 10060 8537 10088 9046
rect 10506 8936 10562 8945
rect 10140 8900 10192 8906
rect 10506 8871 10508 8880
rect 10140 8842 10192 8848
rect 10560 8871 10562 8880
rect 10508 8842 10560 8848
rect 10046 8528 10102 8537
rect 10046 8463 10102 8472
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9692 7342 9720 8366
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9692 7002 9720 7278
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9692 6118 9720 6938
rect 10060 6866 10088 7686
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 9862 6352 9918 6361
rect 9862 6287 9918 6296
rect 9876 6254 9904 6287
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9600 4622 9628 6054
rect 9692 5846 9720 6054
rect 10152 5914 10180 8842
rect 10472 8732 10780 8741
rect 10472 8730 10478 8732
rect 10534 8730 10558 8732
rect 10614 8730 10638 8732
rect 10694 8730 10718 8732
rect 10774 8730 10780 8732
rect 10534 8678 10536 8730
rect 10716 8678 10718 8730
rect 10472 8676 10478 8678
rect 10534 8676 10558 8678
rect 10614 8676 10638 8678
rect 10694 8676 10718 8678
rect 10774 8676 10780 8678
rect 10472 8667 10780 8676
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10472 7644 10780 7653
rect 10472 7642 10478 7644
rect 10534 7642 10558 7644
rect 10614 7642 10638 7644
rect 10694 7642 10718 7644
rect 10774 7642 10780 7644
rect 10534 7590 10536 7642
rect 10716 7590 10718 7642
rect 10472 7588 10478 7590
rect 10534 7588 10558 7590
rect 10614 7588 10638 7590
rect 10694 7588 10718 7590
rect 10774 7588 10780 7590
rect 10472 7579 10780 7588
rect 10888 7002 10916 7958
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10472 6556 10780 6565
rect 10472 6554 10478 6556
rect 10534 6554 10558 6556
rect 10614 6554 10638 6556
rect 10694 6554 10718 6556
rect 10774 6554 10780 6556
rect 10534 6502 10536 6554
rect 10716 6502 10718 6554
rect 10472 6500 10478 6502
rect 10534 6500 10558 6502
rect 10614 6500 10638 6502
rect 10694 6500 10718 6502
rect 10774 6500 10780 6502
rect 10472 6491 10780 6500
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9956 4752 10008 4758
rect 9956 4694 10008 4700
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9968 4282 9996 4694
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9968 3602 9996 4218
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9692 2990 9720 3402
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9862 2952 9918 2961
rect 9862 2887 9918 2896
rect 9508 2746 9628 2774
rect 9220 1760 9272 1766
rect 9220 1702 9272 1708
rect 8392 1556 8444 1562
rect 8392 1498 8444 1504
rect 9232 1494 9260 1702
rect 9220 1488 9272 1494
rect 9220 1430 9272 1436
rect 9600 400 9628 2746
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 2106 9720 2246
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 9876 1834 9904 2887
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10060 2514 10088 2790
rect 10152 2774 10180 5850
rect 10980 5778 11008 6598
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10472 5468 10780 5477
rect 10472 5466 10478 5468
rect 10534 5466 10558 5468
rect 10614 5466 10638 5468
rect 10694 5466 10718 5468
rect 10774 5466 10780 5468
rect 10534 5414 10536 5466
rect 10716 5414 10718 5466
rect 10472 5412 10478 5414
rect 10534 5412 10558 5414
rect 10614 5412 10638 5414
rect 10694 5412 10718 5414
rect 10774 5412 10780 5414
rect 10472 5403 10780 5412
rect 11164 5302 11192 11494
rect 11256 11218 11284 15438
rect 11348 14074 11376 16594
rect 11612 16448 11664 16454
rect 11612 16390 11664 16396
rect 11624 16046 11652 16390
rect 11716 16250 11744 16594
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11980 16108 12032 16114
rect 11900 16068 11980 16096
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11520 15972 11572 15978
rect 11520 15914 11572 15920
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11440 14414 11468 14826
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11532 14006 11560 15914
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 11428 13728 11480 13734
rect 11428 13670 11480 13676
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11348 12782 11376 13126
rect 11440 12782 11468 13670
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11348 11694 11376 12242
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11440 11626 11468 11834
rect 11624 11694 11652 15982
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11716 14958 11744 15030
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11716 12782 11744 14894
rect 11808 14414 11836 15506
rect 11900 15201 11928 16068
rect 11980 16050 12032 16056
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11992 15570 12020 15914
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 11886 15192 11942 15201
rect 11886 15127 11942 15136
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11808 13870 11836 14350
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11900 13462 11928 15127
rect 12084 14958 12112 17070
rect 12164 15972 12216 15978
rect 12164 15914 12216 15920
rect 12176 15502 12204 15914
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11716 11801 11744 12718
rect 12176 12434 12204 15438
rect 12268 14958 12296 15846
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12360 14618 12388 17070
rect 12728 15162 12756 17070
rect 13648 16794 13676 17600
rect 13830 16892 14138 16901
rect 13830 16890 13836 16892
rect 13892 16890 13916 16892
rect 13972 16890 13996 16892
rect 14052 16890 14076 16892
rect 14132 16890 14138 16892
rect 13892 16838 13894 16890
rect 14074 16838 14076 16890
rect 13830 16836 13836 16838
rect 13892 16836 13916 16838
rect 13972 16836 13996 16838
rect 14052 16836 14076 16838
rect 14132 16836 14138 16838
rect 13830 16827 14138 16836
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 14096 16788 14148 16794
rect 14200 16776 14228 17734
rect 14278 17600 14334 17734
rect 14660 17734 14978 17762
rect 14148 16748 14228 16776
rect 14096 16730 14148 16736
rect 14660 16726 14688 17734
rect 14922 17600 14978 17734
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 14648 16720 14700 16726
rect 14648 16662 14700 16668
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12820 14958 12848 15506
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12452 14278 12480 14894
rect 12440 14272 12492 14278
rect 12492 14220 12572 14226
rect 12440 14214 12572 14220
rect 12452 14198 12572 14214
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12268 12753 12296 13670
rect 12452 13530 12480 13670
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12360 12850 12388 13194
rect 12452 12986 12480 13330
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12254 12744 12310 12753
rect 12254 12679 12310 12688
rect 12084 12406 12204 12434
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11992 11898 12020 12106
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11702 11792 11758 11801
rect 11702 11727 11758 11736
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11610 11520 11666 11529
rect 11610 11455 11666 11464
rect 11624 11257 11652 11455
rect 11900 11286 11928 11698
rect 11888 11280 11940 11286
rect 11610 11248 11666 11257
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11428 11212 11480 11218
rect 11888 11222 11940 11228
rect 11610 11183 11666 11192
rect 11704 11212 11756 11218
rect 11428 11154 11480 11160
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11256 10130 11284 10746
rect 11440 10520 11468 11154
rect 11520 10532 11572 10538
rect 11348 10492 11520 10520
rect 11348 10130 11376 10492
rect 11520 10474 11572 10480
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11348 9450 11376 10066
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11440 9518 11468 9998
rect 11428 9512 11480 9518
rect 11624 9489 11652 11183
rect 11704 11154 11756 11160
rect 11716 10606 11744 11154
rect 11704 10600 11756 10606
rect 11980 10600 12032 10606
rect 11704 10542 11756 10548
rect 11978 10568 11980 10577
rect 12032 10568 12034 10577
rect 11716 10130 11744 10542
rect 11978 10503 12034 10512
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11888 10124 11940 10130
rect 11992 10112 12020 10503
rect 11940 10084 12020 10112
rect 11888 10066 11940 10072
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11808 9602 11836 9930
rect 12084 9761 12112 12406
rect 12452 12170 12480 12922
rect 12544 12889 12572 14198
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12636 13433 12664 14010
rect 13004 13938 13032 15098
rect 13096 15008 13124 16050
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13188 15706 13216 15846
rect 13556 15706 13584 16390
rect 13924 16250 13952 16594
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13740 15094 13768 15846
rect 13830 15804 14138 15813
rect 13830 15802 13836 15804
rect 13892 15802 13916 15804
rect 13972 15802 13996 15804
rect 14052 15802 14076 15804
rect 14132 15802 14138 15804
rect 13892 15750 13894 15802
rect 14074 15750 14076 15802
rect 13830 15748 13836 15750
rect 13892 15748 13916 15750
rect 13972 15748 13996 15750
rect 14052 15748 14076 15750
rect 14132 15748 14138 15750
rect 13830 15739 14138 15748
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 14108 15026 14136 15438
rect 13176 15020 13228 15026
rect 13096 14980 13176 15008
rect 13176 14962 13228 14968
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 13188 14414 13216 14962
rect 13832 14906 13860 14962
rect 13740 14878 13860 14906
rect 13910 14920 13966 14929
rect 13740 14414 13768 14878
rect 13910 14855 13912 14864
rect 13964 14855 13966 14864
rect 13912 14826 13964 14832
rect 13830 14716 14138 14725
rect 13830 14714 13836 14716
rect 13892 14714 13916 14716
rect 13972 14714 13996 14716
rect 14052 14714 14076 14716
rect 14132 14714 14138 14716
rect 13892 14662 13894 14714
rect 14074 14662 14076 14714
rect 13830 14660 13836 14662
rect 13892 14660 13916 14662
rect 13972 14660 13996 14662
rect 14052 14660 14076 14662
rect 14132 14660 14138 14662
rect 13830 14651 14138 14660
rect 14200 14618 14228 16594
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14476 15706 14504 15846
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14936 15502 14964 17138
rect 15488 17066 15516 17682
rect 15566 17600 15622 18000
rect 16210 17600 16266 18000
rect 16672 17604 16724 17610
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15120 16794 15148 16934
rect 15580 16794 15608 17600
rect 16854 17600 16910 18000
rect 17498 17600 17554 18000
rect 18142 17762 18198 18000
rect 18142 17734 18276 17762
rect 18142 17600 18198 17734
rect 16672 17546 16724 17552
rect 15936 17264 15988 17270
rect 16120 17264 16172 17270
rect 15988 17224 16120 17252
rect 15936 17206 15988 17212
rect 16120 17206 16172 17212
rect 16684 17134 16712 17546
rect 16868 17202 16896 17600
rect 17512 17524 17540 17600
rect 17512 17496 17632 17524
rect 17188 17436 17496 17445
rect 17188 17434 17194 17436
rect 17250 17434 17274 17436
rect 17330 17434 17354 17436
rect 17410 17434 17434 17436
rect 17490 17434 17496 17436
rect 17250 17382 17252 17434
rect 17432 17382 17434 17434
rect 17188 17380 17194 17382
rect 17250 17380 17274 17382
rect 17330 17380 17354 17382
rect 17410 17380 17434 17382
rect 17490 17380 17496 17382
rect 17188 17371 17496 17380
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 17604 17134 17632 17496
rect 18248 17134 18276 17734
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 16672 17128 16724 17134
rect 17592 17128 17644 17134
rect 16724 17076 17172 17082
rect 16672 17070 17172 17076
rect 17592 17070 17644 17076
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 16684 17054 17172 17070
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15120 16561 15148 16594
rect 15292 16584 15344 16590
rect 15106 16552 15162 16561
rect 15292 16526 15344 16532
rect 15106 16487 15162 16496
rect 15304 16114 15332 16526
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 13176 14408 13228 14414
rect 13544 14408 13596 14414
rect 13228 14368 13308 14396
rect 13176 14350 13228 14356
rect 13280 13938 13308 14368
rect 13544 14350 13596 14356
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 12992 13932 13044 13938
rect 13268 13932 13320 13938
rect 13044 13892 13216 13920
rect 12992 13874 13044 13880
rect 12622 13424 12678 13433
rect 12622 13359 12624 13368
rect 12676 13359 12678 13368
rect 12624 13330 12676 13336
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12530 12880 12586 12889
rect 12530 12815 12532 12824
rect 12584 12815 12586 12824
rect 12532 12786 12584 12792
rect 12728 12782 12756 13126
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12176 10606 12204 10950
rect 12360 10742 12388 11290
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12268 10452 12296 10542
rect 12440 10464 12492 10470
rect 12268 10424 12440 10452
rect 12440 10406 12492 10412
rect 12452 10198 12480 10406
rect 12440 10192 12492 10198
rect 12440 10134 12492 10140
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12070 9752 12126 9761
rect 12070 9687 12126 9696
rect 11716 9574 11836 9602
rect 11716 9518 11744 9574
rect 11704 9512 11756 9518
rect 11428 9454 11480 9460
rect 11610 9480 11666 9489
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 11440 9330 11468 9454
rect 11704 9454 11756 9460
rect 11610 9415 11666 9424
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11808 9330 11836 9386
rect 11980 9376 12032 9382
rect 11348 9302 11468 9330
rect 11716 9302 11836 9330
rect 11900 9324 11980 9330
rect 11900 9318 12032 9324
rect 11900 9302 12020 9318
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11256 8634 11284 8978
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11348 8294 11376 9302
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11428 8424 11480 8430
rect 11532 8412 11560 9046
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11624 8430 11652 8774
rect 11480 8384 11560 8412
rect 11612 8424 11664 8430
rect 11428 8366 11480 8372
rect 11612 8366 11664 8372
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11348 7954 11376 8230
rect 11518 8120 11574 8129
rect 11518 8055 11574 8064
rect 11532 7954 11560 8055
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11716 7886 11744 9302
rect 11900 9110 11928 9302
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11992 8906 12020 9114
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11888 8424 11940 8430
rect 11992 8412 12020 8842
rect 12084 8430 12112 9687
rect 12268 9518 12296 9862
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12176 9110 12204 9318
rect 12164 9104 12216 9110
rect 12268 9081 12296 9454
rect 12360 9178 12388 9454
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12164 9046 12216 9052
rect 12254 9072 12310 9081
rect 12254 9007 12310 9016
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12176 8498 12204 8910
rect 12268 8498 12296 9007
rect 12544 8838 12572 12174
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12636 10810 12664 11154
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12716 10600 12768 10606
rect 12714 10568 12716 10577
rect 12768 10568 12770 10577
rect 12714 10503 12770 10512
rect 12728 9654 12756 10503
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12346 8664 12402 8673
rect 12346 8599 12402 8608
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 11940 8384 12020 8412
rect 12072 8424 12124 8430
rect 11888 8366 11940 8372
rect 12072 8366 12124 8372
rect 12360 8362 12388 8599
rect 12728 8566 12756 9590
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12820 8673 12848 9318
rect 12912 8974 12940 10406
rect 13004 9178 13032 12582
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12806 8664 12862 8673
rect 12806 8599 12862 8608
rect 12716 8560 12768 8566
rect 12768 8520 12940 8548
rect 12716 8502 12768 8508
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12176 7954 12204 8298
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11612 7812 11664 7818
rect 11612 7754 11664 7760
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11256 5642 11284 6734
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11348 5778 11376 6122
rect 11532 5778 11560 6190
rect 11624 6118 11652 7754
rect 11716 7342 11744 7822
rect 12268 7342 12296 8298
rect 12532 8288 12584 8294
rect 12584 8248 12756 8276
rect 12532 8230 12584 8236
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12360 7546 12388 7890
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12544 7002 12572 8026
rect 12636 7342 12664 8026
rect 12728 7954 12756 8248
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12636 6866 12664 7142
rect 12728 6866 12756 7686
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11808 6118 11836 6258
rect 11900 6254 11928 6802
rect 11992 6390 12020 6802
rect 11980 6384 12032 6390
rect 12032 6332 12112 6338
rect 11980 6326 12112 6332
rect 11992 6310 12112 6326
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11624 5778 11652 6054
rect 11716 5846 11744 6054
rect 11992 5914 12020 6190
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12084 5846 12112 6310
rect 12176 5846 12204 6802
rect 12820 6798 12848 7278
rect 12912 6866 12940 8520
rect 13004 6866 13032 9114
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12268 6322 12296 6598
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12348 6248 12400 6254
rect 12254 6216 12310 6225
rect 12348 6190 12400 6196
rect 12254 6151 12256 6160
rect 12308 6151 12310 6160
rect 12256 6122 12308 6128
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11348 5030 11376 5510
rect 11440 5370 11468 5714
rect 11532 5574 11560 5714
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11348 4486 11376 4966
rect 11532 4554 11560 5510
rect 11624 5166 11652 5714
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11612 5160 11664 5166
rect 11612 5102 11664 5108
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 10472 4380 10780 4389
rect 10472 4378 10478 4380
rect 10534 4378 10558 4380
rect 10614 4378 10638 4380
rect 10694 4378 10718 4380
rect 10774 4378 10780 4380
rect 10534 4326 10536 4378
rect 10716 4326 10718 4378
rect 10472 4324 10478 4326
rect 10534 4324 10558 4326
rect 10614 4324 10638 4326
rect 10694 4324 10718 4326
rect 10774 4324 10780 4326
rect 10472 4315 10780 4324
rect 10888 4078 10916 4422
rect 11624 4078 11652 5102
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11624 3602 11652 4014
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 10472 3292 10780 3301
rect 10472 3290 10478 3292
rect 10534 3290 10558 3292
rect 10614 3290 10638 3292
rect 10694 3290 10718 3292
rect 10774 3290 10780 3292
rect 10534 3238 10536 3290
rect 10716 3238 10718 3290
rect 10472 3236 10478 3238
rect 10534 3236 10558 3238
rect 10614 3236 10638 3238
rect 10694 3236 10718 3238
rect 10774 3236 10780 3238
rect 10472 3227 10780 3236
rect 11428 2984 11480 2990
rect 11256 2932 11428 2938
rect 11256 2926 11480 2932
rect 11256 2910 11468 2926
rect 10152 2746 10272 2774
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 9864 1828 9916 1834
rect 9864 1770 9916 1776
rect 9876 1562 9904 1770
rect 10060 1562 10088 2450
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10152 1902 10180 2246
rect 10244 1986 10272 2746
rect 11256 2650 11284 2910
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 10324 2372 10376 2378
rect 10324 2314 10376 2320
rect 10336 2088 10364 2314
rect 10472 2204 10780 2213
rect 10472 2202 10478 2204
rect 10534 2202 10558 2204
rect 10614 2202 10638 2204
rect 10694 2202 10718 2204
rect 10774 2202 10780 2204
rect 10534 2150 10536 2202
rect 10716 2150 10718 2202
rect 10472 2148 10478 2150
rect 10534 2148 10558 2150
rect 10614 2148 10638 2150
rect 10694 2148 10718 2150
rect 10774 2148 10780 2150
rect 10472 2139 10780 2148
rect 10980 2106 11008 2382
rect 11072 2106 11100 2450
rect 11348 2446 11376 2790
rect 11440 2514 11468 2910
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 10968 2100 11020 2106
rect 10336 2060 10640 2088
rect 10244 1958 10548 1986
rect 10612 1970 10640 2060
rect 10968 2042 11020 2048
rect 11060 2100 11112 2106
rect 11060 2042 11112 2048
rect 11532 1970 11560 2586
rect 10520 1902 10548 1958
rect 10600 1964 10652 1970
rect 10600 1906 10652 1912
rect 11520 1964 11572 1970
rect 11520 1906 11572 1912
rect 10140 1896 10192 1902
rect 10140 1838 10192 1844
rect 10508 1896 10560 1902
rect 10508 1838 10560 1844
rect 10612 1562 10640 1906
rect 11152 1760 11204 1766
rect 11152 1702 11204 1708
rect 9864 1556 9916 1562
rect 9864 1498 9916 1504
rect 10048 1556 10100 1562
rect 10048 1498 10100 1504
rect 10600 1556 10652 1562
rect 10600 1498 10652 1504
rect 11164 1494 11192 1702
rect 11152 1488 11204 1494
rect 11152 1430 11204 1436
rect 11624 1222 11652 3538
rect 11716 2774 11744 5238
rect 12268 5098 12296 6122
rect 12360 5370 12388 6190
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12452 5098 12480 6666
rect 13004 5166 13032 6802
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11808 3194 11836 4490
rect 12268 4214 12296 5034
rect 13004 4842 13032 5102
rect 12912 4814 13032 4842
rect 12912 4758 12940 4814
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12900 4752 12952 4758
rect 12900 4694 12952 4700
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 12268 2990 12296 3674
rect 12452 3194 12480 4694
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12544 3058 12572 4218
rect 12728 4078 12756 4626
rect 12820 4554 12848 4626
rect 12808 4548 12860 4554
rect 12808 4490 12860 4496
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 11716 2746 11836 2774
rect 11612 1216 11664 1222
rect 11612 1158 11664 1164
rect 10472 1116 10780 1125
rect 10472 1114 10478 1116
rect 10534 1114 10558 1116
rect 10614 1114 10638 1116
rect 10694 1114 10718 1116
rect 10774 1114 10780 1116
rect 10534 1062 10536 1114
rect 10716 1062 10718 1114
rect 10472 1060 10478 1062
rect 10534 1060 10558 1062
rect 10614 1060 10638 1062
rect 10694 1060 10718 1062
rect 10774 1060 10780 1062
rect 10472 1051 10780 1060
rect 11348 462 11468 490
rect 11348 400 11376 462
rect 5736 326 6040 354
rect 6090 0 6146 400
rect 7838 0 7894 400
rect 9586 0 9642 400
rect 11334 0 11390 400
rect 11440 354 11468 462
rect 11808 354 11836 2746
rect 12268 2650 12296 2926
rect 12912 2774 12940 3334
rect 13004 3194 13032 3606
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 12544 2746 12940 2774
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12544 2582 12572 2746
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 13004 2514 13032 2926
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 11992 1766 12020 2382
rect 12268 1884 12296 2450
rect 12348 1896 12400 1902
rect 12268 1856 12348 1884
rect 12348 1838 12400 1844
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 12360 1222 12388 1838
rect 12728 1494 12756 2450
rect 13004 2378 13032 2450
rect 12992 2372 13044 2378
rect 12992 2314 13044 2320
rect 12716 1488 12768 1494
rect 12716 1430 12768 1436
rect 12808 1420 12860 1426
rect 12808 1362 12860 1368
rect 12348 1216 12400 1222
rect 12348 1158 12400 1164
rect 12820 1018 12848 1362
rect 12808 1012 12860 1018
rect 12808 954 12860 960
rect 13096 400 13124 12038
rect 13188 9042 13216 13892
rect 13268 13874 13320 13880
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13464 12986 13492 13466
rect 13556 13462 13584 14350
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13280 12102 13308 12174
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13372 11014 13400 11630
rect 13464 11626 13492 12582
rect 13452 11620 13504 11626
rect 13452 11562 13504 11568
rect 13556 11354 13584 13398
rect 13740 13326 13768 14350
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 13830 13628 14138 13637
rect 13830 13626 13836 13628
rect 13892 13626 13916 13628
rect 13972 13626 13996 13628
rect 14052 13626 14076 13628
rect 14132 13626 14138 13628
rect 13892 13574 13894 13626
rect 14074 13574 14076 13626
rect 13830 13572 13836 13574
rect 13892 13572 13916 13574
rect 13972 13572 13996 13574
rect 14052 13572 14076 13574
rect 14132 13572 14138 13574
rect 13830 13563 14138 13572
rect 14200 13530 14228 13670
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 14384 12714 14412 13670
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 13830 12540 14138 12549
rect 13830 12538 13836 12540
rect 13892 12538 13916 12540
rect 13972 12538 13996 12540
rect 14052 12538 14076 12540
rect 14132 12538 14138 12540
rect 13892 12486 13894 12538
rect 14074 12486 14076 12538
rect 13830 12484 13836 12486
rect 13892 12484 13916 12486
rect 13972 12484 13996 12486
rect 14052 12484 14076 12486
rect 14132 12484 14138 12486
rect 13830 12475 14138 12484
rect 14200 12374 14228 12582
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14292 11694 14320 12242
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 13830 11452 14138 11461
rect 13830 11450 13836 11452
rect 13892 11450 13916 11452
rect 13972 11450 13996 11452
rect 14052 11450 14076 11452
rect 14132 11450 14138 11452
rect 13892 11398 13894 11450
rect 14074 11398 14076 11450
rect 13830 11396 13836 11398
rect 13892 11396 13916 11398
rect 13972 11396 13996 11398
rect 14052 11396 14076 11398
rect 14132 11396 14138 11398
rect 13634 11384 13690 11393
rect 13830 11387 14138 11396
rect 13544 11348 13596 11354
rect 13820 11348 13872 11354
rect 13690 11328 13820 11336
rect 13634 11319 13820 11328
rect 13648 11308 13820 11319
rect 13544 11290 13596 11296
rect 13820 11290 13872 11296
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13830 10364 14138 10373
rect 13830 10362 13836 10364
rect 13892 10362 13916 10364
rect 13972 10362 13996 10364
rect 14052 10362 14076 10364
rect 14132 10362 14138 10364
rect 13892 10310 13894 10362
rect 14074 10310 14076 10362
rect 13830 10308 13836 10310
rect 13892 10308 13916 10310
rect 13972 10308 13996 10310
rect 14052 10308 14076 10310
rect 14132 10308 14138 10310
rect 13830 10299 14138 10308
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 14002 9616 14058 9625
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13188 7342 13216 8978
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13280 8294 13308 8910
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13176 7200 13228 7206
rect 13280 7188 13308 8230
rect 13228 7160 13308 7188
rect 13176 7142 13228 7148
rect 13372 6458 13400 9454
rect 13464 9178 13492 9522
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13556 9042 13584 9590
rect 14002 9551 14004 9560
rect 14056 9551 14058 9560
rect 14004 9522 14056 9528
rect 13830 9276 14138 9285
rect 13830 9274 13836 9276
rect 13892 9274 13916 9276
rect 13972 9274 13996 9276
rect 14052 9274 14076 9276
rect 14132 9274 14138 9276
rect 13892 9222 13894 9274
rect 14074 9222 14076 9274
rect 13830 9220 13836 9222
rect 13892 9220 13916 9222
rect 13972 9220 13996 9222
rect 14052 9220 14076 9222
rect 14132 9220 14138 9222
rect 13830 9211 14138 9220
rect 14004 9104 14056 9110
rect 13726 9072 13782 9081
rect 13544 9036 13596 9042
rect 14004 9046 14056 9052
rect 13726 9007 13782 9016
rect 13544 8978 13596 8984
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13464 8129 13492 8366
rect 13556 8294 13584 8978
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13648 8129 13676 8570
rect 13450 8120 13506 8129
rect 13450 8055 13506 8064
rect 13634 8120 13690 8129
rect 13634 8055 13690 8064
rect 13740 8072 13768 9007
rect 13818 8664 13874 8673
rect 13818 8599 13874 8608
rect 13832 8362 13860 8599
rect 13910 8528 13966 8537
rect 13910 8463 13966 8472
rect 13924 8362 13952 8463
rect 14016 8362 14044 9046
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13830 8188 14138 8197
rect 13830 8186 13836 8188
rect 13892 8186 13916 8188
rect 13972 8186 13996 8188
rect 14052 8186 14076 8188
rect 14132 8186 14138 8188
rect 13892 8134 13894 8186
rect 14074 8134 14076 8186
rect 13830 8132 13836 8134
rect 13892 8132 13916 8134
rect 13972 8132 13996 8134
rect 14052 8132 14076 8134
rect 14132 8132 14138 8134
rect 13830 8123 14138 8132
rect 13740 8044 14044 8072
rect 14016 7954 14044 8044
rect 13728 7948 13780 7954
rect 13648 7908 13728 7936
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13556 7410 13584 7686
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13648 7274 13676 7908
rect 13728 7890 13780 7896
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 13924 7478 13952 7890
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 13648 6934 13676 7210
rect 13830 7100 14138 7109
rect 13830 7098 13836 7100
rect 13892 7098 13916 7100
rect 13972 7098 13996 7100
rect 14052 7098 14076 7100
rect 14132 7098 14138 7100
rect 13892 7046 13894 7098
rect 14074 7046 14076 7098
rect 13830 7044 13836 7046
rect 13892 7044 13916 7046
rect 13972 7044 13996 7046
rect 14052 7044 14076 7046
rect 14132 7044 14138 7046
rect 13830 7035 14138 7044
rect 13636 6928 13688 6934
rect 13636 6870 13688 6876
rect 14096 6860 14148 6866
rect 14200 6848 14228 11494
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10606 14320 10950
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14292 10198 14320 10542
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 14292 9042 14320 10134
rect 14384 10130 14412 12650
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14476 9994 14504 14962
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14568 12442 14596 13262
rect 14660 13138 14688 14214
rect 14752 14074 14780 14350
rect 14936 14074 14964 15438
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14660 13110 14780 13138
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14568 11694 14596 12378
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14660 11694 14688 12310
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 14752 9110 14780 13110
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 14936 12306 14964 12378
rect 15028 12374 15056 15914
rect 15304 15638 15332 16050
rect 15292 15632 15344 15638
rect 15292 15574 15344 15580
rect 15672 15570 15700 16594
rect 15764 16114 15792 16934
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15568 15088 15620 15094
rect 15568 15030 15620 15036
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 15120 13938 15148 14350
rect 15212 14006 15240 14418
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15120 12782 15148 13262
rect 15212 12918 15240 13330
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15120 12442 15148 12718
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15016 12368 15068 12374
rect 15016 12310 15068 12316
rect 15212 12306 15240 12854
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 14844 11626 14872 12242
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 14832 11620 14884 11626
rect 14832 11562 14884 11568
rect 14740 9104 14792 9110
rect 14740 9046 14792 9052
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14384 8022 14412 8230
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 14568 7954 14596 8230
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14844 7342 14872 7686
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14148 6820 14228 6848
rect 14096 6802 14148 6808
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13372 5914 13400 6394
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 13188 4282 13216 4626
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13188 3670 13216 3878
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13188 1766 13216 2790
rect 13280 2582 13308 3470
rect 13372 3058 13400 5850
rect 13556 5574 13584 6734
rect 13830 6012 14138 6021
rect 13830 6010 13836 6012
rect 13892 6010 13916 6012
rect 13972 6010 13996 6012
rect 14052 6010 14076 6012
rect 14132 6010 14138 6012
rect 13892 5958 13894 6010
rect 14074 5958 14076 6010
rect 13830 5956 13836 5958
rect 13892 5956 13916 5958
rect 13972 5956 13996 5958
rect 14052 5956 14076 5958
rect 14132 5956 14138 5958
rect 13830 5947 14138 5956
rect 14200 5828 14228 6820
rect 14384 6254 14412 7142
rect 14568 6798 14596 7278
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14108 5800 14228 5828
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13648 5370 13676 5646
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 14108 5234 14136 5800
rect 14384 5778 14412 6190
rect 14568 6186 14596 6734
rect 14844 6458 14872 6802
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14372 5772 14424 5778
rect 14200 5732 14372 5760
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 13648 4690 13676 5170
rect 13830 4924 14138 4933
rect 13830 4922 13836 4924
rect 13892 4922 13916 4924
rect 13972 4922 13996 4924
rect 14052 4922 14076 4924
rect 14132 4922 14138 4924
rect 13892 4870 13894 4922
rect 14074 4870 14076 4922
rect 13830 4868 13836 4870
rect 13892 4868 13916 4870
rect 13972 4868 13996 4870
rect 14052 4868 14076 4870
rect 14132 4868 14138 4870
rect 13830 4859 14138 4868
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 14004 4684 14056 4690
rect 14200 4672 14228 5732
rect 14372 5714 14424 5720
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14476 5681 14504 5714
rect 14462 5672 14518 5681
rect 14462 5607 14518 5616
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14476 4690 14504 4966
rect 14056 4644 14228 4672
rect 14004 4626 14056 4632
rect 13648 4554 13676 4626
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 13556 3602 13584 4150
rect 14200 4078 14228 4644
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14476 4078 14504 4626
rect 14568 4622 14596 6122
rect 14660 5778 14688 6190
rect 14936 5914 14964 6190
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14660 5030 14688 5714
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14844 4282 14872 4626
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 15028 4162 15056 12106
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15198 9752 15254 9761
rect 15198 9687 15254 9696
rect 15212 9654 15240 9687
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15212 5778 15240 6598
rect 15304 5778 15332 6938
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15396 5778 15424 6054
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 14844 4134 15056 4162
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 13452 3596 13504 3602
rect 13452 3538 13504 3544
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13464 3126 13492 3538
rect 13648 3398 13676 4014
rect 13830 3836 14138 3845
rect 13830 3834 13836 3836
rect 13892 3834 13916 3836
rect 13972 3834 13996 3836
rect 14052 3834 14076 3836
rect 14132 3834 14138 3836
rect 13892 3782 13894 3834
rect 14074 3782 14076 3834
rect 13830 3780 13836 3782
rect 13892 3780 13916 3782
rect 13972 3780 13996 3782
rect 14052 3780 14076 3782
rect 14132 3780 14138 3782
rect 13830 3771 14138 3780
rect 14200 3602 14228 4014
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13358 2952 13414 2961
rect 13358 2887 13414 2896
rect 13372 2650 13400 2887
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13268 2576 13320 2582
rect 13464 2553 13492 3062
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13740 2564 13768 2790
rect 13830 2748 14138 2757
rect 13830 2746 13836 2748
rect 13892 2746 13916 2748
rect 13972 2746 13996 2748
rect 14052 2746 14076 2748
rect 14132 2746 14138 2748
rect 13892 2694 13894 2746
rect 14074 2694 14076 2746
rect 13830 2692 13836 2694
rect 13892 2692 13916 2694
rect 13972 2692 13996 2694
rect 14052 2692 14076 2694
rect 14132 2692 14138 2694
rect 13830 2683 14138 2692
rect 14200 2650 14228 3130
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 13912 2576 13964 2582
rect 13268 2518 13320 2524
rect 13450 2544 13506 2553
rect 13280 2310 13308 2518
rect 13740 2536 13912 2564
rect 14280 2576 14332 2582
rect 13912 2518 13964 2524
rect 14094 2544 14150 2553
rect 13450 2479 13506 2488
rect 14280 2518 14332 2524
rect 14094 2479 14096 2488
rect 14148 2479 14150 2488
rect 14096 2450 14148 2456
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13176 1760 13228 1766
rect 13176 1702 13228 1708
rect 13372 814 13400 2246
rect 13556 2106 13584 2246
rect 13544 2100 13596 2106
rect 13544 2042 13596 2048
rect 13648 1902 13676 2246
rect 14292 2106 14320 2518
rect 14752 2514 14780 3538
rect 14844 3505 14872 4134
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 15108 4072 15160 4078
rect 15212 4060 15240 4626
rect 15304 4570 15332 5714
rect 15304 4542 15424 4570
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15304 4078 15332 4422
rect 15396 4146 15424 4542
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15160 4032 15240 4060
rect 15292 4072 15344 4078
rect 15108 4014 15160 4020
rect 15292 4014 15344 4020
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14830 3496 14886 3505
rect 14830 3431 14886 3440
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14280 2100 14332 2106
rect 14280 2042 14332 2048
rect 14384 1902 14412 2382
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14476 1902 14504 2246
rect 14660 1902 14688 2314
rect 13636 1896 13688 1902
rect 13636 1838 13688 1844
rect 14372 1896 14424 1902
rect 14372 1838 14424 1844
rect 14464 1896 14516 1902
rect 14464 1838 14516 1844
rect 14648 1896 14700 1902
rect 14648 1838 14700 1844
rect 14384 1766 14412 1838
rect 14372 1760 14424 1766
rect 14372 1702 14424 1708
rect 14832 1760 14884 1766
rect 14832 1702 14884 1708
rect 13830 1660 14138 1669
rect 13830 1658 13836 1660
rect 13892 1658 13916 1660
rect 13972 1658 13996 1660
rect 14052 1658 14076 1660
rect 14132 1658 14138 1660
rect 13892 1606 13894 1658
rect 14074 1606 14076 1658
rect 13830 1604 13836 1606
rect 13892 1604 13916 1606
rect 13972 1604 13996 1606
rect 14052 1604 14076 1606
rect 14132 1604 14138 1606
rect 13830 1595 14138 1604
rect 14384 1426 14412 1702
rect 14844 1562 14872 1702
rect 14832 1556 14884 1562
rect 14832 1498 14884 1504
rect 14936 1442 14964 3878
rect 15028 3602 15056 4014
rect 15396 3738 15424 4082
rect 15488 3942 15516 11494
rect 15580 10810 15608 15030
rect 15672 14958 15700 15506
rect 15948 14958 15976 15642
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15948 14278 15976 14894
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15856 13870 15884 14214
rect 16040 13938 16068 14758
rect 16132 14482 16160 16594
rect 16592 16046 16620 16594
rect 16684 16182 16712 16934
rect 16776 16726 16804 16934
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16672 16176 16724 16182
rect 16672 16118 16724 16124
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16224 15570 16252 15846
rect 16776 15570 16804 16390
rect 16960 16114 16988 16730
rect 17038 16552 17094 16561
rect 17144 16522 17172 17054
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17512 16794 17540 16934
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17328 16590 17356 16730
rect 17696 16726 17724 16934
rect 17684 16720 17736 16726
rect 17684 16662 17736 16668
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17604 16522 17816 16538
rect 17038 16487 17094 16496
rect 17132 16516 17184 16522
rect 17052 16114 17080 16487
rect 17132 16458 17184 16464
rect 17604 16516 17828 16522
rect 17604 16510 17776 16516
rect 17188 16348 17496 16357
rect 17188 16346 17194 16348
rect 17250 16346 17274 16348
rect 17330 16346 17354 16348
rect 17410 16346 17434 16348
rect 17490 16346 17496 16348
rect 17250 16294 17252 16346
rect 17432 16294 17434 16346
rect 17188 16292 17194 16294
rect 17250 16292 17274 16294
rect 17330 16292 17354 16294
rect 17410 16292 17434 16294
rect 17490 16292 17496 16294
rect 17188 16283 17496 16292
rect 17604 16232 17632 16510
rect 17776 16458 17828 16464
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17328 16204 17632 16232
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 17328 16046 17356 16204
rect 16856 16040 16908 16046
rect 16856 15982 16908 15988
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16776 15473 16804 15506
rect 16762 15464 16818 15473
rect 16762 15399 16818 15408
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16408 15201 16436 15302
rect 16394 15192 16450 15201
rect 16394 15127 16450 15136
rect 16408 15094 16436 15127
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16316 14958 16344 15030
rect 16408 14958 16436 15030
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 16120 13728 16172 13734
rect 16120 13670 16172 13676
rect 16132 13394 16160 13670
rect 16316 13462 16344 14010
rect 16408 14006 16436 14894
rect 16868 14770 16896 15982
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16960 14890 16988 15846
rect 17040 15428 17092 15434
rect 17040 15370 17092 15376
rect 17052 14958 17080 15370
rect 17188 15260 17496 15269
rect 17188 15258 17194 15260
rect 17250 15258 17274 15260
rect 17330 15258 17354 15260
rect 17410 15258 17434 15260
rect 17490 15258 17496 15260
rect 17250 15206 17252 15258
rect 17432 15206 17434 15258
rect 17188 15204 17194 15206
rect 17250 15204 17274 15206
rect 17330 15204 17354 15206
rect 17410 15204 17434 15206
rect 17490 15204 17496 15206
rect 17188 15195 17496 15204
rect 17604 15026 17632 15982
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 16948 14884 17000 14890
rect 16948 14826 17000 14832
rect 17132 14816 17184 14822
rect 16868 14742 17080 14770
rect 17132 14758 17184 14764
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16304 13456 16356 13462
rect 16304 13398 16356 13404
rect 16120 13388 16172 13394
rect 16408 13376 16436 13942
rect 16868 13870 16896 14282
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16672 13796 16724 13802
rect 16672 13738 16724 13744
rect 16684 13462 16712 13738
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 16488 13388 16540 13394
rect 16408 13348 16488 13376
rect 16120 13330 16172 13336
rect 16488 13330 16540 13336
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15948 12782 15976 13126
rect 16132 12986 16160 13330
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16316 11218 16344 12718
rect 16592 12714 16620 13194
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16856 12368 16908 12374
rect 16856 12310 16908 12316
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15672 9450 15700 10542
rect 15750 9480 15806 9489
rect 15660 9444 15712 9450
rect 15750 9415 15752 9424
rect 15660 9386 15712 9392
rect 15804 9415 15806 9424
rect 15752 9386 15804 9392
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16132 9042 16160 9318
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 15948 7546 15976 7822
rect 16132 7818 16160 8978
rect 16316 8090 16344 8978
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 16028 7336 16080 7342
rect 16132 7324 16160 7754
rect 16080 7296 16160 7324
rect 16028 7278 16080 7284
rect 16316 7274 16344 8026
rect 16408 7528 16436 12038
rect 16592 11286 16620 12106
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16500 10810 16528 11154
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16592 10742 16620 11222
rect 16684 10742 16712 11494
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 16672 10736 16724 10742
rect 16672 10678 16724 10684
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16684 10266 16712 10542
rect 16776 10266 16804 10542
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16868 10146 16896 12310
rect 16960 11558 16988 12582
rect 17052 12306 17080 14742
rect 17144 14482 17172 14758
rect 17236 14482 17264 14962
rect 17408 14884 17460 14890
rect 17460 14844 17632 14872
rect 17408 14826 17460 14832
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 17188 14172 17496 14181
rect 17188 14170 17194 14172
rect 17250 14170 17274 14172
rect 17330 14170 17354 14172
rect 17410 14170 17434 14172
rect 17490 14170 17496 14172
rect 17250 14118 17252 14170
rect 17432 14118 17434 14170
rect 17188 14116 17194 14118
rect 17250 14116 17274 14118
rect 17330 14116 17354 14118
rect 17410 14116 17434 14118
rect 17490 14116 17496 14118
rect 17188 14107 17496 14116
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17144 13802 17172 14010
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 17328 13870 17356 13942
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 17188 13084 17496 13093
rect 17188 13082 17194 13084
rect 17250 13082 17274 13084
rect 17330 13082 17354 13084
rect 17410 13082 17434 13084
rect 17490 13082 17496 13084
rect 17250 13030 17252 13082
rect 17432 13030 17434 13082
rect 17188 13028 17194 13030
rect 17250 13028 17274 13030
rect 17330 13028 17354 13030
rect 17410 13028 17434 13030
rect 17490 13028 17496 13030
rect 17188 13019 17496 13028
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 17512 12714 17540 12854
rect 17500 12708 17552 12714
rect 17500 12650 17552 12656
rect 17604 12374 17632 14844
rect 17696 14550 17724 16390
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17788 15570 17816 15982
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17880 15638 17908 15846
rect 17868 15632 17920 15638
rect 17868 15574 17920 15580
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17684 14544 17736 14550
rect 17684 14486 17736 14492
rect 17788 13802 17816 14758
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17880 13802 17908 14418
rect 17776 13796 17828 13802
rect 17776 13738 17828 13744
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17696 12306 17724 12922
rect 17788 12782 17816 13738
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17880 12374 17908 13262
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17972 12322 18000 16390
rect 18524 16250 18552 16594
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 18156 15094 18184 16050
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 18156 13433 18184 15030
rect 18248 14482 18276 15438
rect 18616 15162 18644 15506
rect 18708 15162 18736 17614
rect 18786 17600 18842 18000
rect 19430 17600 19486 18000
rect 20074 17600 20130 18000
rect 20718 17600 20774 18000
rect 21362 17762 21418 18000
rect 21362 17734 21680 17762
rect 21362 17600 21418 17734
rect 19444 17134 19472 17600
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19628 16726 19656 17206
rect 21652 17134 21680 17734
rect 22006 17600 22062 18000
rect 22650 17600 22706 18000
rect 23294 17600 23350 18000
rect 23938 17600 23994 18000
rect 24582 17600 24638 18000
rect 25226 17600 25282 18000
rect 25870 17600 25926 18000
rect 26514 17762 26570 18000
rect 26514 17734 26832 17762
rect 26514 17600 26570 17734
rect 22020 17134 22048 17600
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 22008 17128 22060 17134
rect 22008 17070 22060 17076
rect 22664 17066 22692 17600
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23112 17128 23164 17134
rect 23032 17088 23112 17116
rect 22652 17060 22704 17066
rect 22652 17002 22704 17008
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 19616 16720 19668 16726
rect 19616 16662 19668 16668
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 18880 15972 18932 15978
rect 18880 15914 18932 15920
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18340 14618 18368 14894
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18248 13870 18276 14418
rect 18340 14074 18368 14418
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18142 13424 18198 13433
rect 18142 13359 18198 13368
rect 18708 13258 18736 13806
rect 18696 13252 18748 13258
rect 18696 13194 18748 13200
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18052 12776 18104 12782
rect 18236 12776 18288 12782
rect 18052 12718 18104 12724
rect 18142 12744 18198 12753
rect 18064 12617 18092 12718
rect 18236 12718 18288 12724
rect 18142 12679 18144 12688
rect 18196 12679 18198 12688
rect 18144 12650 18196 12656
rect 18050 12608 18106 12617
rect 18050 12543 18106 12552
rect 18156 12442 18184 12650
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17592 12164 17644 12170
rect 17592 12106 17644 12112
rect 17684 12164 17736 12170
rect 17684 12106 17736 12112
rect 17188 11996 17496 12005
rect 17188 11994 17194 11996
rect 17250 11994 17274 11996
rect 17330 11994 17354 11996
rect 17410 11994 17434 11996
rect 17490 11994 17496 11996
rect 17250 11942 17252 11994
rect 17432 11942 17434 11994
rect 17188 11940 17194 11942
rect 17250 11940 17274 11942
rect 17330 11940 17354 11942
rect 17410 11940 17434 11942
rect 17490 11940 17496 11942
rect 17188 11931 17496 11940
rect 17604 11937 17632 12106
rect 17590 11928 17646 11937
rect 17590 11863 17646 11872
rect 17590 11792 17646 11801
rect 17696 11762 17724 12106
rect 17590 11727 17646 11736
rect 17684 11756 17736 11762
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 17604 11218 17632 11727
rect 17684 11698 17736 11704
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16960 10606 16988 10950
rect 17188 10908 17496 10917
rect 17188 10906 17194 10908
rect 17250 10906 17274 10908
rect 17330 10906 17354 10908
rect 17410 10906 17434 10908
rect 17490 10906 17496 10908
rect 17250 10854 17252 10906
rect 17432 10854 17434 10906
rect 17188 10852 17194 10854
rect 17250 10852 17274 10854
rect 17330 10852 17354 10854
rect 17410 10852 17434 10854
rect 17490 10852 17496 10854
rect 17188 10843 17496 10852
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16684 10118 16896 10146
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16500 8498 16528 9454
rect 16592 9353 16620 9658
rect 16578 9344 16634 9353
rect 16578 9279 16634 9288
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16684 7993 16712 10118
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16868 9602 16896 9658
rect 16776 9574 16896 9602
rect 16776 9450 16804 9574
rect 16764 9444 16816 9450
rect 16764 9386 16816 9392
rect 16856 9444 16908 9450
rect 16856 9386 16908 9392
rect 16868 9178 16896 9386
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16854 9072 16910 9081
rect 16776 8294 16804 9046
rect 16854 9007 16856 9016
rect 16908 9007 16910 9016
rect 16856 8978 16908 8984
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16670 7984 16726 7993
rect 16670 7919 16726 7928
rect 16868 7886 16896 8978
rect 16960 8838 16988 10542
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17236 10198 17264 10406
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17188 9820 17496 9829
rect 17188 9818 17194 9820
rect 17250 9818 17274 9820
rect 17330 9818 17354 9820
rect 17410 9818 17434 9820
rect 17490 9818 17496 9820
rect 17250 9766 17252 9818
rect 17432 9766 17434 9818
rect 17188 9764 17194 9766
rect 17250 9764 17274 9766
rect 17330 9764 17354 9766
rect 17410 9764 17434 9766
rect 17490 9764 17496 9766
rect 17188 9755 17496 9764
rect 17130 9344 17186 9353
rect 17130 9279 17186 9288
rect 17144 9042 17172 9279
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 17188 8732 17496 8741
rect 17188 8730 17194 8732
rect 17250 8730 17274 8732
rect 17330 8730 17354 8732
rect 17410 8730 17434 8732
rect 17490 8730 17496 8732
rect 17250 8678 17252 8730
rect 17432 8678 17434 8730
rect 17188 8676 17194 8678
rect 17250 8676 17274 8678
rect 17330 8676 17354 8678
rect 17410 8676 17434 8678
rect 17490 8676 17496 8678
rect 17188 8667 17496 8676
rect 17604 8634 17632 11154
rect 17696 10198 17724 11494
rect 17684 10192 17736 10198
rect 17684 10134 17736 10140
rect 17696 9042 17724 10134
rect 17788 9353 17816 12310
rect 17972 12294 18184 12322
rect 18156 11694 18184 12294
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 18248 11558 18276 12718
rect 18616 12628 18644 12854
rect 18708 12782 18736 13194
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18800 12628 18828 12718
rect 18616 12600 18828 12628
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17972 10674 18000 11018
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17972 10266 18000 10610
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18064 10130 18092 10406
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 17868 9376 17920 9382
rect 17774 9344 17830 9353
rect 17868 9318 17920 9324
rect 17774 9279 17830 9288
rect 17880 9042 17908 9318
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16408 7500 16528 7528
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15580 5778 15608 7142
rect 16316 6662 16344 7210
rect 16408 7002 16436 7210
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 16132 5914 16160 6122
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 15568 5772 15620 5778
rect 15620 5732 15700 5760
rect 15568 5714 15620 5720
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15580 4078 15608 4966
rect 15672 4146 15700 5732
rect 16500 4162 16528 7500
rect 16868 7410 16896 7822
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16856 7268 16908 7274
rect 16856 7210 16908 7216
rect 16868 6798 16896 7210
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16592 5234 16620 6190
rect 16960 5846 16988 8230
rect 17052 7954 17080 8366
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 17052 7342 17080 7890
rect 17188 7644 17496 7653
rect 17188 7642 17194 7644
rect 17250 7642 17274 7644
rect 17330 7642 17354 7644
rect 17410 7642 17434 7644
rect 17490 7642 17496 7644
rect 17250 7590 17252 7642
rect 17432 7590 17434 7642
rect 17188 7588 17194 7590
rect 17250 7588 17274 7590
rect 17330 7588 17354 7590
rect 17410 7588 17434 7590
rect 17490 7588 17496 7590
rect 17188 7579 17496 7588
rect 17604 7342 17632 8570
rect 17696 8537 17724 8978
rect 17682 8528 17738 8537
rect 17682 8463 17738 8472
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17788 8022 17816 8366
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 17052 6322 17080 7278
rect 17788 7206 17816 7958
rect 17880 7954 17908 8978
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17972 8430 18000 8842
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17960 7336 18012 7342
rect 18064 7324 18092 8910
rect 18156 8566 18184 10474
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18156 8090 18184 8366
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18012 7296 18184 7324
rect 17960 7278 18012 7284
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17188 6556 17496 6565
rect 17188 6554 17194 6556
rect 17250 6554 17274 6556
rect 17330 6554 17354 6556
rect 17410 6554 17434 6556
rect 17490 6554 17496 6556
rect 17250 6502 17252 6554
rect 17432 6502 17434 6554
rect 17188 6500 17194 6502
rect 17250 6500 17274 6502
rect 17330 6500 17354 6502
rect 17410 6500 17434 6502
rect 17490 6500 17496 6502
rect 17188 6491 17496 6500
rect 17604 6390 17632 7142
rect 17972 6866 18000 7142
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17696 6458 17724 6734
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17592 6384 17644 6390
rect 17512 6332 17592 6338
rect 17512 6326 17644 6332
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17512 6310 17632 6326
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16868 4622 16896 5102
rect 16948 5092 17000 5098
rect 17052 5080 17080 6258
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17236 5914 17264 6054
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17512 5778 17540 6310
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17188 5468 17496 5477
rect 17188 5466 17194 5468
rect 17250 5466 17274 5468
rect 17330 5466 17354 5468
rect 17410 5466 17434 5468
rect 17490 5466 17496 5468
rect 17250 5414 17252 5466
rect 17432 5414 17434 5466
rect 17188 5412 17194 5414
rect 17250 5412 17274 5414
rect 17330 5412 17354 5414
rect 17410 5412 17434 5414
rect 17490 5412 17496 5414
rect 17188 5403 17496 5412
rect 17604 5250 17632 5714
rect 17000 5052 17080 5080
rect 17512 5222 17632 5250
rect 16948 5034 17000 5040
rect 17512 5030 17540 5222
rect 17972 5166 18000 6802
rect 18156 5778 18184 7296
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18064 5370 18092 5714
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17222 4720 17278 4729
rect 17512 4690 17540 4966
rect 18156 4729 18184 5714
rect 18142 4720 18198 4729
rect 17222 4655 17224 4664
rect 17276 4655 17278 4664
rect 17500 4684 17552 4690
rect 17224 4626 17276 4632
rect 17500 4626 17552 4632
rect 18064 4678 18142 4706
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 17188 4380 17496 4389
rect 17188 4378 17194 4380
rect 17250 4378 17274 4380
rect 17330 4378 17354 4380
rect 17410 4378 17434 4380
rect 17490 4378 17496 4380
rect 17250 4326 17252 4378
rect 17432 4326 17434 4378
rect 17188 4324 17194 4326
rect 17250 4324 17274 4326
rect 17330 4324 17354 4326
rect 17410 4324 17434 4326
rect 17490 4324 17496 4326
rect 17188 4315 17496 4324
rect 15660 4140 15712 4146
rect 16500 4134 16620 4162
rect 15660 4082 15712 4088
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15384 3732 15436 3738
rect 15212 3692 15384 3720
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 15028 2514 15056 3538
rect 15212 2854 15240 3692
rect 15384 3674 15436 3680
rect 15292 3596 15344 3602
rect 15580 3584 15608 4014
rect 16500 3670 16528 4014
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 15344 3556 15608 3584
rect 15660 3596 15712 3602
rect 15292 3538 15344 3544
rect 15660 3538 15712 3544
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 15304 2990 15332 3538
rect 15672 3194 15700 3538
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 15028 2378 15056 2450
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 14372 1420 14424 1426
rect 14372 1362 14424 1368
rect 14844 1414 14964 1442
rect 15028 1426 15056 2314
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 15120 1902 15148 2246
rect 15212 1902 15240 2790
rect 15108 1896 15160 1902
rect 15108 1838 15160 1844
rect 15200 1896 15252 1902
rect 15200 1838 15252 1844
rect 15304 1766 15332 2926
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 15292 1760 15344 1766
rect 15292 1702 15344 1708
rect 15396 1494 15424 2450
rect 15936 2304 15988 2310
rect 15936 2246 15988 2252
rect 15660 1964 15712 1970
rect 15660 1906 15712 1912
rect 15384 1488 15436 1494
rect 15384 1430 15436 1436
rect 15672 1426 15700 1906
rect 15948 1902 15976 2246
rect 15936 1896 15988 1902
rect 15936 1838 15988 1844
rect 16040 1426 16068 3538
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 16132 2650 16160 2790
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 15016 1420 15068 1426
rect 13360 808 13412 814
rect 13360 750 13412 756
rect 13830 572 14138 581
rect 13830 570 13836 572
rect 13892 570 13916 572
rect 13972 570 13996 572
rect 14052 570 14076 572
rect 14132 570 14138 572
rect 13892 518 13894 570
rect 14074 518 14076 570
rect 13830 516 13836 518
rect 13892 516 13916 518
rect 13972 516 13996 518
rect 14052 516 14076 518
rect 14132 516 14138 518
rect 13830 507 14138 516
rect 14844 400 14872 1414
rect 15016 1362 15068 1368
rect 15660 1420 15712 1426
rect 15660 1362 15712 1368
rect 16028 1420 16080 1426
rect 16028 1362 16080 1368
rect 16592 400 16620 4134
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 17592 4004 17644 4010
rect 17592 3946 17644 3952
rect 16776 3194 16804 3946
rect 17604 3738 17632 3946
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17972 3602 18000 3878
rect 18064 3670 18092 4678
rect 18142 4655 18198 4664
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18052 3664 18104 3670
rect 18052 3606 18104 3612
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17188 3292 17496 3301
rect 17188 3290 17194 3292
rect 17250 3290 17274 3292
rect 17330 3290 17354 3292
rect 17410 3290 17434 3292
rect 17490 3290 17496 3292
rect 17250 3238 17252 3290
rect 17432 3238 17434 3290
rect 17188 3236 17194 3238
rect 17250 3236 17274 3238
rect 17330 3236 17354 3238
rect 17410 3236 17434 3238
rect 17490 3236 17496 3238
rect 17188 3227 17496 3236
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 17880 2990 17908 3470
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 3058 18092 3334
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 17236 2650 17264 2790
rect 17880 2650 17908 2926
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 17236 2514 17264 2586
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 16684 2106 16712 2382
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 16672 2100 16724 2106
rect 16672 2042 16724 2048
rect 16868 1494 16896 2246
rect 17188 2204 17496 2213
rect 17188 2202 17194 2204
rect 17250 2202 17274 2204
rect 17330 2202 17354 2204
rect 17410 2202 17434 2204
rect 17490 2202 17496 2204
rect 17250 2150 17252 2202
rect 17432 2150 17434 2202
rect 17188 2148 17194 2150
rect 17250 2148 17274 2150
rect 17330 2148 17354 2150
rect 17410 2148 17434 2150
rect 17490 2148 17496 2150
rect 17188 2139 17496 2148
rect 16856 1488 16908 1494
rect 16856 1430 16908 1436
rect 17604 1222 17632 2246
rect 17880 1902 17908 2586
rect 18064 2514 18092 2994
rect 18156 2990 18184 3878
rect 18144 2984 18196 2990
rect 18248 2961 18276 11494
rect 18340 10538 18368 12378
rect 18432 11121 18460 12378
rect 18512 12300 18564 12306
rect 18512 12242 18564 12248
rect 18524 11665 18552 12242
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18510 11656 18566 11665
rect 18800 11626 18828 11698
rect 18510 11591 18566 11600
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 18708 11529 18736 11562
rect 18694 11520 18750 11529
rect 18694 11455 18750 11464
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 18418 11112 18474 11121
rect 18418 11047 18474 11056
rect 18328 10532 18380 10538
rect 18328 10474 18380 10480
rect 18524 10266 18552 11154
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18616 10849 18644 11086
rect 18602 10840 18658 10849
rect 18602 10775 18658 10784
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18708 10062 18736 10202
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18340 9042 18368 9522
rect 18800 9518 18828 11562
rect 18892 11218 18920 15914
rect 19064 15428 19116 15434
rect 19064 15370 19116 15376
rect 19076 14822 19104 15370
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18984 12306 19012 12582
rect 19352 12434 19380 15914
rect 19536 15502 19564 16526
rect 19628 16046 19656 16662
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19536 14958 19564 15438
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19708 15088 19760 15094
rect 19628 15036 19708 15042
rect 19628 15030 19760 15036
rect 19628 15014 19748 15030
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19444 14385 19472 14486
rect 19536 14414 19564 14894
rect 19524 14408 19576 14414
rect 19430 14376 19486 14385
rect 19524 14350 19576 14356
rect 19430 14311 19486 14320
rect 19432 14272 19484 14278
rect 19628 14226 19656 15014
rect 19484 14220 19656 14226
rect 19432 14214 19656 14220
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19444 14198 19656 14214
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19444 12442 19472 12650
rect 19168 12406 19380 12434
rect 19432 12436 19484 12442
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 19168 11830 19196 12406
rect 19432 12378 19484 12384
rect 19628 12306 19656 14198
rect 19812 13870 19840 14214
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19812 12782 19840 13806
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19904 12434 19932 15302
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 19720 12406 19932 12434
rect 19616 12300 19668 12306
rect 19616 12242 19668 12248
rect 19156 11824 19208 11830
rect 19156 11766 19208 11772
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 18892 10810 18920 11154
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 18420 9104 18472 9110
rect 18420 9046 18472 9052
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18432 7818 18460 9046
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 19076 7750 19104 9114
rect 19168 9042 19196 11766
rect 19720 11370 19748 12406
rect 19996 11558 20024 12718
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 20088 11898 20116 12038
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19444 11342 19748 11370
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19260 10198 19288 11222
rect 19248 10192 19300 10198
rect 19248 10134 19300 10140
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19260 9382 19288 9590
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19260 9042 19288 9318
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19352 8634 19380 9862
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18708 6322 18736 7414
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18984 6254 19012 6598
rect 19076 6254 19104 7686
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 19352 6866 19380 7210
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 18984 5778 19012 6190
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18524 4486 18552 5102
rect 18984 5098 19012 5510
rect 19076 5370 19104 6190
rect 19168 5778 19196 6734
rect 19444 6361 19472 11342
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19536 9382 19564 11154
rect 19628 9654 19656 11154
rect 19720 10810 19748 11154
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19720 10130 19748 10202
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19720 9450 19748 10066
rect 19904 9602 19932 11154
rect 19996 10588 20024 11494
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 20088 10742 20116 11018
rect 20076 10736 20128 10742
rect 20076 10678 20128 10684
rect 20076 10600 20128 10606
rect 19996 10560 20076 10588
rect 20076 10542 20128 10548
rect 20088 9926 20116 10542
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 19904 9574 20024 9602
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19708 9444 19760 9450
rect 19708 9386 19760 9392
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19536 8906 19564 9318
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19904 8634 19932 9454
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19800 7948 19852 7954
rect 19904 7936 19932 8570
rect 19852 7908 19932 7936
rect 19800 7890 19852 7896
rect 19996 7818 20024 9574
rect 20180 9450 20208 16934
rect 20546 16892 20854 16901
rect 20546 16890 20552 16892
rect 20608 16890 20632 16892
rect 20688 16890 20712 16892
rect 20768 16890 20792 16892
rect 20848 16890 20854 16892
rect 20608 16838 20610 16890
rect 20790 16838 20792 16890
rect 20546 16836 20552 16838
rect 20608 16836 20632 16838
rect 20688 16836 20712 16838
rect 20768 16836 20792 16838
rect 20848 16836 20854 16838
rect 20546 16827 20854 16836
rect 21468 16658 21496 16934
rect 22112 16658 22140 16934
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 20824 16250 20852 16594
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20456 15366 20484 15982
rect 20546 15804 20854 15813
rect 20546 15802 20552 15804
rect 20608 15802 20632 15804
rect 20688 15802 20712 15804
rect 20768 15802 20792 15804
rect 20848 15802 20854 15804
rect 20608 15750 20610 15802
rect 20790 15750 20792 15802
rect 20546 15748 20552 15750
rect 20608 15748 20632 15750
rect 20688 15748 20712 15750
rect 20768 15748 20792 15750
rect 20848 15748 20854 15750
rect 20546 15739 20854 15748
rect 21100 15570 21128 16526
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 21100 14822 21128 15302
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 20546 14716 20854 14725
rect 20546 14714 20552 14716
rect 20608 14714 20632 14716
rect 20688 14714 20712 14716
rect 20768 14714 20792 14716
rect 20848 14714 20854 14716
rect 20608 14662 20610 14714
rect 20790 14662 20792 14714
rect 20546 14660 20552 14662
rect 20608 14660 20632 14662
rect 20688 14660 20712 14662
rect 20768 14660 20792 14662
rect 20848 14660 20854 14662
rect 20546 14651 20854 14660
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20916 14074 20944 14214
rect 21192 14074 21220 14418
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 20546 13628 20854 13637
rect 20546 13626 20552 13628
rect 20608 13626 20632 13628
rect 20688 13626 20712 13628
rect 20768 13626 20792 13628
rect 20848 13626 20854 13628
rect 20608 13574 20610 13626
rect 20790 13574 20792 13626
rect 20546 13572 20552 13574
rect 20608 13572 20632 13574
rect 20688 13572 20712 13574
rect 20768 13572 20792 13574
rect 20848 13572 20854 13574
rect 20546 13563 20854 13572
rect 20916 13394 20944 14010
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20364 12306 20392 12378
rect 20456 12306 20484 12922
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 20546 12540 20854 12549
rect 20546 12538 20552 12540
rect 20608 12538 20632 12540
rect 20688 12538 20712 12540
rect 20768 12538 20792 12540
rect 20848 12538 20854 12540
rect 20608 12486 20610 12538
rect 20790 12486 20792 12538
rect 20546 12484 20552 12486
rect 20608 12484 20632 12486
rect 20688 12484 20712 12486
rect 20768 12484 20792 12486
rect 20848 12484 20854 12486
rect 20546 12475 20854 12484
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20168 9444 20220 9450
rect 20168 9386 20220 9392
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19904 6866 19932 7142
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19430 6352 19486 6361
rect 19430 6287 19486 6296
rect 19248 6180 19300 6186
rect 19248 6122 19300 6128
rect 19260 5778 19288 6122
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 19352 5098 19380 6054
rect 19708 5908 19760 5914
rect 19708 5850 19760 5856
rect 19720 5710 19748 5850
rect 20272 5760 20300 12038
rect 20364 11830 20392 12242
rect 21008 12238 21036 12786
rect 21100 12345 21128 13194
rect 21192 12782 21220 14010
rect 21284 13870 21312 15846
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21284 13326 21312 13806
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21284 12850 21312 13262
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 21086 12336 21142 12345
rect 21086 12271 21142 12280
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 20352 11824 20404 11830
rect 20352 11766 20404 11772
rect 20546 11452 20854 11461
rect 20546 11450 20552 11452
rect 20608 11450 20632 11452
rect 20688 11450 20712 11452
rect 20768 11450 20792 11452
rect 20848 11450 20854 11452
rect 20608 11398 20610 11450
rect 20790 11398 20792 11450
rect 20546 11396 20552 11398
rect 20608 11396 20632 11398
rect 20688 11396 20712 11398
rect 20768 11396 20792 11398
rect 20848 11396 20854 11398
rect 20546 11387 20854 11396
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20548 10713 20576 11086
rect 21284 10810 21312 11834
rect 21376 11257 21404 13874
rect 21468 13870 21496 14758
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 21548 13864 21600 13870
rect 21548 13806 21600 13812
rect 21560 13462 21588 13806
rect 21548 13456 21600 13462
rect 21548 13398 21600 13404
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21468 11354 21496 12786
rect 21560 12782 21588 13398
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 21560 12374 21588 12718
rect 21548 12368 21600 12374
rect 21548 12310 21600 12316
rect 21652 12238 21680 16594
rect 21928 13938 21956 16594
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22112 14618 22140 15506
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 22192 14476 22244 14482
rect 22192 14418 22244 14424
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 22204 12434 22232 14418
rect 22296 13326 22324 16662
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 22388 14074 22416 14418
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22388 13841 22416 13874
rect 22374 13832 22430 13841
rect 22374 13767 22430 13776
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 22480 12850 22508 16594
rect 22756 15994 22784 16934
rect 22940 16658 22968 16934
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 23032 16590 23060 17088
rect 23112 17070 23164 17076
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 23032 16046 23060 16526
rect 22664 15966 22784 15994
rect 23020 16040 23072 16046
rect 23020 15982 23072 15988
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22572 12434 22600 13262
rect 22112 12406 22232 12434
rect 22296 12406 22600 12434
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21652 11830 21680 12174
rect 21640 11824 21692 11830
rect 21640 11766 21692 11772
rect 21546 11656 21602 11665
rect 21546 11591 21602 11600
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21560 11286 21588 11591
rect 21548 11280 21600 11286
rect 21362 11248 21418 11257
rect 21548 11222 21600 11228
rect 21362 11183 21418 11192
rect 22112 10810 22140 12406
rect 22192 11620 22244 11626
rect 22192 11562 22244 11568
rect 22204 10810 22232 11562
rect 21272 10804 21324 10810
rect 22100 10804 22152 10810
rect 21324 10764 21496 10792
rect 21272 10746 21324 10752
rect 20534 10704 20590 10713
rect 21468 10674 21496 10764
rect 22100 10746 22152 10752
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 20534 10639 20590 10648
rect 21456 10668 21508 10674
rect 20548 10606 20576 10639
rect 21456 10610 21508 10616
rect 20352 10600 20404 10606
rect 20536 10600 20588 10606
rect 20352 10542 20404 10548
rect 20456 10560 20536 10588
rect 20364 9994 20392 10542
rect 20352 9988 20404 9994
rect 20352 9930 20404 9936
rect 20456 8090 20484 10560
rect 20536 10542 20588 10548
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20546 10364 20854 10373
rect 20546 10362 20552 10364
rect 20608 10362 20632 10364
rect 20688 10362 20712 10364
rect 20768 10362 20792 10364
rect 20848 10362 20854 10364
rect 20608 10310 20610 10362
rect 20790 10310 20792 10362
rect 20546 10308 20552 10310
rect 20608 10308 20632 10310
rect 20688 10308 20712 10310
rect 20768 10308 20792 10310
rect 20848 10308 20854 10310
rect 20546 10299 20854 10308
rect 20916 10198 20944 10406
rect 20904 10192 20956 10198
rect 20956 10152 21036 10180
rect 20904 10134 20956 10140
rect 20902 9616 20958 9625
rect 20902 9551 20958 9560
rect 20916 9518 20944 9551
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20546 9276 20854 9285
rect 20546 9274 20552 9276
rect 20608 9274 20632 9276
rect 20688 9274 20712 9276
rect 20768 9274 20792 9276
rect 20848 9274 20854 9276
rect 20608 9222 20610 9274
rect 20790 9222 20792 9274
rect 20546 9220 20552 9222
rect 20608 9220 20632 9222
rect 20688 9220 20712 9222
rect 20768 9220 20792 9222
rect 20848 9220 20854 9222
rect 20546 9211 20854 9220
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20640 8362 20668 8774
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 20546 8188 20854 8197
rect 20546 8186 20552 8188
rect 20608 8186 20632 8188
rect 20688 8186 20712 8188
rect 20768 8186 20792 8188
rect 20848 8186 20854 8188
rect 20608 8134 20610 8186
rect 20790 8134 20792 8186
rect 20546 8132 20552 8134
rect 20608 8132 20632 8134
rect 20688 8132 20712 8134
rect 20768 8132 20792 8134
rect 20848 8132 20854 8134
rect 20546 8123 20854 8132
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 20364 7954 20392 8026
rect 20916 7954 20944 8298
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 20640 7546 20668 7890
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 21008 7478 21036 10152
rect 21100 9926 21128 10542
rect 21456 10532 21508 10538
rect 21456 10474 21508 10480
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21088 9920 21140 9926
rect 21088 9862 21140 9868
rect 21100 9382 21128 9862
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 21192 8945 21220 9454
rect 21178 8936 21234 8945
rect 21178 8871 21234 8880
rect 21192 8634 21220 8871
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21284 8294 21312 10406
rect 21468 9518 21496 10474
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21560 9722 21588 10066
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21456 9512 21508 9518
rect 21456 9454 21508 9460
rect 21836 9110 21864 10406
rect 22192 9716 22244 9722
rect 22192 9658 22244 9664
rect 22204 9518 22232 9658
rect 22192 9512 22244 9518
rect 22192 9454 22244 9460
rect 21548 9104 21600 9110
rect 21548 9046 21600 9052
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 21284 7818 21312 8230
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 21100 7546 21128 7754
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20996 7472 21048 7478
rect 20996 7414 21048 7420
rect 20546 7100 20854 7109
rect 20546 7098 20552 7100
rect 20608 7098 20632 7100
rect 20688 7098 20712 7100
rect 20768 7098 20792 7100
rect 20848 7098 20854 7100
rect 20608 7046 20610 7098
rect 20790 7046 20792 7098
rect 20546 7044 20552 7046
rect 20608 7044 20632 7046
rect 20688 7044 20712 7046
rect 20768 7044 20792 7046
rect 20848 7044 20854 7046
rect 20546 7035 20854 7044
rect 21008 6866 21036 7414
rect 21560 7342 21588 9046
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 21456 6860 21508 6866
rect 21456 6802 21508 6808
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20364 5778 20392 6054
rect 20456 5914 20484 6054
rect 20546 6012 20854 6021
rect 20546 6010 20552 6012
rect 20608 6010 20632 6012
rect 20688 6010 20712 6012
rect 20768 6010 20792 6012
rect 20848 6010 20854 6012
rect 20608 5958 20610 6010
rect 20790 5958 20792 6010
rect 20546 5956 20552 5958
rect 20608 5956 20632 5958
rect 20688 5956 20712 5958
rect 20768 5956 20792 5958
rect 20848 5956 20854 5958
rect 20546 5947 20854 5956
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20180 5732 20300 5760
rect 20352 5772 20404 5778
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19430 5264 19486 5273
rect 19430 5199 19486 5208
rect 18972 5092 19024 5098
rect 18972 5034 19024 5040
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18524 4078 18552 4422
rect 18512 4072 18564 4078
rect 18326 4040 18382 4049
rect 18512 4014 18564 4020
rect 18326 3975 18382 3984
rect 18144 2926 18196 2932
rect 18234 2952 18290 2961
rect 18234 2887 18290 2896
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 18064 1902 18092 2314
rect 18144 2032 18196 2038
rect 18144 1974 18196 1980
rect 18156 1902 18184 1974
rect 17868 1896 17920 1902
rect 17682 1864 17738 1873
rect 17868 1838 17920 1844
rect 18052 1896 18104 1902
rect 18052 1838 18104 1844
rect 18144 1896 18196 1902
rect 18144 1838 18196 1844
rect 17682 1799 17738 1808
rect 17960 1828 18012 1834
rect 17696 1222 17724 1799
rect 17960 1770 18012 1776
rect 17972 1290 18000 1770
rect 17960 1284 18012 1290
rect 17960 1226 18012 1232
rect 17592 1216 17644 1222
rect 17592 1158 17644 1164
rect 17684 1216 17736 1222
rect 17684 1158 17736 1164
rect 17188 1116 17496 1125
rect 17188 1114 17194 1116
rect 17250 1114 17274 1116
rect 17330 1114 17354 1116
rect 17410 1114 17434 1116
rect 17490 1114 17496 1116
rect 17250 1062 17252 1114
rect 17432 1062 17434 1114
rect 17188 1060 17194 1062
rect 17250 1060 17274 1062
rect 17330 1060 17354 1062
rect 17410 1060 17434 1062
rect 17490 1060 17496 1062
rect 17188 1051 17496 1060
rect 17696 882 17724 1158
rect 17684 876 17736 882
rect 17684 818 17736 824
rect 18340 400 18368 3975
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 18432 2990 18460 3674
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 18432 2038 18460 2926
rect 18524 2446 18552 4014
rect 18616 3602 18644 4762
rect 19444 4758 19472 5199
rect 19892 5160 19944 5166
rect 19892 5102 19944 5108
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19904 4570 19932 5102
rect 19996 5030 20024 5510
rect 20088 5370 20116 5646
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19996 4690 20024 4966
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19904 4542 20024 4570
rect 19996 4146 20024 4542
rect 20074 4176 20130 4185
rect 19984 4140 20036 4146
rect 20074 4111 20130 4120
rect 19984 4082 20036 4088
rect 19064 4004 19116 4010
rect 19064 3946 19116 3952
rect 19076 3738 19104 3946
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 19996 2990 20024 4082
rect 20088 3942 20116 4111
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18420 2032 18472 2038
rect 18418 2000 18420 2009
rect 18472 2000 18474 2009
rect 18418 1935 18474 1944
rect 18524 1494 18552 2382
rect 18708 2106 18736 2926
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19352 2582 19380 2790
rect 19996 2774 20024 2926
rect 20180 2774 20208 5732
rect 20352 5714 20404 5720
rect 20260 5636 20312 5642
rect 20260 5578 20312 5584
rect 20272 5166 20300 5578
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20272 4690 20300 4966
rect 20364 4690 20392 5714
rect 20456 5386 20484 5850
rect 20904 5840 20956 5846
rect 20904 5782 20956 5788
rect 20456 5358 20576 5386
rect 20548 5030 20576 5358
rect 20916 5030 20944 5782
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 21008 5166 21036 5510
rect 21086 5264 21142 5273
rect 21086 5199 21142 5208
rect 21100 5166 21128 5199
rect 21284 5166 21312 6394
rect 21468 5760 21496 6802
rect 21560 5953 21588 7278
rect 21652 7002 21680 7278
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21744 6322 21772 6598
rect 22112 6390 22140 7958
rect 21916 6384 21968 6390
rect 21916 6326 21968 6332
rect 22100 6384 22152 6390
rect 22100 6326 22152 6332
rect 21732 6316 21784 6322
rect 21732 6258 21784 6264
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 21546 5944 21602 5953
rect 21546 5879 21548 5888
rect 21600 5879 21602 5888
rect 21548 5850 21600 5856
rect 21548 5772 21600 5778
rect 21468 5732 21548 5760
rect 21548 5714 21600 5720
rect 21560 5642 21588 5714
rect 21548 5636 21600 5642
rect 21548 5578 21600 5584
rect 21652 5370 21680 6190
rect 21640 5364 21692 5370
rect 21640 5306 21692 5312
rect 21744 5302 21772 6258
rect 21928 5914 21956 6326
rect 22112 6254 22140 6326
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 21916 5908 21968 5914
rect 21916 5850 21968 5856
rect 21836 5778 22140 5794
rect 21824 5772 22140 5778
rect 21876 5766 22140 5772
rect 21824 5714 21876 5720
rect 22112 5710 22140 5766
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 21732 5296 21784 5302
rect 21732 5238 21784 5244
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 21364 5092 21416 5098
rect 21364 5034 21416 5040
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20546 4924 20854 4933
rect 20546 4922 20552 4924
rect 20608 4922 20632 4924
rect 20688 4922 20712 4924
rect 20768 4922 20792 4924
rect 20848 4922 20854 4924
rect 20608 4870 20610 4922
rect 20790 4870 20792 4922
rect 20546 4868 20552 4870
rect 20608 4868 20632 4870
rect 20688 4868 20712 4870
rect 20768 4868 20792 4870
rect 20848 4868 20854 4870
rect 20546 4859 20854 4868
rect 20916 4690 20944 4966
rect 20260 4684 20312 4690
rect 20260 4626 20312 4632
rect 20352 4684 20404 4690
rect 20352 4626 20404 4632
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 21376 4486 21404 5034
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21100 4078 21128 4422
rect 21744 4282 21772 5238
rect 21916 4480 21968 4486
rect 21916 4422 21968 4428
rect 21732 4276 21784 4282
rect 21732 4218 21784 4224
rect 21088 4072 21140 4078
rect 21088 4014 21140 4020
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20272 3602 20300 3878
rect 20546 3836 20854 3845
rect 20546 3834 20552 3836
rect 20608 3834 20632 3836
rect 20688 3834 20712 3836
rect 20768 3834 20792 3836
rect 20848 3834 20854 3836
rect 20608 3782 20610 3834
rect 20790 3782 20792 3834
rect 20546 3780 20552 3782
rect 20608 3780 20632 3782
rect 20688 3780 20712 3782
rect 20768 3780 20792 3782
rect 20848 3780 20854 3782
rect 20546 3771 20854 3780
rect 21928 3602 21956 4422
rect 22204 4078 22232 6054
rect 22192 4072 22244 4078
rect 22112 4020 22192 4026
rect 22112 4014 22244 4020
rect 22112 3998 22232 4014
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 21548 3596 21600 3602
rect 21548 3538 21600 3544
rect 21732 3596 21784 3602
rect 21732 3538 21784 3544
rect 21916 3596 21968 3602
rect 21968 3556 22048 3584
rect 21916 3538 21968 3544
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 20364 2922 20392 3334
rect 21560 3194 21588 3538
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 20352 2916 20404 2922
rect 20352 2858 20404 2864
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 19904 2746 20024 2774
rect 20088 2746 20208 2774
rect 20546 2748 20854 2757
rect 20546 2746 20552 2748
rect 20608 2746 20632 2748
rect 20688 2746 20712 2748
rect 20768 2746 20792 2748
rect 20848 2746 20854 2748
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19340 2576 19392 2582
rect 19340 2518 19392 2524
rect 18696 2100 18748 2106
rect 18696 2042 18748 2048
rect 19062 2000 19118 2009
rect 19062 1935 19118 1944
rect 19076 1902 19104 1935
rect 19444 1902 19472 2586
rect 19904 1970 19932 2746
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19996 2038 20024 2246
rect 19984 2032 20036 2038
rect 19984 1974 20036 1980
rect 19892 1964 19944 1970
rect 19892 1906 19944 1912
rect 18972 1896 19024 1902
rect 18972 1838 19024 1844
rect 19064 1896 19116 1902
rect 19064 1838 19116 1844
rect 19432 1896 19484 1902
rect 19432 1838 19484 1844
rect 18696 1760 18748 1766
rect 18696 1702 18748 1708
rect 18512 1488 18564 1494
rect 18512 1430 18564 1436
rect 18708 882 18736 1702
rect 18984 1018 19012 1838
rect 18972 1012 19024 1018
rect 18972 954 19024 960
rect 19076 882 19104 1838
rect 19340 1216 19392 1222
rect 19340 1158 19392 1164
rect 19352 1018 19380 1158
rect 19340 1012 19392 1018
rect 19340 954 19392 960
rect 18696 876 18748 882
rect 18696 818 18748 824
rect 19064 876 19116 882
rect 19064 818 19116 824
rect 19444 814 19472 1838
rect 19616 1556 19668 1562
rect 19616 1498 19668 1504
rect 19628 814 19656 1498
rect 19904 1426 19932 1906
rect 19800 1420 19852 1426
rect 19800 1362 19852 1368
rect 19892 1420 19944 1426
rect 19892 1362 19944 1368
rect 19812 1018 19840 1362
rect 19800 1012 19852 1018
rect 19800 954 19852 960
rect 19432 808 19484 814
rect 19432 750 19484 756
rect 19616 808 19668 814
rect 19616 750 19668 756
rect 20088 400 20116 2746
rect 20608 2694 20610 2746
rect 20790 2694 20792 2746
rect 20546 2692 20552 2694
rect 20608 2692 20632 2694
rect 20688 2692 20712 2694
rect 20768 2692 20792 2694
rect 20848 2692 20854 2694
rect 20546 2683 20854 2692
rect 21468 2514 21496 2790
rect 21456 2508 21508 2514
rect 21456 2450 21508 2456
rect 20904 1896 20956 1902
rect 20904 1838 20956 1844
rect 20546 1660 20854 1669
rect 20546 1658 20552 1660
rect 20608 1658 20632 1660
rect 20688 1658 20712 1660
rect 20768 1658 20792 1660
rect 20848 1658 20854 1660
rect 20608 1606 20610 1658
rect 20790 1606 20792 1658
rect 20546 1604 20552 1606
rect 20608 1604 20632 1606
rect 20688 1604 20712 1606
rect 20768 1604 20792 1606
rect 20848 1604 20854 1606
rect 20546 1595 20854 1604
rect 20916 814 20944 1838
rect 21652 814 21680 3130
rect 21744 2650 21772 3538
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 21836 2990 21864 3402
rect 21916 3392 21968 3398
rect 21916 3334 21968 3340
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 21732 2644 21784 2650
rect 21732 2586 21784 2592
rect 21836 2514 21864 2926
rect 21824 2508 21876 2514
rect 21824 2450 21876 2456
rect 21928 2394 21956 3334
rect 22020 3126 22048 3556
rect 22008 3120 22060 3126
rect 22008 3062 22060 3068
rect 22112 2530 22140 3998
rect 22296 3398 22324 12406
rect 22664 12050 22692 15966
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 22756 12442 22784 15846
rect 23124 15706 23152 15982
rect 23216 15706 23244 17478
rect 23308 17202 23336 17600
rect 23952 17542 23980 17600
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 24308 17536 24360 17542
rect 24308 17478 24360 17484
rect 23904 17436 24212 17445
rect 23904 17434 23910 17436
rect 23966 17434 23990 17436
rect 24046 17434 24070 17436
rect 24126 17434 24150 17436
rect 24206 17434 24212 17436
rect 23966 17382 23968 17434
rect 24148 17382 24150 17434
rect 23904 17380 23910 17382
rect 23966 17380 23990 17382
rect 24046 17380 24070 17382
rect 24126 17380 24150 17382
rect 24206 17380 24212 17382
rect 23904 17371 24212 17380
rect 23296 17196 23348 17202
rect 23296 17138 23348 17144
rect 24320 17134 24348 17478
rect 24596 17134 24624 17600
rect 25240 17134 25268 17600
rect 25884 17134 25912 17600
rect 26804 17134 26832 17734
rect 27158 17600 27214 18000
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 25228 17128 25280 17134
rect 25228 17070 25280 17076
rect 25872 17128 25924 17134
rect 25872 17070 25924 17076
rect 26792 17128 26844 17134
rect 26792 17070 26844 17076
rect 23664 17060 23716 17066
rect 23664 17002 23716 17008
rect 26608 17060 26660 17066
rect 26608 17002 26660 17008
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23480 16788 23532 16794
rect 23480 16730 23532 16736
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 22836 15428 22888 15434
rect 22836 15370 22888 15376
rect 22848 14482 22876 15370
rect 22836 14476 22888 14482
rect 22836 14418 22888 14424
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 23020 12436 23072 12442
rect 23020 12378 23072 12384
rect 22572 12022 22692 12050
rect 22572 11665 22600 12022
rect 23032 11762 23060 12378
rect 23124 12102 23152 15642
rect 23216 15570 23244 15642
rect 23204 15564 23256 15570
rect 23204 15506 23256 15512
rect 23492 15065 23520 16730
rect 23584 16658 23612 16934
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23584 15994 23612 16186
rect 23676 16114 23704 17002
rect 25320 16992 25372 16998
rect 25320 16934 25372 16940
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 25332 16726 25360 16934
rect 25320 16720 25372 16726
rect 25320 16662 25372 16668
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23584 15966 23704 15994
rect 23676 15910 23704 15966
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23478 15056 23534 15065
rect 23478 14991 23534 15000
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23308 14346 23336 14418
rect 23478 14376 23534 14385
rect 23296 14340 23348 14346
rect 23478 14311 23534 14320
rect 23296 14282 23348 14288
rect 23308 13870 23336 14282
rect 23492 14074 23520 14311
rect 23676 14278 23704 15846
rect 23768 15162 23796 16594
rect 24584 16448 24636 16454
rect 24584 16390 24636 16396
rect 23904 16348 24212 16357
rect 23904 16346 23910 16348
rect 23966 16346 23990 16348
rect 24046 16346 24070 16348
rect 24126 16346 24150 16348
rect 24206 16346 24212 16348
rect 23966 16294 23968 16346
rect 24148 16294 24150 16346
rect 23904 16292 23910 16294
rect 23966 16292 23990 16294
rect 24046 16292 24070 16294
rect 24126 16292 24150 16294
rect 24206 16292 24212 16294
rect 23904 16283 24212 16292
rect 23904 15260 24212 15269
rect 23904 15258 23910 15260
rect 23966 15258 23990 15260
rect 24046 15258 24070 15260
rect 24126 15258 24150 15260
rect 24206 15258 24212 15260
rect 23966 15206 23968 15258
rect 24148 15206 24150 15258
rect 23904 15204 23910 15206
rect 23966 15204 23990 15206
rect 24046 15204 24070 15206
rect 24126 15204 24150 15206
rect 24206 15204 24212 15206
rect 23904 15195 24212 15204
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 24492 15020 24544 15026
rect 24492 14962 24544 14968
rect 24032 14952 24084 14958
rect 24032 14894 24084 14900
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23952 14550 23980 14758
rect 23940 14544 23992 14550
rect 23940 14486 23992 14492
rect 24044 14414 24072 14894
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24032 14408 24084 14414
rect 24032 14350 24084 14356
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23904 14172 24212 14181
rect 23904 14170 23910 14172
rect 23966 14170 23990 14172
rect 24046 14170 24070 14172
rect 24126 14170 24150 14172
rect 24206 14170 24212 14172
rect 23966 14118 23968 14170
rect 24148 14118 24150 14170
rect 23904 14116 23910 14118
rect 23966 14116 23990 14118
rect 24046 14116 24070 14118
rect 24126 14116 24150 14118
rect 24206 14116 24212 14118
rect 23904 14107 24212 14116
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 24044 13394 24072 14010
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 24308 13320 24360 13326
rect 24308 13262 24360 13268
rect 23768 12986 23796 13262
rect 23904 13084 24212 13093
rect 23904 13082 23910 13084
rect 23966 13082 23990 13084
rect 24046 13082 24070 13084
rect 24126 13082 24150 13084
rect 24206 13082 24212 13084
rect 23966 13030 23968 13082
rect 24148 13030 24150 13082
rect 23904 13028 23910 13030
rect 23966 13028 23990 13030
rect 24046 13028 24070 13030
rect 24126 13028 24150 13030
rect 24206 13028 24212 13030
rect 23904 13019 24212 13028
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23296 12708 23348 12714
rect 23296 12650 23348 12656
rect 23308 12434 23336 12650
rect 23308 12406 23428 12434
rect 23296 12232 23348 12238
rect 23296 12174 23348 12180
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 22652 11688 22704 11694
rect 22558 11656 22614 11665
rect 22652 11630 22704 11636
rect 22558 11591 22614 11600
rect 22664 11218 22692 11630
rect 23124 11626 23152 12038
rect 23308 11694 23336 12174
rect 23296 11688 23348 11694
rect 23296 11630 23348 11636
rect 23112 11620 23164 11626
rect 23112 11562 23164 11568
rect 22744 11552 22796 11558
rect 22744 11494 22796 11500
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22558 11112 22614 11121
rect 22558 11047 22614 11056
rect 22572 11014 22600 11047
rect 22560 11008 22612 11014
rect 22560 10950 22612 10956
rect 22572 10674 22600 10950
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22388 8378 22416 10542
rect 22664 10198 22692 11154
rect 22756 10606 22784 11494
rect 23308 11354 23336 11630
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 22928 10736 22980 10742
rect 22928 10678 22980 10684
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 22652 10192 22704 10198
rect 22652 10134 22704 10140
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22572 9926 22600 9998
rect 22560 9920 22612 9926
rect 22560 9862 22612 9868
rect 22572 9722 22600 9862
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22468 9512 22520 9518
rect 22468 9454 22520 9460
rect 22480 9042 22508 9454
rect 22468 9036 22520 9042
rect 22468 8978 22520 8984
rect 22480 8634 22508 8978
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22664 8498 22692 10134
rect 22756 9926 22784 10202
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22848 9654 22876 10406
rect 22940 10062 22968 10678
rect 23308 10266 23336 11290
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 22928 10056 22980 10062
rect 22928 9998 22980 10004
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22836 9648 22888 9654
rect 22836 9590 22888 9596
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22388 8350 22508 8378
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22388 7954 22416 8230
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22480 7750 22508 8350
rect 22664 7954 22692 8434
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22480 7478 22508 7686
rect 22468 7472 22520 7478
rect 22468 7414 22520 7420
rect 22940 7426 22968 9862
rect 23032 9722 23060 10066
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 23020 8424 23072 8430
rect 23020 8366 23072 8372
rect 23032 8090 23060 8366
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 23032 7546 23060 7890
rect 23216 7546 23244 7890
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 22940 7398 23060 7426
rect 22376 7268 22428 7274
rect 22376 7210 22428 7216
rect 22388 6322 22416 7210
rect 23032 7206 23060 7398
rect 23020 7200 23072 7206
rect 23020 7142 23072 7148
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 22376 6180 22428 6186
rect 22376 6122 22428 6128
rect 22388 5953 22416 6122
rect 22374 5944 22430 5953
rect 22374 5879 22430 5888
rect 22388 5778 22416 5879
rect 23032 5778 23060 7142
rect 23296 6792 23348 6798
rect 23296 6734 23348 6740
rect 23308 6458 23336 6734
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23204 6112 23256 6118
rect 23204 6054 23256 6060
rect 22376 5772 22428 5778
rect 22376 5714 22428 5720
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 23020 5772 23072 5778
rect 23020 5714 23072 5720
rect 22664 5574 22692 5714
rect 22756 5642 22784 5714
rect 22744 5636 22796 5642
rect 22744 5578 22796 5584
rect 22652 5568 22704 5574
rect 22652 5510 22704 5516
rect 22376 5092 22428 5098
rect 22376 5034 22428 5040
rect 22388 4690 22416 5034
rect 22664 4826 22692 5510
rect 22928 5160 22980 5166
rect 22928 5102 22980 5108
rect 22836 5024 22888 5030
rect 22836 4966 22888 4972
rect 22652 4820 22704 4826
rect 22652 4762 22704 4768
rect 22376 4684 22428 4690
rect 22376 4626 22428 4632
rect 22388 4026 22416 4626
rect 22664 4214 22692 4762
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22756 4282 22784 4558
rect 22848 4282 22876 4966
rect 22940 4826 22968 5102
rect 22928 4820 22980 4826
rect 22928 4762 22980 4768
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 22652 4208 22704 4214
rect 22652 4150 22704 4156
rect 22560 4072 22612 4078
rect 22388 3998 22508 4026
rect 22560 4014 22612 4020
rect 22376 3596 22428 3602
rect 22376 3538 22428 3544
rect 22284 3392 22336 3398
rect 22284 3334 22336 3340
rect 22388 3194 22416 3538
rect 22480 3534 22508 3998
rect 22572 3777 22600 4014
rect 22664 4010 22692 4150
rect 22848 4078 22876 4218
rect 23032 4078 23060 5714
rect 23112 5568 23164 5574
rect 23112 5510 23164 5516
rect 23124 5166 23152 5510
rect 23216 5166 23244 6054
rect 23112 5160 23164 5166
rect 23112 5102 23164 5108
rect 23204 5160 23256 5166
rect 23204 5102 23256 5108
rect 23296 4276 23348 4282
rect 23296 4218 23348 4224
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 22652 4004 22704 4010
rect 22652 3946 22704 3952
rect 22558 3768 22614 3777
rect 22558 3703 22614 3712
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22376 3188 22428 3194
rect 22376 3130 22428 3136
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 22192 2848 22244 2854
rect 22192 2790 22244 2796
rect 22020 2514 22140 2530
rect 22204 2514 22232 2790
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 22388 2514 22416 2586
rect 22480 2514 22508 2994
rect 22664 2650 22692 3946
rect 22848 2854 22876 4014
rect 23216 3942 23244 4082
rect 23308 4078 23336 4218
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 23400 4026 23428 12406
rect 23492 12238 23520 12854
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23664 12640 23716 12646
rect 23584 12588 23664 12594
rect 23584 12582 23716 12588
rect 23584 12566 23704 12582
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23584 12102 23612 12566
rect 23768 12434 23796 12718
rect 23676 12406 23796 12434
rect 23676 12374 23704 12406
rect 23664 12368 23716 12374
rect 23664 12310 23716 12316
rect 23676 12102 23704 12310
rect 23756 12300 23808 12306
rect 23756 12242 23808 12248
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23664 12096 23716 12102
rect 23664 12038 23716 12044
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23492 11286 23520 11834
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23492 10198 23520 11222
rect 23584 11150 23612 12038
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23572 11008 23624 11014
rect 23572 10950 23624 10956
rect 23584 10538 23612 10950
rect 23572 10532 23624 10538
rect 23572 10474 23624 10480
rect 23480 10192 23532 10198
rect 23480 10134 23532 10140
rect 23676 9994 23704 12038
rect 23768 11898 23796 12242
rect 23904 11996 24212 12005
rect 23904 11994 23910 11996
rect 23966 11994 23990 11996
rect 24046 11994 24070 11996
rect 24126 11994 24150 11996
rect 24206 11994 24212 11996
rect 23966 11942 23968 11994
rect 24148 11942 24150 11994
rect 23904 11940 23910 11942
rect 23966 11940 23990 11942
rect 24046 11940 24070 11942
rect 24126 11940 24150 11942
rect 24206 11940 24212 11942
rect 23904 11931 24212 11940
rect 23756 11892 23808 11898
rect 24320 11880 24348 13262
rect 24412 12714 24440 14758
rect 24504 14482 24532 14962
rect 24492 14476 24544 14482
rect 24492 14418 24544 14424
rect 24400 12708 24452 12714
rect 24400 12650 24452 12656
rect 23756 11834 23808 11840
rect 24136 11852 24348 11880
rect 24136 11150 24164 11852
rect 24412 11762 24440 12650
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24228 11286 24256 11698
rect 24308 11552 24360 11558
rect 24308 11494 24360 11500
rect 24216 11280 24268 11286
rect 24216 11222 24268 11228
rect 24228 11150 24256 11222
rect 24320 11150 24348 11494
rect 24504 11354 24532 12242
rect 24596 12209 24624 16390
rect 24688 14890 24716 16594
rect 24768 15564 24820 15570
rect 24768 15506 24820 15512
rect 24780 15162 24808 15506
rect 25056 15366 25084 16594
rect 25976 16182 26004 16934
rect 25964 16176 26016 16182
rect 25964 16118 26016 16124
rect 26620 16046 26648 17002
rect 26608 16040 26660 16046
rect 26608 15982 26660 15988
rect 25228 15632 25280 15638
rect 25228 15574 25280 15580
rect 25044 15360 25096 15366
rect 25044 15302 25096 15308
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24860 14952 24912 14958
rect 24860 14894 24912 14900
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 24688 14346 24716 14826
rect 24676 14340 24728 14346
rect 24676 14282 24728 14288
rect 24872 13920 24900 14894
rect 24964 14618 24992 14894
rect 25056 14822 25084 15302
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 24872 13892 24992 13920
rect 24860 13796 24912 13802
rect 24860 13738 24912 13744
rect 24872 13530 24900 13738
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 24964 13326 24992 13892
rect 25056 13394 25084 14758
rect 25240 14550 25268 15574
rect 25412 15088 25464 15094
rect 25412 15030 25464 15036
rect 25228 14544 25280 14550
rect 25228 14486 25280 14492
rect 25240 13938 25268 14486
rect 25424 14074 25452 15030
rect 25504 14476 25556 14482
rect 25504 14418 25556 14424
rect 25516 14074 25544 14418
rect 25596 14272 25648 14278
rect 25596 14214 25648 14220
rect 25608 14074 25636 14214
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 24768 13184 24820 13190
rect 24768 13126 24820 13132
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 24582 12200 24638 12209
rect 24582 12135 24638 12144
rect 24492 11348 24544 11354
rect 24492 11290 24544 11296
rect 24780 11268 24808 13126
rect 24964 12986 24992 13126
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 25044 12912 25096 12918
rect 24964 12860 25044 12866
rect 24964 12854 25096 12860
rect 24964 12838 25084 12854
rect 25148 12850 25176 13806
rect 25240 12850 25268 13874
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 25424 13394 25452 13806
rect 25596 13796 25648 13802
rect 25596 13738 25648 13744
rect 25412 13388 25464 13394
rect 25412 13330 25464 13336
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25136 12844 25188 12850
rect 24964 12442 24992 12838
rect 25136 12786 25188 12792
rect 25228 12844 25280 12850
rect 25228 12786 25280 12792
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 24952 12436 25004 12442
rect 24952 12378 25004 12384
rect 25056 12374 25084 12582
rect 25240 12434 25268 12786
rect 25332 12753 25360 13262
rect 25424 12918 25452 13330
rect 25412 12912 25464 12918
rect 25412 12854 25464 12860
rect 25424 12782 25452 12854
rect 25412 12776 25464 12782
rect 25318 12744 25374 12753
rect 25412 12718 25464 12724
rect 25608 12714 25636 13738
rect 25792 13394 25820 13874
rect 25872 13864 25924 13870
rect 27172 13841 27200 17600
rect 27262 16892 27570 16901
rect 27262 16890 27268 16892
rect 27324 16890 27348 16892
rect 27404 16890 27428 16892
rect 27484 16890 27508 16892
rect 27564 16890 27570 16892
rect 27324 16838 27326 16890
rect 27506 16838 27508 16890
rect 27262 16836 27268 16838
rect 27324 16836 27348 16838
rect 27404 16836 27428 16838
rect 27484 16836 27508 16838
rect 27564 16836 27570 16838
rect 27262 16827 27570 16836
rect 27262 15804 27570 15813
rect 27262 15802 27268 15804
rect 27324 15802 27348 15804
rect 27404 15802 27428 15804
rect 27484 15802 27508 15804
rect 27564 15802 27570 15804
rect 27324 15750 27326 15802
rect 27506 15750 27508 15802
rect 27262 15748 27268 15750
rect 27324 15748 27348 15750
rect 27404 15748 27428 15750
rect 27484 15748 27508 15750
rect 27564 15748 27570 15750
rect 27262 15739 27570 15748
rect 27262 14716 27570 14725
rect 27262 14714 27268 14716
rect 27324 14714 27348 14716
rect 27404 14714 27428 14716
rect 27484 14714 27508 14716
rect 27564 14714 27570 14716
rect 27324 14662 27326 14714
rect 27506 14662 27508 14714
rect 27262 14660 27268 14662
rect 27324 14660 27348 14662
rect 27404 14660 27428 14662
rect 27484 14660 27508 14662
rect 27564 14660 27570 14662
rect 27262 14651 27570 14660
rect 26238 13832 26294 13841
rect 25872 13806 25924 13812
rect 25884 13530 25912 13806
rect 26160 13790 26238 13818
rect 25872 13524 25924 13530
rect 25872 13466 25924 13472
rect 25780 13388 25832 13394
rect 25780 13330 25832 13336
rect 25792 13274 25820 13330
rect 25700 13246 25820 13274
rect 25884 13258 25912 13466
rect 25872 13252 25924 13258
rect 25318 12679 25374 12688
rect 25596 12708 25648 12714
rect 25596 12650 25648 12656
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25332 12442 25360 12582
rect 25410 12472 25466 12481
rect 25148 12406 25268 12434
rect 25320 12436 25372 12442
rect 25044 12368 25096 12374
rect 25044 12310 25096 12316
rect 25148 12306 25176 12406
rect 25608 12458 25636 12650
rect 25410 12407 25466 12416
rect 25516 12430 25636 12458
rect 25320 12378 25372 12384
rect 25136 12300 25188 12306
rect 25136 12242 25188 12248
rect 25148 11778 25176 12242
rect 25424 12102 25452 12407
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 25412 12096 25464 12102
rect 25412 12038 25464 12044
rect 25056 11750 25176 11778
rect 25056 11694 25084 11750
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 24860 11280 24912 11286
rect 24780 11240 24860 11268
rect 24124 11144 24176 11150
rect 24122 11112 24124 11121
rect 24216 11144 24268 11150
rect 24176 11112 24178 11121
rect 24216 11086 24268 11092
rect 24308 11144 24360 11150
rect 24308 11086 24360 11092
rect 24122 11047 24178 11056
rect 24228 11014 24256 11086
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 23904 10908 24212 10917
rect 23904 10906 23910 10908
rect 23966 10906 23990 10908
rect 24046 10906 24070 10908
rect 24126 10906 24150 10908
rect 24206 10906 24212 10908
rect 23966 10854 23968 10906
rect 24148 10854 24150 10906
rect 23904 10852 23910 10854
rect 23966 10852 23990 10854
rect 24046 10852 24070 10854
rect 24126 10852 24150 10854
rect 24206 10852 24212 10854
rect 23754 10840 23810 10849
rect 23904 10843 24212 10852
rect 23754 10775 23756 10784
rect 23808 10775 23810 10784
rect 23756 10746 23808 10752
rect 24124 10736 24176 10742
rect 24122 10704 24124 10713
rect 24176 10704 24178 10713
rect 24122 10639 24178 10648
rect 24780 10606 24808 11240
rect 24860 11222 24912 11228
rect 25056 11218 25084 11630
rect 25044 11212 25096 11218
rect 25044 11154 25096 11160
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 24032 10600 24084 10606
rect 24032 10542 24084 10548
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24768 10600 24820 10606
rect 24768 10542 24820 10548
rect 23664 9988 23716 9994
rect 23664 9930 23716 9936
rect 24044 9926 24072 10542
rect 24688 10266 24716 10542
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24308 10192 24360 10198
rect 24308 10134 24360 10140
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 23904 9820 24212 9829
rect 23904 9818 23910 9820
rect 23966 9818 23990 9820
rect 24046 9818 24070 9820
rect 24126 9818 24150 9820
rect 24206 9818 24212 9820
rect 23966 9766 23968 9818
rect 24148 9766 24150 9818
rect 23904 9764 23910 9766
rect 23966 9764 23990 9766
rect 24046 9764 24070 9766
rect 24126 9764 24150 9766
rect 24206 9764 24212 9766
rect 23904 9755 24212 9764
rect 24032 9512 24084 9518
rect 24084 9472 24164 9500
rect 24032 9454 24084 9460
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 24136 9330 24164 9472
rect 24320 9466 24348 10134
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24400 9580 24452 9586
rect 24400 9522 24452 9528
rect 24228 9450 24348 9466
rect 24216 9444 24348 9450
rect 24268 9438 24348 9444
rect 24216 9386 24268 9392
rect 24412 9330 24440 9522
rect 24492 9512 24544 9518
rect 24780 9466 24808 9862
rect 24872 9625 24900 9862
rect 24858 9616 24914 9625
rect 24858 9551 24914 9560
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 24860 9512 24912 9518
rect 24492 9454 24544 9460
rect 24596 9460 24860 9466
rect 24596 9454 24912 9460
rect 24044 8838 24072 9318
rect 24136 9302 24440 9330
rect 24504 9178 24532 9454
rect 24596 9438 24900 9454
rect 24596 9178 24624 9438
rect 24492 9172 24544 9178
rect 24492 9114 24544 9120
rect 24584 9172 24636 9178
rect 24584 9114 24636 9120
rect 24308 8968 24360 8974
rect 24308 8910 24360 8916
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 23904 8732 24212 8741
rect 23904 8730 23910 8732
rect 23966 8730 23990 8732
rect 24046 8730 24070 8732
rect 24126 8730 24150 8732
rect 24206 8730 24212 8732
rect 23966 8678 23968 8730
rect 24148 8678 24150 8730
rect 23904 8676 23910 8678
rect 23966 8676 23990 8678
rect 24046 8676 24070 8678
rect 24126 8676 24150 8678
rect 24206 8676 24212 8678
rect 23904 8667 24212 8676
rect 23664 8356 23716 8362
rect 23664 8298 23716 8304
rect 23676 8090 23704 8298
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23904 7644 24212 7653
rect 23904 7642 23910 7644
rect 23966 7642 23990 7644
rect 24046 7642 24070 7644
rect 24126 7642 24150 7644
rect 24206 7642 24212 7644
rect 23966 7590 23968 7642
rect 24148 7590 24150 7642
rect 23904 7588 23910 7590
rect 23966 7588 23990 7590
rect 24046 7588 24070 7590
rect 24126 7588 24150 7590
rect 24206 7588 24212 7590
rect 23904 7579 24212 7588
rect 24320 7206 24348 8910
rect 24492 8900 24544 8906
rect 24492 8842 24544 8848
rect 24504 8362 24532 8842
rect 24492 8356 24544 8362
rect 24492 8298 24544 8304
rect 24596 7342 24624 9114
rect 24964 9110 24992 9522
rect 24952 9104 25004 9110
rect 24952 9046 25004 9052
rect 25148 9042 25176 11154
rect 25240 10130 25268 12038
rect 25320 11620 25372 11626
rect 25320 11562 25372 11568
rect 25332 11354 25360 11562
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25516 10198 25544 12430
rect 25700 11218 25728 13246
rect 25872 13194 25924 13200
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25792 12782 25820 13126
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 25884 12646 25912 13194
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 26160 12345 26188 13790
rect 26238 13767 26294 13776
rect 27158 13832 27214 13841
rect 27158 13767 27214 13776
rect 27262 13628 27570 13637
rect 27262 13626 27268 13628
rect 27324 13626 27348 13628
rect 27404 13626 27428 13628
rect 27484 13626 27508 13628
rect 27564 13626 27570 13628
rect 27324 13574 27326 13626
rect 27506 13574 27508 13626
rect 27262 13572 27268 13574
rect 27324 13572 27348 13574
rect 27404 13572 27428 13574
rect 27484 13572 27508 13574
rect 27564 13572 27570 13574
rect 27262 13563 27570 13572
rect 26884 12640 26936 12646
rect 26884 12582 26936 12588
rect 26146 12336 26202 12345
rect 26146 12271 26202 12280
rect 26896 12238 26924 12582
rect 27262 12540 27570 12549
rect 27262 12538 27268 12540
rect 27324 12538 27348 12540
rect 27404 12538 27428 12540
rect 27484 12538 27508 12540
rect 27564 12538 27570 12540
rect 27324 12486 27326 12538
rect 27506 12486 27508 12538
rect 27262 12484 27268 12486
rect 27324 12484 27348 12486
rect 27404 12484 27428 12486
rect 27484 12484 27508 12486
rect 27564 12484 27570 12486
rect 27262 12475 27570 12484
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 27068 11892 27120 11898
rect 27068 11834 27120 11840
rect 26148 11552 26200 11558
rect 26148 11494 26200 11500
rect 26160 11218 26188 11494
rect 25688 11212 25740 11218
rect 25688 11154 25740 11160
rect 26148 11212 26200 11218
rect 26148 11154 26200 11160
rect 25596 11144 25648 11150
rect 25596 11086 25648 11092
rect 25608 10606 25636 11086
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25872 11008 25924 11014
rect 25872 10950 25924 10956
rect 26056 11008 26108 11014
rect 26056 10950 26108 10956
rect 25792 10742 25820 10950
rect 25780 10736 25832 10742
rect 25780 10678 25832 10684
rect 25884 10606 25912 10950
rect 25596 10600 25648 10606
rect 25596 10542 25648 10548
rect 25872 10600 25924 10606
rect 25872 10542 25924 10548
rect 25780 10464 25832 10470
rect 25780 10406 25832 10412
rect 25504 10192 25556 10198
rect 25504 10134 25556 10140
rect 25228 10124 25280 10130
rect 25228 10066 25280 10072
rect 25320 10124 25372 10130
rect 25320 10066 25372 10072
rect 25332 9625 25360 10066
rect 25792 9722 25820 10406
rect 26068 10266 26096 10950
rect 26056 10260 26108 10266
rect 26056 10202 26108 10208
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 25318 9616 25374 9625
rect 25318 9551 25374 9560
rect 25332 9518 25360 9551
rect 25792 9518 25820 9658
rect 26792 9580 26844 9586
rect 26792 9522 26844 9528
rect 25320 9512 25372 9518
rect 25240 9472 25320 9500
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 25136 9036 25188 9042
rect 25136 8978 25188 8984
rect 24872 8922 24900 8978
rect 24688 8894 24900 8922
rect 24688 8838 24716 8894
rect 24676 8832 24728 8838
rect 24676 8774 24728 8780
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24780 7818 24808 8774
rect 24872 7954 24900 8894
rect 25148 8566 25176 8978
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 24952 8356 25004 8362
rect 24952 8298 25004 8304
rect 24964 7954 24992 8298
rect 25148 8090 25176 8502
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 24952 7948 25004 7954
rect 24952 7890 25004 7896
rect 24768 7812 24820 7818
rect 24768 7754 24820 7760
rect 24780 7410 24808 7754
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 24308 7200 24360 7206
rect 24308 7142 24360 7148
rect 24584 7200 24636 7206
rect 24584 7142 24636 7148
rect 24596 6934 24624 7142
rect 24872 7002 24900 7890
rect 25044 7744 25096 7750
rect 25044 7686 25096 7692
rect 25056 7342 25084 7686
rect 25148 7342 25176 8026
rect 25240 7886 25268 9472
rect 25320 9454 25372 9460
rect 25780 9512 25832 9518
rect 25780 9454 25832 9460
rect 25320 9376 25372 9382
rect 25320 9318 25372 9324
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25332 9042 25360 9318
rect 25424 9042 25452 9318
rect 25792 9042 25820 9454
rect 25320 9036 25372 9042
rect 25320 8978 25372 8984
rect 25412 9036 25464 9042
rect 25412 8978 25464 8984
rect 25596 9036 25648 9042
rect 25596 8978 25648 8984
rect 25780 9036 25832 9042
rect 25780 8978 25832 8984
rect 25964 9036 26016 9042
rect 25964 8978 26016 8984
rect 25608 7954 25636 8978
rect 25976 8906 26004 8978
rect 26804 8974 26832 9522
rect 26792 8968 26844 8974
rect 26792 8910 26844 8916
rect 25964 8900 26016 8906
rect 25964 8842 26016 8848
rect 25780 8832 25832 8838
rect 25780 8774 25832 8780
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 25792 8430 25820 8774
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25596 7948 25648 7954
rect 25596 7890 25648 7896
rect 25228 7880 25280 7886
rect 25228 7822 25280 7828
rect 25608 7546 25636 7890
rect 25884 7750 25912 8774
rect 25976 7818 26004 8842
rect 26804 8294 26832 8910
rect 26792 8288 26844 8294
rect 26792 8230 26844 8236
rect 26804 7954 26832 8230
rect 26976 8016 27028 8022
rect 26976 7958 27028 7964
rect 26792 7948 26844 7954
rect 26792 7890 26844 7896
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 25964 7812 26016 7818
rect 25964 7754 26016 7760
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25872 7744 25924 7750
rect 25872 7686 25924 7692
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 25136 7336 25188 7342
rect 25136 7278 25188 7284
rect 24860 6996 24912 7002
rect 24860 6938 24912 6944
rect 24584 6928 24636 6934
rect 24584 6870 24636 6876
rect 25608 6866 25636 7482
rect 25596 6860 25648 6866
rect 25596 6802 25648 6808
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 23904 6556 24212 6565
rect 23904 6554 23910 6556
rect 23966 6554 23990 6556
rect 24046 6554 24070 6556
rect 24126 6554 24150 6556
rect 24206 6554 24212 6556
rect 23966 6502 23968 6554
rect 24148 6502 24150 6554
rect 23904 6500 23910 6502
rect 23966 6500 23990 6502
rect 24046 6500 24070 6502
rect 24126 6500 24150 6502
rect 24206 6500 24212 6502
rect 23904 6491 24212 6500
rect 24320 6322 24348 6734
rect 24308 6316 24360 6322
rect 24308 6258 24360 6264
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23492 5166 23520 6054
rect 24320 5846 24348 6258
rect 25700 6254 25728 7686
rect 25884 7478 25912 7686
rect 26068 7546 26096 7822
rect 26056 7540 26108 7546
rect 26056 7482 26108 7488
rect 25872 7472 25924 7478
rect 25872 7414 25924 7420
rect 25872 7336 25924 7342
rect 25872 7278 25924 7284
rect 26608 7336 26660 7342
rect 26608 7278 26660 7284
rect 25884 7002 25912 7278
rect 26620 7002 26648 7278
rect 25872 6996 25924 7002
rect 25872 6938 25924 6944
rect 26608 6996 26660 7002
rect 26608 6938 26660 6944
rect 26804 6798 26832 7890
rect 26988 6798 27016 7958
rect 26792 6792 26844 6798
rect 26792 6734 26844 6740
rect 26976 6792 27028 6798
rect 26976 6734 27028 6740
rect 26988 6458 27016 6734
rect 26976 6452 27028 6458
rect 26976 6394 27028 6400
rect 24400 6248 24452 6254
rect 24400 6190 24452 6196
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 24412 5914 24440 6190
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 23756 5840 23808 5846
rect 23756 5782 23808 5788
rect 24308 5840 24360 5846
rect 24308 5782 24360 5788
rect 24676 5840 24728 5846
rect 24676 5782 24728 5788
rect 23768 5302 23796 5782
rect 23904 5468 24212 5477
rect 23904 5466 23910 5468
rect 23966 5466 23990 5468
rect 24046 5466 24070 5468
rect 24126 5466 24150 5468
rect 24206 5466 24212 5468
rect 23966 5414 23968 5466
rect 24148 5414 24150 5466
rect 23904 5412 23910 5414
rect 23966 5412 23990 5414
rect 24046 5412 24070 5414
rect 24126 5412 24150 5414
rect 24206 5412 24212 5414
rect 23904 5403 24212 5412
rect 23756 5296 23808 5302
rect 23756 5238 23808 5244
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 23572 5092 23624 5098
rect 23572 5034 23624 5040
rect 23584 4622 23612 5034
rect 23768 4826 23796 5238
rect 24688 5166 24716 5782
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25424 5370 25452 5646
rect 25412 5364 25464 5370
rect 25412 5306 25464 5312
rect 24676 5160 24728 5166
rect 24676 5102 24728 5108
rect 25872 5160 25924 5166
rect 25872 5102 25924 5108
rect 25884 4826 25912 5102
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 25872 4820 25924 4826
rect 25872 4762 25924 4768
rect 23664 4684 23716 4690
rect 23664 4626 23716 4632
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23676 4146 23704 4626
rect 24308 4480 24360 4486
rect 24308 4422 24360 4428
rect 23904 4380 24212 4389
rect 23904 4378 23910 4380
rect 23966 4378 23990 4380
rect 24046 4378 24070 4380
rect 24126 4378 24150 4380
rect 24206 4378 24212 4380
rect 23966 4326 23968 4378
rect 24148 4326 24150 4378
rect 23904 4324 23910 4326
rect 23966 4324 23990 4326
rect 24046 4324 24070 4326
rect 24126 4324 24150 4326
rect 24206 4324 24212 4326
rect 23904 4315 24212 4324
rect 24122 4176 24178 4185
rect 23664 4140 23716 4146
rect 24122 4111 24178 4120
rect 23664 4082 23716 4088
rect 24136 4078 24164 4111
rect 24320 4078 24348 4422
rect 24124 4072 24176 4078
rect 23400 3998 23520 4026
rect 24124 4014 24176 4020
rect 24308 4072 24360 4078
rect 24308 4014 24360 4020
rect 25136 4072 25188 4078
rect 25136 4014 25188 4020
rect 25318 4040 25374 4049
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23400 3670 23428 3878
rect 23388 3664 23440 3670
rect 23388 3606 23440 3612
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 23124 3176 23152 3470
rect 23296 3188 23348 3194
rect 23124 3148 23296 3176
rect 23296 3130 23348 3136
rect 22836 2848 22888 2854
rect 22836 2790 22888 2796
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 22652 2644 22704 2650
rect 22572 2604 22652 2632
rect 22008 2508 22140 2514
rect 22060 2502 22140 2508
rect 22008 2450 22060 2456
rect 21836 2366 21956 2394
rect 21732 2304 21784 2310
rect 21732 2246 21784 2252
rect 21744 814 21772 2246
rect 20904 808 20956 814
rect 20904 750 20956 756
rect 21640 808 21692 814
rect 21640 750 21692 756
rect 21732 808 21784 814
rect 21732 750 21784 756
rect 20546 572 20854 581
rect 20546 570 20552 572
rect 20608 570 20632 572
rect 20688 570 20712 572
rect 20768 570 20792 572
rect 20848 570 20854 572
rect 20608 518 20610 570
rect 20790 518 20792 570
rect 20546 516 20552 518
rect 20608 516 20632 518
rect 20688 516 20712 518
rect 20768 516 20792 518
rect 20848 516 20854 518
rect 20546 507 20854 516
rect 21836 400 21864 2366
rect 22112 2310 22140 2502
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 22376 2508 22428 2514
rect 22376 2450 22428 2456
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22100 2304 22152 2310
rect 22100 2246 22152 2252
rect 22112 814 22140 2246
rect 22296 2106 22324 2450
rect 22284 2100 22336 2106
rect 22284 2042 22336 2048
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 22388 1970 22416 2042
rect 22192 1964 22244 1970
rect 22192 1906 22244 1912
rect 22376 1964 22428 1970
rect 22376 1906 22428 1912
rect 22204 1562 22232 1906
rect 22468 1760 22520 1766
rect 22468 1702 22520 1708
rect 22192 1556 22244 1562
rect 22192 1498 22244 1504
rect 22480 814 22508 1702
rect 22572 814 22600 2604
rect 22652 2586 22704 2592
rect 23020 2644 23072 2650
rect 23020 2586 23072 2592
rect 23032 2514 23060 2586
rect 23216 2514 23244 2790
rect 23020 2508 23072 2514
rect 23204 2508 23256 2514
rect 23020 2450 23072 2456
rect 23124 2468 23204 2496
rect 22652 2372 22704 2378
rect 22652 2314 22704 2320
rect 22664 814 22692 2314
rect 23032 2310 23060 2450
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 22836 1896 22888 1902
rect 22836 1838 22888 1844
rect 22848 1018 22876 1838
rect 23124 1766 23152 2468
rect 23204 2450 23256 2456
rect 23112 1760 23164 1766
rect 23112 1702 23164 1708
rect 22836 1012 22888 1018
rect 22836 954 22888 960
rect 22744 944 22796 950
rect 22744 886 22796 892
rect 22100 808 22152 814
rect 22100 750 22152 756
rect 22468 808 22520 814
rect 22468 750 22520 756
rect 22560 808 22612 814
rect 22560 750 22612 756
rect 22652 808 22704 814
rect 22652 750 22704 756
rect 22756 678 22784 886
rect 22928 808 22980 814
rect 23124 796 23152 1702
rect 23204 1420 23256 1426
rect 23204 1362 23256 1368
rect 23216 1018 23244 1362
rect 23204 1012 23256 1018
rect 23204 954 23256 960
rect 23308 950 23336 3130
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23400 2378 23428 2790
rect 23492 2774 23520 3998
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23492 2746 23612 2774
rect 23388 2372 23440 2378
rect 23388 2314 23440 2320
rect 23400 1902 23428 2314
rect 23388 1896 23440 1902
rect 23388 1838 23440 1844
rect 23480 1828 23532 1834
rect 23480 1770 23532 1776
rect 23492 1222 23520 1770
rect 23480 1216 23532 1222
rect 23480 1158 23532 1164
rect 23296 944 23348 950
rect 23296 886 23348 892
rect 23308 814 23336 886
rect 23492 814 23520 1158
rect 22980 768 23152 796
rect 23296 808 23348 814
rect 22928 750 22980 756
rect 23296 750 23348 756
rect 23480 808 23532 814
rect 23480 750 23532 756
rect 22744 672 22796 678
rect 22744 614 22796 620
rect 23584 400 23612 2746
rect 23768 2446 23796 3334
rect 23904 3292 24212 3301
rect 23904 3290 23910 3292
rect 23966 3290 23990 3292
rect 24046 3290 24070 3292
rect 24126 3290 24150 3292
rect 24206 3290 24212 3292
rect 23966 3238 23968 3290
rect 24148 3238 24150 3290
rect 23904 3236 23910 3238
rect 23966 3236 23990 3238
rect 24046 3236 24070 3238
rect 24126 3236 24150 3238
rect 24206 3236 24212 3238
rect 23904 3227 24212 3236
rect 24032 2984 24084 2990
rect 24412 2972 24440 3878
rect 24688 3670 24716 3878
rect 25148 3738 25176 4014
rect 25318 3975 25374 3984
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 24676 3664 24728 3670
rect 24676 3606 24728 3612
rect 24492 3596 24544 3602
rect 24492 3538 24544 3544
rect 24504 3194 24532 3538
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 24412 2944 24532 2972
rect 24032 2926 24084 2932
rect 24044 2650 24072 2926
rect 24504 2854 24532 2944
rect 25228 2916 25280 2922
rect 25228 2858 25280 2864
rect 24492 2848 24544 2854
rect 24492 2790 24544 2796
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23768 1290 23796 2382
rect 24308 2304 24360 2310
rect 24308 2246 24360 2252
rect 23904 2204 24212 2213
rect 23904 2202 23910 2204
rect 23966 2202 23990 2204
rect 24046 2202 24070 2204
rect 24126 2202 24150 2204
rect 24206 2202 24212 2204
rect 23966 2150 23968 2202
rect 24148 2150 24150 2202
rect 23904 2148 23910 2150
rect 23966 2148 23990 2150
rect 24046 2148 24070 2150
rect 24126 2148 24150 2150
rect 24206 2148 24212 2150
rect 23904 2139 24212 2148
rect 24320 2038 24348 2246
rect 24308 2032 24360 2038
rect 24308 1974 24360 1980
rect 24504 1902 24532 2790
rect 25240 2310 25268 2858
rect 25228 2304 25280 2310
rect 25228 2246 25280 2252
rect 25240 1902 25268 2246
rect 24492 1896 24544 1902
rect 24214 1864 24270 1873
rect 24492 1838 24544 1844
rect 24768 1896 24820 1902
rect 24768 1838 24820 1844
rect 25228 1896 25280 1902
rect 25228 1838 25280 1844
rect 24214 1799 24216 1808
rect 24268 1799 24270 1808
rect 24216 1770 24268 1776
rect 24780 1562 24808 1838
rect 24768 1556 24820 1562
rect 24768 1498 24820 1504
rect 23756 1284 23808 1290
rect 23756 1226 23808 1232
rect 23904 1116 24212 1125
rect 23904 1114 23910 1116
rect 23966 1114 23990 1116
rect 24046 1114 24070 1116
rect 24126 1114 24150 1116
rect 24206 1114 24212 1116
rect 23966 1062 23968 1114
rect 24148 1062 24150 1114
rect 23904 1060 23910 1062
rect 23966 1060 23990 1062
rect 24046 1060 24070 1062
rect 24126 1060 24150 1062
rect 24206 1060 24212 1062
rect 23904 1051 24212 1060
rect 24780 950 24808 1498
rect 24768 944 24820 950
rect 24768 886 24820 892
rect 25332 400 25360 3975
rect 25594 3768 25650 3777
rect 25650 3712 25728 3720
rect 25594 3703 25596 3712
rect 25648 3692 25728 3712
rect 25596 3674 25648 3680
rect 25596 3120 25648 3126
rect 25596 3062 25648 3068
rect 25608 1902 25636 3062
rect 25700 3058 25728 3692
rect 25688 3052 25740 3058
rect 25688 2994 25740 3000
rect 25688 2576 25740 2582
rect 25688 2518 25740 2524
rect 25700 1902 25728 2518
rect 25964 2440 26016 2446
rect 25964 2382 26016 2388
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25884 1902 25912 2246
rect 25976 2106 26004 2382
rect 25964 2100 26016 2106
rect 25964 2042 26016 2048
rect 25596 1896 25648 1902
rect 25596 1838 25648 1844
rect 25688 1896 25740 1902
rect 25688 1838 25740 1844
rect 25872 1896 25924 1902
rect 25872 1838 25924 1844
rect 25780 1760 25832 1766
rect 25780 1702 25832 1708
rect 26700 1760 26752 1766
rect 26700 1702 26752 1708
rect 25792 1018 25820 1702
rect 26712 1426 26740 1702
rect 26700 1420 26752 1426
rect 26700 1362 26752 1368
rect 25780 1012 25832 1018
rect 25780 954 25832 960
rect 27080 400 27108 11834
rect 27262 11452 27570 11461
rect 27262 11450 27268 11452
rect 27324 11450 27348 11452
rect 27404 11450 27428 11452
rect 27484 11450 27508 11452
rect 27564 11450 27570 11452
rect 27324 11398 27326 11450
rect 27506 11398 27508 11450
rect 27262 11396 27268 11398
rect 27324 11396 27348 11398
rect 27404 11396 27428 11398
rect 27484 11396 27508 11398
rect 27564 11396 27570 11398
rect 27262 11387 27570 11396
rect 27262 10364 27570 10373
rect 27262 10362 27268 10364
rect 27324 10362 27348 10364
rect 27404 10362 27428 10364
rect 27484 10362 27508 10364
rect 27564 10362 27570 10364
rect 27324 10310 27326 10362
rect 27506 10310 27508 10362
rect 27262 10308 27268 10310
rect 27324 10308 27348 10310
rect 27404 10308 27428 10310
rect 27484 10308 27508 10310
rect 27564 10308 27570 10310
rect 27262 10299 27570 10308
rect 27262 9276 27570 9285
rect 27262 9274 27268 9276
rect 27324 9274 27348 9276
rect 27404 9274 27428 9276
rect 27484 9274 27508 9276
rect 27564 9274 27570 9276
rect 27324 9222 27326 9274
rect 27506 9222 27508 9274
rect 27262 9220 27268 9222
rect 27324 9220 27348 9222
rect 27404 9220 27428 9222
rect 27484 9220 27508 9222
rect 27564 9220 27570 9222
rect 27262 9211 27570 9220
rect 27262 8188 27570 8197
rect 27262 8186 27268 8188
rect 27324 8186 27348 8188
rect 27404 8186 27428 8188
rect 27484 8186 27508 8188
rect 27564 8186 27570 8188
rect 27324 8134 27326 8186
rect 27506 8134 27508 8186
rect 27262 8132 27268 8134
rect 27324 8132 27348 8134
rect 27404 8132 27428 8134
rect 27484 8132 27508 8134
rect 27564 8132 27570 8134
rect 27262 8123 27570 8132
rect 27262 7100 27570 7109
rect 27262 7098 27268 7100
rect 27324 7098 27348 7100
rect 27404 7098 27428 7100
rect 27484 7098 27508 7100
rect 27564 7098 27570 7100
rect 27324 7046 27326 7098
rect 27506 7046 27508 7098
rect 27262 7044 27268 7046
rect 27324 7044 27348 7046
rect 27404 7044 27428 7046
rect 27484 7044 27508 7046
rect 27564 7044 27570 7046
rect 27262 7035 27570 7044
rect 27262 6012 27570 6021
rect 27262 6010 27268 6012
rect 27324 6010 27348 6012
rect 27404 6010 27428 6012
rect 27484 6010 27508 6012
rect 27564 6010 27570 6012
rect 27324 5958 27326 6010
rect 27506 5958 27508 6010
rect 27262 5956 27268 5958
rect 27324 5956 27348 5958
rect 27404 5956 27428 5958
rect 27484 5956 27508 5958
rect 27564 5956 27570 5958
rect 27262 5947 27570 5956
rect 27262 4924 27570 4933
rect 27262 4922 27268 4924
rect 27324 4922 27348 4924
rect 27404 4922 27428 4924
rect 27484 4922 27508 4924
rect 27564 4922 27570 4924
rect 27324 4870 27326 4922
rect 27506 4870 27508 4922
rect 27262 4868 27268 4870
rect 27324 4868 27348 4870
rect 27404 4868 27428 4870
rect 27484 4868 27508 4870
rect 27564 4868 27570 4870
rect 27262 4859 27570 4868
rect 27262 3836 27570 3845
rect 27262 3834 27268 3836
rect 27324 3834 27348 3836
rect 27404 3834 27428 3836
rect 27484 3834 27508 3836
rect 27564 3834 27570 3836
rect 27324 3782 27326 3834
rect 27506 3782 27508 3834
rect 27262 3780 27268 3782
rect 27324 3780 27348 3782
rect 27404 3780 27428 3782
rect 27484 3780 27508 3782
rect 27564 3780 27570 3782
rect 27262 3771 27570 3780
rect 27262 2748 27570 2757
rect 27262 2746 27268 2748
rect 27324 2746 27348 2748
rect 27404 2746 27428 2748
rect 27484 2746 27508 2748
rect 27564 2746 27570 2748
rect 27324 2694 27326 2746
rect 27506 2694 27508 2746
rect 27262 2692 27268 2694
rect 27324 2692 27348 2694
rect 27404 2692 27428 2694
rect 27484 2692 27508 2694
rect 27564 2692 27570 2694
rect 27262 2683 27570 2692
rect 27262 1660 27570 1669
rect 27262 1658 27268 1660
rect 27324 1658 27348 1660
rect 27404 1658 27428 1660
rect 27484 1658 27508 1660
rect 27564 1658 27570 1660
rect 27324 1606 27326 1658
rect 27506 1606 27508 1658
rect 27262 1604 27268 1606
rect 27324 1604 27348 1606
rect 27404 1604 27428 1606
rect 27484 1604 27508 1606
rect 27564 1604 27570 1606
rect 27262 1595 27570 1604
rect 27262 572 27570 581
rect 27262 570 27268 572
rect 27324 570 27348 572
rect 27404 570 27428 572
rect 27484 570 27508 572
rect 27564 570 27570 572
rect 27324 518 27326 570
rect 27506 518 27508 570
rect 27262 516 27268 518
rect 27324 516 27348 518
rect 27404 516 27428 518
rect 27484 516 27508 518
rect 27564 516 27570 518
rect 27262 507 27570 516
rect 11440 326 11836 354
rect 13082 0 13138 400
rect 14830 0 14886 400
rect 16578 0 16634 400
rect 18326 0 18382 400
rect 20074 0 20130 400
rect 21822 0 21878 400
rect 23570 0 23626 400
rect 25318 0 25374 400
rect 27066 0 27122 400
<< via2 >>
rect 3762 17434 3818 17436
rect 3842 17434 3898 17436
rect 3922 17434 3978 17436
rect 4002 17434 4058 17436
rect 3762 17382 3808 17434
rect 3808 17382 3818 17434
rect 3842 17382 3872 17434
rect 3872 17382 3884 17434
rect 3884 17382 3898 17434
rect 3922 17382 3936 17434
rect 3936 17382 3948 17434
rect 3948 17382 3978 17434
rect 4002 17382 4012 17434
rect 4012 17382 4058 17434
rect 3762 17380 3818 17382
rect 3842 17380 3898 17382
rect 3922 17380 3978 17382
rect 4002 17380 4058 17382
rect 7120 16890 7176 16892
rect 7200 16890 7256 16892
rect 7280 16890 7336 16892
rect 7360 16890 7416 16892
rect 7120 16838 7166 16890
rect 7166 16838 7176 16890
rect 7200 16838 7230 16890
rect 7230 16838 7242 16890
rect 7242 16838 7256 16890
rect 7280 16838 7294 16890
rect 7294 16838 7306 16890
rect 7306 16838 7336 16890
rect 7360 16838 7370 16890
rect 7370 16838 7416 16890
rect 7120 16836 7176 16838
rect 7200 16836 7256 16838
rect 7280 16836 7336 16838
rect 7360 16836 7416 16838
rect 3762 16346 3818 16348
rect 3842 16346 3898 16348
rect 3922 16346 3978 16348
rect 4002 16346 4058 16348
rect 3762 16294 3808 16346
rect 3808 16294 3818 16346
rect 3842 16294 3872 16346
rect 3872 16294 3884 16346
rect 3884 16294 3898 16346
rect 3922 16294 3936 16346
rect 3936 16294 3948 16346
rect 3948 16294 3978 16346
rect 4002 16294 4012 16346
rect 4012 16294 4058 16346
rect 3762 16292 3818 16294
rect 3842 16292 3898 16294
rect 3922 16292 3978 16294
rect 4002 16292 4058 16294
rect 3762 15258 3818 15260
rect 3842 15258 3898 15260
rect 3922 15258 3978 15260
rect 4002 15258 4058 15260
rect 3762 15206 3808 15258
rect 3808 15206 3818 15258
rect 3842 15206 3872 15258
rect 3872 15206 3884 15258
rect 3884 15206 3898 15258
rect 3922 15206 3936 15258
rect 3936 15206 3948 15258
rect 3948 15206 3978 15258
rect 4002 15206 4012 15258
rect 4012 15206 4058 15258
rect 3762 15204 3818 15206
rect 3842 15204 3898 15206
rect 3922 15204 3978 15206
rect 4002 15204 4058 15206
rect 4894 14864 4950 14920
rect 3762 14170 3818 14172
rect 3842 14170 3898 14172
rect 3922 14170 3978 14172
rect 4002 14170 4058 14172
rect 3762 14118 3808 14170
rect 3808 14118 3818 14170
rect 3842 14118 3872 14170
rect 3872 14118 3884 14170
rect 3884 14118 3898 14170
rect 3922 14118 3936 14170
rect 3936 14118 3948 14170
rect 3948 14118 3978 14170
rect 4002 14118 4012 14170
rect 4012 14118 4058 14170
rect 3762 14116 3818 14118
rect 3842 14116 3898 14118
rect 3922 14116 3978 14118
rect 4002 14116 4058 14118
rect 3762 13082 3818 13084
rect 3842 13082 3898 13084
rect 3922 13082 3978 13084
rect 4002 13082 4058 13084
rect 3762 13030 3808 13082
rect 3808 13030 3818 13082
rect 3842 13030 3872 13082
rect 3872 13030 3884 13082
rect 3884 13030 3898 13082
rect 3922 13030 3936 13082
rect 3936 13030 3948 13082
rect 3948 13030 3978 13082
rect 4002 13030 4012 13082
rect 4012 13030 4058 13082
rect 3762 13028 3818 13030
rect 3842 13028 3898 13030
rect 3922 13028 3978 13030
rect 4002 13028 4058 13030
rect 3762 11994 3818 11996
rect 3842 11994 3898 11996
rect 3922 11994 3978 11996
rect 4002 11994 4058 11996
rect 3762 11942 3808 11994
rect 3808 11942 3818 11994
rect 3842 11942 3872 11994
rect 3872 11942 3884 11994
rect 3884 11942 3898 11994
rect 3922 11942 3936 11994
rect 3936 11942 3948 11994
rect 3948 11942 3978 11994
rect 4002 11942 4012 11994
rect 4012 11942 4058 11994
rect 3762 11940 3818 11942
rect 3842 11940 3898 11942
rect 3922 11940 3978 11942
rect 4002 11940 4058 11942
rect 3762 10906 3818 10908
rect 3842 10906 3898 10908
rect 3922 10906 3978 10908
rect 4002 10906 4058 10908
rect 3762 10854 3808 10906
rect 3808 10854 3818 10906
rect 3842 10854 3872 10906
rect 3872 10854 3884 10906
rect 3884 10854 3898 10906
rect 3922 10854 3936 10906
rect 3936 10854 3948 10906
rect 3948 10854 3978 10906
rect 4002 10854 4012 10906
rect 4012 10854 4058 10906
rect 3762 10852 3818 10854
rect 3842 10852 3898 10854
rect 3922 10852 3978 10854
rect 4002 10852 4058 10854
rect 3762 9818 3818 9820
rect 3842 9818 3898 9820
rect 3922 9818 3978 9820
rect 4002 9818 4058 9820
rect 3762 9766 3808 9818
rect 3808 9766 3818 9818
rect 3842 9766 3872 9818
rect 3872 9766 3884 9818
rect 3884 9766 3898 9818
rect 3922 9766 3936 9818
rect 3936 9766 3948 9818
rect 3948 9766 3978 9818
rect 4002 9766 4012 9818
rect 4012 9766 4058 9818
rect 3762 9764 3818 9766
rect 3842 9764 3898 9766
rect 3922 9764 3978 9766
rect 4002 9764 4058 9766
rect 3762 8730 3818 8732
rect 3842 8730 3898 8732
rect 3922 8730 3978 8732
rect 4002 8730 4058 8732
rect 3762 8678 3808 8730
rect 3808 8678 3818 8730
rect 3842 8678 3872 8730
rect 3872 8678 3884 8730
rect 3884 8678 3898 8730
rect 3922 8678 3936 8730
rect 3936 8678 3948 8730
rect 3948 8678 3978 8730
rect 4002 8678 4012 8730
rect 4012 8678 4058 8730
rect 3762 8676 3818 8678
rect 3842 8676 3898 8678
rect 3922 8676 3978 8678
rect 4002 8676 4058 8678
rect 3762 7642 3818 7644
rect 3842 7642 3898 7644
rect 3922 7642 3978 7644
rect 4002 7642 4058 7644
rect 3762 7590 3808 7642
rect 3808 7590 3818 7642
rect 3842 7590 3872 7642
rect 3872 7590 3884 7642
rect 3884 7590 3898 7642
rect 3922 7590 3936 7642
rect 3936 7590 3948 7642
rect 3948 7590 3978 7642
rect 4002 7590 4012 7642
rect 4012 7590 4058 7642
rect 3762 7588 3818 7590
rect 3842 7588 3898 7590
rect 3922 7588 3978 7590
rect 4002 7588 4058 7590
rect 3762 6554 3818 6556
rect 3842 6554 3898 6556
rect 3922 6554 3978 6556
rect 4002 6554 4058 6556
rect 3762 6502 3808 6554
rect 3808 6502 3818 6554
rect 3842 6502 3872 6554
rect 3872 6502 3884 6554
rect 3884 6502 3898 6554
rect 3922 6502 3936 6554
rect 3936 6502 3948 6554
rect 3948 6502 3978 6554
rect 4002 6502 4012 6554
rect 4012 6502 4058 6554
rect 3762 6500 3818 6502
rect 3842 6500 3898 6502
rect 3922 6500 3978 6502
rect 4002 6500 4058 6502
rect 3762 5466 3818 5468
rect 3842 5466 3898 5468
rect 3922 5466 3978 5468
rect 4002 5466 4058 5468
rect 3762 5414 3808 5466
rect 3808 5414 3818 5466
rect 3842 5414 3872 5466
rect 3872 5414 3884 5466
rect 3884 5414 3898 5466
rect 3922 5414 3936 5466
rect 3936 5414 3948 5466
rect 3948 5414 3978 5466
rect 4002 5414 4012 5466
rect 4012 5414 4058 5466
rect 3762 5412 3818 5414
rect 3842 5412 3898 5414
rect 3922 5412 3978 5414
rect 4002 5412 4058 5414
rect 3762 4378 3818 4380
rect 3842 4378 3898 4380
rect 3922 4378 3978 4380
rect 4002 4378 4058 4380
rect 3762 4326 3808 4378
rect 3808 4326 3818 4378
rect 3842 4326 3872 4378
rect 3872 4326 3884 4378
rect 3884 4326 3898 4378
rect 3922 4326 3936 4378
rect 3936 4326 3948 4378
rect 3948 4326 3978 4378
rect 4002 4326 4012 4378
rect 4012 4326 4058 4378
rect 3762 4324 3818 4326
rect 3842 4324 3898 4326
rect 3922 4324 3978 4326
rect 4002 4324 4058 4326
rect 846 3440 902 3496
rect 3762 3290 3818 3292
rect 3842 3290 3898 3292
rect 3922 3290 3978 3292
rect 4002 3290 4058 3292
rect 3762 3238 3808 3290
rect 3808 3238 3818 3290
rect 3842 3238 3872 3290
rect 3872 3238 3884 3290
rect 3884 3238 3898 3290
rect 3922 3238 3936 3290
rect 3936 3238 3948 3290
rect 3948 3238 3978 3290
rect 4002 3238 4012 3290
rect 4012 3238 4058 3290
rect 3762 3236 3818 3238
rect 3842 3236 3898 3238
rect 3922 3236 3978 3238
rect 4002 3236 4058 3238
rect 3762 2202 3818 2204
rect 3842 2202 3898 2204
rect 3922 2202 3978 2204
rect 4002 2202 4058 2204
rect 3762 2150 3808 2202
rect 3808 2150 3818 2202
rect 3842 2150 3872 2202
rect 3872 2150 3884 2202
rect 3884 2150 3898 2202
rect 3922 2150 3936 2202
rect 3936 2150 3948 2202
rect 3948 2150 3978 2202
rect 4002 2150 4012 2202
rect 4012 2150 4058 2202
rect 3762 2148 3818 2150
rect 3842 2148 3898 2150
rect 3922 2148 3978 2150
rect 4002 2148 4058 2150
rect 3762 1114 3818 1116
rect 3842 1114 3898 1116
rect 3922 1114 3978 1116
rect 4002 1114 4058 1116
rect 3762 1062 3808 1114
rect 3808 1062 3818 1114
rect 3842 1062 3872 1114
rect 3872 1062 3884 1114
rect 3884 1062 3898 1114
rect 3922 1062 3936 1114
rect 3936 1062 3948 1114
rect 3948 1062 3978 1114
rect 4002 1062 4012 1114
rect 4012 1062 4058 1114
rect 3762 1060 3818 1062
rect 3842 1060 3898 1062
rect 3922 1060 3978 1062
rect 4002 1060 4058 1062
rect 5814 13912 5870 13968
rect 7120 15802 7176 15804
rect 7200 15802 7256 15804
rect 7280 15802 7336 15804
rect 7360 15802 7416 15804
rect 7120 15750 7166 15802
rect 7166 15750 7176 15802
rect 7200 15750 7230 15802
rect 7230 15750 7242 15802
rect 7242 15750 7256 15802
rect 7280 15750 7294 15802
rect 7294 15750 7306 15802
rect 7306 15750 7336 15802
rect 7360 15750 7370 15802
rect 7370 15750 7416 15802
rect 7120 15748 7176 15750
rect 7200 15748 7256 15750
rect 7280 15748 7336 15750
rect 7360 15748 7416 15750
rect 7120 14714 7176 14716
rect 7200 14714 7256 14716
rect 7280 14714 7336 14716
rect 7360 14714 7416 14716
rect 7120 14662 7166 14714
rect 7166 14662 7176 14714
rect 7200 14662 7230 14714
rect 7230 14662 7242 14714
rect 7242 14662 7256 14714
rect 7280 14662 7294 14714
rect 7294 14662 7306 14714
rect 7306 14662 7336 14714
rect 7360 14662 7370 14714
rect 7370 14662 7416 14714
rect 7120 14660 7176 14662
rect 7200 14660 7256 14662
rect 7280 14660 7336 14662
rect 7360 14660 7416 14662
rect 10478 17434 10534 17436
rect 10558 17434 10614 17436
rect 10638 17434 10694 17436
rect 10718 17434 10774 17436
rect 10478 17382 10524 17434
rect 10524 17382 10534 17434
rect 10558 17382 10588 17434
rect 10588 17382 10600 17434
rect 10600 17382 10614 17434
rect 10638 17382 10652 17434
rect 10652 17382 10664 17434
rect 10664 17382 10694 17434
rect 10718 17382 10728 17434
rect 10728 17382 10774 17434
rect 10478 17380 10534 17382
rect 10558 17380 10614 17382
rect 10638 17380 10694 17382
rect 10718 17380 10774 17382
rect 8482 15000 8538 15056
rect 8482 14864 8538 14920
rect 8022 13812 8024 13832
rect 8024 13812 8076 13832
rect 8076 13812 8078 13832
rect 8022 13776 8078 13812
rect 7120 13626 7176 13628
rect 7200 13626 7256 13628
rect 7280 13626 7336 13628
rect 7360 13626 7416 13628
rect 7120 13574 7166 13626
rect 7166 13574 7176 13626
rect 7200 13574 7230 13626
rect 7230 13574 7242 13626
rect 7242 13574 7256 13626
rect 7280 13574 7294 13626
rect 7294 13574 7306 13626
rect 7306 13574 7336 13626
rect 7360 13574 7370 13626
rect 7370 13574 7416 13626
rect 7120 13572 7176 13574
rect 7200 13572 7256 13574
rect 7280 13572 7336 13574
rect 7360 13572 7416 13574
rect 7120 12538 7176 12540
rect 7200 12538 7256 12540
rect 7280 12538 7336 12540
rect 7360 12538 7416 12540
rect 7120 12486 7166 12538
rect 7166 12486 7176 12538
rect 7200 12486 7230 12538
rect 7230 12486 7242 12538
rect 7242 12486 7256 12538
rect 7280 12486 7294 12538
rect 7294 12486 7306 12538
rect 7306 12486 7336 12538
rect 7360 12486 7370 12538
rect 7370 12486 7416 12538
rect 7120 12484 7176 12486
rect 7200 12484 7256 12486
rect 7280 12484 7336 12486
rect 7360 12484 7416 12486
rect 8206 12416 8262 12472
rect 7838 12300 7894 12336
rect 9126 13776 9182 13832
rect 7838 12280 7840 12300
rect 7840 12280 7892 12300
rect 7892 12280 7894 12300
rect 7470 11636 7472 11656
rect 7472 11636 7524 11656
rect 7524 11636 7526 11656
rect 7470 11600 7526 11636
rect 7120 11450 7176 11452
rect 7200 11450 7256 11452
rect 7280 11450 7336 11452
rect 7360 11450 7416 11452
rect 7120 11398 7166 11450
rect 7166 11398 7176 11450
rect 7200 11398 7230 11450
rect 7230 11398 7242 11450
rect 7242 11398 7256 11450
rect 7280 11398 7294 11450
rect 7294 11398 7306 11450
rect 7306 11398 7336 11450
rect 7360 11398 7370 11450
rect 7370 11398 7416 11450
rect 7120 11396 7176 11398
rect 7200 11396 7256 11398
rect 7280 11396 7336 11398
rect 7360 11396 7416 11398
rect 7120 10362 7176 10364
rect 7200 10362 7256 10364
rect 7280 10362 7336 10364
rect 7360 10362 7416 10364
rect 7120 10310 7166 10362
rect 7166 10310 7176 10362
rect 7200 10310 7230 10362
rect 7230 10310 7242 10362
rect 7242 10310 7256 10362
rect 7280 10310 7294 10362
rect 7294 10310 7306 10362
rect 7306 10310 7336 10362
rect 7360 10310 7370 10362
rect 7370 10310 7416 10362
rect 7120 10308 7176 10310
rect 7200 10308 7256 10310
rect 7280 10308 7336 10310
rect 7360 10308 7416 10310
rect 7120 9274 7176 9276
rect 7200 9274 7256 9276
rect 7280 9274 7336 9276
rect 7360 9274 7416 9276
rect 7120 9222 7166 9274
rect 7166 9222 7176 9274
rect 7200 9222 7230 9274
rect 7230 9222 7242 9274
rect 7242 9222 7256 9274
rect 7280 9222 7294 9274
rect 7294 9222 7306 9274
rect 7306 9222 7336 9274
rect 7360 9222 7370 9274
rect 7370 9222 7416 9274
rect 7120 9220 7176 9222
rect 7200 9220 7256 9222
rect 7280 9220 7336 9222
rect 7360 9220 7416 9222
rect 5814 8336 5870 8392
rect 7120 8186 7176 8188
rect 7200 8186 7256 8188
rect 7280 8186 7336 8188
rect 7360 8186 7416 8188
rect 7120 8134 7166 8186
rect 7166 8134 7176 8186
rect 7200 8134 7230 8186
rect 7230 8134 7242 8186
rect 7242 8134 7256 8186
rect 7280 8134 7294 8186
rect 7294 8134 7306 8186
rect 7306 8134 7336 8186
rect 7360 8134 7370 8186
rect 7370 8134 7416 8186
rect 7120 8132 7176 8134
rect 7200 8132 7256 8134
rect 7280 8132 7336 8134
rect 7360 8132 7416 8134
rect 7120 7098 7176 7100
rect 7200 7098 7256 7100
rect 7280 7098 7336 7100
rect 7360 7098 7416 7100
rect 7120 7046 7166 7098
rect 7166 7046 7176 7098
rect 7200 7046 7230 7098
rect 7230 7046 7242 7098
rect 7242 7046 7256 7098
rect 7280 7046 7294 7098
rect 7294 7046 7306 7098
rect 7306 7046 7336 7098
rect 7360 7046 7370 7098
rect 7370 7046 7416 7098
rect 7120 7044 7176 7046
rect 7200 7044 7256 7046
rect 7280 7044 7336 7046
rect 7360 7044 7416 7046
rect 6642 5636 6698 5672
rect 6642 5616 6644 5636
rect 6644 5616 6696 5636
rect 6696 5616 6698 5636
rect 7120 6010 7176 6012
rect 7200 6010 7256 6012
rect 7280 6010 7336 6012
rect 7360 6010 7416 6012
rect 7120 5958 7166 6010
rect 7166 5958 7176 6010
rect 7200 5958 7230 6010
rect 7230 5958 7242 6010
rect 7242 5958 7256 6010
rect 7280 5958 7294 6010
rect 7294 5958 7306 6010
rect 7306 5958 7336 6010
rect 7360 5958 7370 6010
rect 7370 5958 7416 6010
rect 7120 5956 7176 5958
rect 7200 5956 7256 5958
rect 7280 5956 7336 5958
rect 7360 5956 7416 5958
rect 7120 4922 7176 4924
rect 7200 4922 7256 4924
rect 7280 4922 7336 4924
rect 7360 4922 7416 4924
rect 7120 4870 7166 4922
rect 7166 4870 7176 4922
rect 7200 4870 7230 4922
rect 7230 4870 7242 4922
rect 7242 4870 7256 4922
rect 7280 4870 7294 4922
rect 7294 4870 7306 4922
rect 7306 4870 7336 4922
rect 7360 4870 7370 4922
rect 7370 4870 7416 4922
rect 7120 4868 7176 4870
rect 7200 4868 7256 4870
rect 7280 4868 7336 4870
rect 7360 4868 7416 4870
rect 7120 3834 7176 3836
rect 7200 3834 7256 3836
rect 7280 3834 7336 3836
rect 7360 3834 7416 3836
rect 7120 3782 7166 3834
rect 7166 3782 7176 3834
rect 7200 3782 7230 3834
rect 7230 3782 7242 3834
rect 7242 3782 7256 3834
rect 7280 3782 7294 3834
rect 7294 3782 7306 3834
rect 7306 3782 7336 3834
rect 7360 3782 7370 3834
rect 7370 3782 7416 3834
rect 7120 3780 7176 3782
rect 7200 3780 7256 3782
rect 7280 3780 7336 3782
rect 7360 3780 7416 3782
rect 7120 2746 7176 2748
rect 7200 2746 7256 2748
rect 7280 2746 7336 2748
rect 7360 2746 7416 2748
rect 7120 2694 7166 2746
rect 7166 2694 7176 2746
rect 7200 2694 7230 2746
rect 7230 2694 7242 2746
rect 7242 2694 7256 2746
rect 7280 2694 7294 2746
rect 7294 2694 7306 2746
rect 7306 2694 7336 2746
rect 7360 2694 7370 2746
rect 7370 2694 7416 2746
rect 7120 2692 7176 2694
rect 7200 2692 7256 2694
rect 7280 2692 7336 2694
rect 7360 2692 7416 2694
rect 7838 9424 7894 9480
rect 9586 13932 9642 13968
rect 9586 13912 9588 13932
rect 9588 13912 9640 13932
rect 9640 13912 9642 13932
rect 11242 16496 11298 16552
rect 10478 16346 10534 16348
rect 10558 16346 10614 16348
rect 10638 16346 10694 16348
rect 10718 16346 10774 16348
rect 10478 16294 10524 16346
rect 10524 16294 10534 16346
rect 10558 16294 10588 16346
rect 10588 16294 10600 16346
rect 10600 16294 10614 16346
rect 10638 16294 10652 16346
rect 10652 16294 10664 16346
rect 10664 16294 10694 16346
rect 10718 16294 10728 16346
rect 10728 16294 10774 16346
rect 10478 16292 10534 16294
rect 10558 16292 10614 16294
rect 10638 16292 10694 16294
rect 10718 16292 10774 16294
rect 10478 15258 10534 15260
rect 10558 15258 10614 15260
rect 10638 15258 10694 15260
rect 10718 15258 10774 15260
rect 10478 15206 10524 15258
rect 10524 15206 10534 15258
rect 10558 15206 10588 15258
rect 10588 15206 10600 15258
rect 10600 15206 10614 15258
rect 10638 15206 10652 15258
rect 10652 15206 10664 15258
rect 10664 15206 10694 15258
rect 10718 15206 10728 15258
rect 10728 15206 10774 15258
rect 10478 15204 10534 15206
rect 10558 15204 10614 15206
rect 10638 15204 10694 15206
rect 10718 15204 10774 15206
rect 8114 6296 8170 6352
rect 8850 7948 8906 7984
rect 8850 7928 8852 7948
rect 8852 7928 8904 7948
rect 8904 7928 8906 7948
rect 7120 1658 7176 1660
rect 7200 1658 7256 1660
rect 7280 1658 7336 1660
rect 7360 1658 7416 1660
rect 7120 1606 7166 1658
rect 7166 1606 7176 1658
rect 7200 1606 7230 1658
rect 7230 1606 7242 1658
rect 7242 1606 7256 1658
rect 7280 1606 7294 1658
rect 7294 1606 7306 1658
rect 7306 1606 7336 1658
rect 7360 1606 7370 1658
rect 7370 1606 7416 1658
rect 7120 1604 7176 1606
rect 7200 1604 7256 1606
rect 7280 1604 7336 1606
rect 7360 1604 7416 1606
rect 7120 570 7176 572
rect 7200 570 7256 572
rect 7280 570 7336 572
rect 7360 570 7416 572
rect 7120 518 7166 570
rect 7166 518 7176 570
rect 7200 518 7230 570
rect 7230 518 7242 570
rect 7242 518 7256 570
rect 7280 518 7294 570
rect 7294 518 7306 570
rect 7306 518 7336 570
rect 7360 518 7370 570
rect 7370 518 7416 570
rect 7120 516 7176 518
rect 7200 516 7256 518
rect 7280 516 7336 518
rect 7360 516 7416 518
rect 9678 11328 9734 11384
rect 10478 14170 10534 14172
rect 10558 14170 10614 14172
rect 10638 14170 10694 14172
rect 10718 14170 10774 14172
rect 10478 14118 10524 14170
rect 10524 14118 10534 14170
rect 10558 14118 10588 14170
rect 10588 14118 10600 14170
rect 10600 14118 10614 14170
rect 10638 14118 10652 14170
rect 10652 14118 10664 14170
rect 10664 14118 10694 14170
rect 10718 14118 10728 14170
rect 10728 14118 10774 14170
rect 10478 14116 10534 14118
rect 10558 14116 10614 14118
rect 10638 14116 10694 14118
rect 10718 14116 10774 14118
rect 10478 13082 10534 13084
rect 10558 13082 10614 13084
rect 10638 13082 10694 13084
rect 10718 13082 10774 13084
rect 10478 13030 10524 13082
rect 10524 13030 10534 13082
rect 10558 13030 10588 13082
rect 10588 13030 10600 13082
rect 10600 13030 10614 13082
rect 10638 13030 10652 13082
rect 10652 13030 10664 13082
rect 10664 13030 10694 13082
rect 10718 13030 10728 13082
rect 10728 13030 10774 13082
rect 10478 13028 10534 13030
rect 10558 13028 10614 13030
rect 10638 13028 10694 13030
rect 10718 13028 10774 13030
rect 10506 12824 10562 12880
rect 10874 12416 10930 12472
rect 10874 12144 10930 12200
rect 10478 11994 10534 11996
rect 10558 11994 10614 11996
rect 10638 11994 10694 11996
rect 10718 11994 10774 11996
rect 10478 11942 10524 11994
rect 10524 11942 10534 11994
rect 10558 11942 10588 11994
rect 10588 11942 10600 11994
rect 10600 11942 10614 11994
rect 10638 11942 10652 11994
rect 10652 11942 10664 11994
rect 10664 11942 10694 11994
rect 10718 11942 10728 11994
rect 10728 11942 10774 11994
rect 10478 11940 10534 11942
rect 10558 11940 10614 11942
rect 10638 11940 10694 11942
rect 10718 11940 10774 11942
rect 11058 11464 11114 11520
rect 10478 10906 10534 10908
rect 10558 10906 10614 10908
rect 10638 10906 10694 10908
rect 10718 10906 10774 10908
rect 10478 10854 10524 10906
rect 10524 10854 10534 10906
rect 10558 10854 10588 10906
rect 10588 10854 10600 10906
rect 10600 10854 10614 10906
rect 10638 10854 10652 10906
rect 10652 10854 10664 10906
rect 10664 10854 10694 10906
rect 10718 10854 10728 10906
rect 10728 10854 10774 10906
rect 10478 10852 10534 10854
rect 10558 10852 10614 10854
rect 10638 10852 10694 10854
rect 10718 10852 10774 10854
rect 10478 9818 10534 9820
rect 10558 9818 10614 9820
rect 10638 9818 10694 9820
rect 10718 9818 10774 9820
rect 10478 9766 10524 9818
rect 10524 9766 10534 9818
rect 10558 9766 10588 9818
rect 10588 9766 10600 9818
rect 10600 9766 10614 9818
rect 10638 9766 10652 9818
rect 10652 9766 10664 9818
rect 10664 9766 10694 9818
rect 10718 9766 10728 9818
rect 10728 9766 10774 9818
rect 10478 9764 10534 9766
rect 10558 9764 10614 9766
rect 10638 9764 10694 9766
rect 10718 9764 10774 9766
rect 10506 8900 10562 8936
rect 10506 8880 10508 8900
rect 10508 8880 10560 8900
rect 10560 8880 10562 8900
rect 10046 8472 10102 8528
rect 9862 6296 9918 6352
rect 10478 8730 10534 8732
rect 10558 8730 10614 8732
rect 10638 8730 10694 8732
rect 10718 8730 10774 8732
rect 10478 8678 10524 8730
rect 10524 8678 10534 8730
rect 10558 8678 10588 8730
rect 10588 8678 10600 8730
rect 10600 8678 10614 8730
rect 10638 8678 10652 8730
rect 10652 8678 10664 8730
rect 10664 8678 10694 8730
rect 10718 8678 10728 8730
rect 10728 8678 10774 8730
rect 10478 8676 10534 8678
rect 10558 8676 10614 8678
rect 10638 8676 10694 8678
rect 10718 8676 10774 8678
rect 10478 7642 10534 7644
rect 10558 7642 10614 7644
rect 10638 7642 10694 7644
rect 10718 7642 10774 7644
rect 10478 7590 10524 7642
rect 10524 7590 10534 7642
rect 10558 7590 10588 7642
rect 10588 7590 10600 7642
rect 10600 7590 10614 7642
rect 10638 7590 10652 7642
rect 10652 7590 10664 7642
rect 10664 7590 10694 7642
rect 10718 7590 10728 7642
rect 10728 7590 10774 7642
rect 10478 7588 10534 7590
rect 10558 7588 10614 7590
rect 10638 7588 10694 7590
rect 10718 7588 10774 7590
rect 10478 6554 10534 6556
rect 10558 6554 10614 6556
rect 10638 6554 10694 6556
rect 10718 6554 10774 6556
rect 10478 6502 10524 6554
rect 10524 6502 10534 6554
rect 10558 6502 10588 6554
rect 10588 6502 10600 6554
rect 10600 6502 10614 6554
rect 10638 6502 10652 6554
rect 10652 6502 10664 6554
rect 10664 6502 10694 6554
rect 10718 6502 10728 6554
rect 10728 6502 10774 6554
rect 10478 6500 10534 6502
rect 10558 6500 10614 6502
rect 10638 6500 10694 6502
rect 10718 6500 10774 6502
rect 9862 2896 9918 2952
rect 10478 5466 10534 5468
rect 10558 5466 10614 5468
rect 10638 5466 10694 5468
rect 10718 5466 10774 5468
rect 10478 5414 10524 5466
rect 10524 5414 10534 5466
rect 10558 5414 10588 5466
rect 10588 5414 10600 5466
rect 10600 5414 10614 5466
rect 10638 5414 10652 5466
rect 10652 5414 10664 5466
rect 10664 5414 10694 5466
rect 10718 5414 10728 5466
rect 10728 5414 10774 5466
rect 10478 5412 10534 5414
rect 10558 5412 10614 5414
rect 10638 5412 10694 5414
rect 10718 5412 10774 5414
rect 11886 15136 11942 15192
rect 13836 16890 13892 16892
rect 13916 16890 13972 16892
rect 13996 16890 14052 16892
rect 14076 16890 14132 16892
rect 13836 16838 13882 16890
rect 13882 16838 13892 16890
rect 13916 16838 13946 16890
rect 13946 16838 13958 16890
rect 13958 16838 13972 16890
rect 13996 16838 14010 16890
rect 14010 16838 14022 16890
rect 14022 16838 14052 16890
rect 14076 16838 14086 16890
rect 14086 16838 14132 16890
rect 13836 16836 13892 16838
rect 13916 16836 13972 16838
rect 13996 16836 14052 16838
rect 14076 16836 14132 16838
rect 12254 12688 12310 12744
rect 11702 11736 11758 11792
rect 11610 11464 11666 11520
rect 11610 11192 11666 11248
rect 11978 10548 11980 10568
rect 11980 10548 12032 10568
rect 12032 10548 12034 10568
rect 11978 10512 12034 10548
rect 13836 15802 13892 15804
rect 13916 15802 13972 15804
rect 13996 15802 14052 15804
rect 14076 15802 14132 15804
rect 13836 15750 13882 15802
rect 13882 15750 13892 15802
rect 13916 15750 13946 15802
rect 13946 15750 13958 15802
rect 13958 15750 13972 15802
rect 13996 15750 14010 15802
rect 14010 15750 14022 15802
rect 14022 15750 14052 15802
rect 14076 15750 14086 15802
rect 14086 15750 14132 15802
rect 13836 15748 13892 15750
rect 13916 15748 13972 15750
rect 13996 15748 14052 15750
rect 14076 15748 14132 15750
rect 13910 14884 13966 14920
rect 13910 14864 13912 14884
rect 13912 14864 13964 14884
rect 13964 14864 13966 14884
rect 13836 14714 13892 14716
rect 13916 14714 13972 14716
rect 13996 14714 14052 14716
rect 14076 14714 14132 14716
rect 13836 14662 13882 14714
rect 13882 14662 13892 14714
rect 13916 14662 13946 14714
rect 13946 14662 13958 14714
rect 13958 14662 13972 14714
rect 13996 14662 14010 14714
rect 14010 14662 14022 14714
rect 14022 14662 14052 14714
rect 14076 14662 14086 14714
rect 14086 14662 14132 14714
rect 13836 14660 13892 14662
rect 13916 14660 13972 14662
rect 13996 14660 14052 14662
rect 14076 14660 14132 14662
rect 17194 17434 17250 17436
rect 17274 17434 17330 17436
rect 17354 17434 17410 17436
rect 17434 17434 17490 17436
rect 17194 17382 17240 17434
rect 17240 17382 17250 17434
rect 17274 17382 17304 17434
rect 17304 17382 17316 17434
rect 17316 17382 17330 17434
rect 17354 17382 17368 17434
rect 17368 17382 17380 17434
rect 17380 17382 17410 17434
rect 17434 17382 17444 17434
rect 17444 17382 17490 17434
rect 17194 17380 17250 17382
rect 17274 17380 17330 17382
rect 17354 17380 17410 17382
rect 17434 17380 17490 17382
rect 15106 16496 15162 16552
rect 12622 13388 12678 13424
rect 12622 13368 12624 13388
rect 12624 13368 12676 13388
rect 12676 13368 12678 13388
rect 12530 12844 12586 12880
rect 12530 12824 12532 12844
rect 12532 12824 12584 12844
rect 12584 12824 12586 12844
rect 12070 9696 12126 9752
rect 11610 9424 11666 9480
rect 11518 8064 11574 8120
rect 12254 9016 12310 9072
rect 12714 10548 12716 10568
rect 12716 10548 12768 10568
rect 12768 10548 12770 10568
rect 12714 10512 12770 10548
rect 12346 8608 12402 8664
rect 12806 8608 12862 8664
rect 12254 6180 12310 6216
rect 12254 6160 12256 6180
rect 12256 6160 12308 6180
rect 12308 6160 12310 6180
rect 10478 4378 10534 4380
rect 10558 4378 10614 4380
rect 10638 4378 10694 4380
rect 10718 4378 10774 4380
rect 10478 4326 10524 4378
rect 10524 4326 10534 4378
rect 10558 4326 10588 4378
rect 10588 4326 10600 4378
rect 10600 4326 10614 4378
rect 10638 4326 10652 4378
rect 10652 4326 10664 4378
rect 10664 4326 10694 4378
rect 10718 4326 10728 4378
rect 10728 4326 10774 4378
rect 10478 4324 10534 4326
rect 10558 4324 10614 4326
rect 10638 4324 10694 4326
rect 10718 4324 10774 4326
rect 10478 3290 10534 3292
rect 10558 3290 10614 3292
rect 10638 3290 10694 3292
rect 10718 3290 10774 3292
rect 10478 3238 10524 3290
rect 10524 3238 10534 3290
rect 10558 3238 10588 3290
rect 10588 3238 10600 3290
rect 10600 3238 10614 3290
rect 10638 3238 10652 3290
rect 10652 3238 10664 3290
rect 10664 3238 10694 3290
rect 10718 3238 10728 3290
rect 10728 3238 10774 3290
rect 10478 3236 10534 3238
rect 10558 3236 10614 3238
rect 10638 3236 10694 3238
rect 10718 3236 10774 3238
rect 10478 2202 10534 2204
rect 10558 2202 10614 2204
rect 10638 2202 10694 2204
rect 10718 2202 10774 2204
rect 10478 2150 10524 2202
rect 10524 2150 10534 2202
rect 10558 2150 10588 2202
rect 10588 2150 10600 2202
rect 10600 2150 10614 2202
rect 10638 2150 10652 2202
rect 10652 2150 10664 2202
rect 10664 2150 10694 2202
rect 10718 2150 10728 2202
rect 10728 2150 10774 2202
rect 10478 2148 10534 2150
rect 10558 2148 10614 2150
rect 10638 2148 10694 2150
rect 10718 2148 10774 2150
rect 10478 1114 10534 1116
rect 10558 1114 10614 1116
rect 10638 1114 10694 1116
rect 10718 1114 10774 1116
rect 10478 1062 10524 1114
rect 10524 1062 10534 1114
rect 10558 1062 10588 1114
rect 10588 1062 10600 1114
rect 10600 1062 10614 1114
rect 10638 1062 10652 1114
rect 10652 1062 10664 1114
rect 10664 1062 10694 1114
rect 10718 1062 10728 1114
rect 10728 1062 10774 1114
rect 10478 1060 10534 1062
rect 10558 1060 10614 1062
rect 10638 1060 10694 1062
rect 10718 1060 10774 1062
rect 13836 13626 13892 13628
rect 13916 13626 13972 13628
rect 13996 13626 14052 13628
rect 14076 13626 14132 13628
rect 13836 13574 13882 13626
rect 13882 13574 13892 13626
rect 13916 13574 13946 13626
rect 13946 13574 13958 13626
rect 13958 13574 13972 13626
rect 13996 13574 14010 13626
rect 14010 13574 14022 13626
rect 14022 13574 14052 13626
rect 14076 13574 14086 13626
rect 14086 13574 14132 13626
rect 13836 13572 13892 13574
rect 13916 13572 13972 13574
rect 13996 13572 14052 13574
rect 14076 13572 14132 13574
rect 13836 12538 13892 12540
rect 13916 12538 13972 12540
rect 13996 12538 14052 12540
rect 14076 12538 14132 12540
rect 13836 12486 13882 12538
rect 13882 12486 13892 12538
rect 13916 12486 13946 12538
rect 13946 12486 13958 12538
rect 13958 12486 13972 12538
rect 13996 12486 14010 12538
rect 14010 12486 14022 12538
rect 14022 12486 14052 12538
rect 14076 12486 14086 12538
rect 14086 12486 14132 12538
rect 13836 12484 13892 12486
rect 13916 12484 13972 12486
rect 13996 12484 14052 12486
rect 14076 12484 14132 12486
rect 13836 11450 13892 11452
rect 13916 11450 13972 11452
rect 13996 11450 14052 11452
rect 14076 11450 14132 11452
rect 13836 11398 13882 11450
rect 13882 11398 13892 11450
rect 13916 11398 13946 11450
rect 13946 11398 13958 11450
rect 13958 11398 13972 11450
rect 13996 11398 14010 11450
rect 14010 11398 14022 11450
rect 14022 11398 14052 11450
rect 14076 11398 14086 11450
rect 14086 11398 14132 11450
rect 13836 11396 13892 11398
rect 13916 11396 13972 11398
rect 13996 11396 14052 11398
rect 14076 11396 14132 11398
rect 13634 11328 13690 11384
rect 13836 10362 13892 10364
rect 13916 10362 13972 10364
rect 13996 10362 14052 10364
rect 14076 10362 14132 10364
rect 13836 10310 13882 10362
rect 13882 10310 13892 10362
rect 13916 10310 13946 10362
rect 13946 10310 13958 10362
rect 13958 10310 13972 10362
rect 13996 10310 14010 10362
rect 14010 10310 14022 10362
rect 14022 10310 14052 10362
rect 14076 10310 14086 10362
rect 14086 10310 14132 10362
rect 13836 10308 13892 10310
rect 13916 10308 13972 10310
rect 13996 10308 14052 10310
rect 14076 10308 14132 10310
rect 14002 9580 14058 9616
rect 14002 9560 14004 9580
rect 14004 9560 14056 9580
rect 14056 9560 14058 9580
rect 13836 9274 13892 9276
rect 13916 9274 13972 9276
rect 13996 9274 14052 9276
rect 14076 9274 14132 9276
rect 13836 9222 13882 9274
rect 13882 9222 13892 9274
rect 13916 9222 13946 9274
rect 13946 9222 13958 9274
rect 13958 9222 13972 9274
rect 13996 9222 14010 9274
rect 14010 9222 14022 9274
rect 14022 9222 14052 9274
rect 14076 9222 14086 9274
rect 14086 9222 14132 9274
rect 13836 9220 13892 9222
rect 13916 9220 13972 9222
rect 13996 9220 14052 9222
rect 14076 9220 14132 9222
rect 13726 9016 13782 9072
rect 13450 8064 13506 8120
rect 13634 8064 13690 8120
rect 13818 8608 13874 8664
rect 13910 8472 13966 8528
rect 13836 8186 13892 8188
rect 13916 8186 13972 8188
rect 13996 8186 14052 8188
rect 14076 8186 14132 8188
rect 13836 8134 13882 8186
rect 13882 8134 13892 8186
rect 13916 8134 13946 8186
rect 13946 8134 13958 8186
rect 13958 8134 13972 8186
rect 13996 8134 14010 8186
rect 14010 8134 14022 8186
rect 14022 8134 14052 8186
rect 14076 8134 14086 8186
rect 14086 8134 14132 8186
rect 13836 8132 13892 8134
rect 13916 8132 13972 8134
rect 13996 8132 14052 8134
rect 14076 8132 14132 8134
rect 13836 7098 13892 7100
rect 13916 7098 13972 7100
rect 13996 7098 14052 7100
rect 14076 7098 14132 7100
rect 13836 7046 13882 7098
rect 13882 7046 13892 7098
rect 13916 7046 13946 7098
rect 13946 7046 13958 7098
rect 13958 7046 13972 7098
rect 13996 7046 14010 7098
rect 14010 7046 14022 7098
rect 14022 7046 14052 7098
rect 14076 7046 14086 7098
rect 14086 7046 14132 7098
rect 13836 7044 13892 7046
rect 13916 7044 13972 7046
rect 13996 7044 14052 7046
rect 14076 7044 14132 7046
rect 13836 6010 13892 6012
rect 13916 6010 13972 6012
rect 13996 6010 14052 6012
rect 14076 6010 14132 6012
rect 13836 5958 13882 6010
rect 13882 5958 13892 6010
rect 13916 5958 13946 6010
rect 13946 5958 13958 6010
rect 13958 5958 13972 6010
rect 13996 5958 14010 6010
rect 14010 5958 14022 6010
rect 14022 5958 14052 6010
rect 14076 5958 14086 6010
rect 14086 5958 14132 6010
rect 13836 5956 13892 5958
rect 13916 5956 13972 5958
rect 13996 5956 14052 5958
rect 14076 5956 14132 5958
rect 13836 4922 13892 4924
rect 13916 4922 13972 4924
rect 13996 4922 14052 4924
rect 14076 4922 14132 4924
rect 13836 4870 13882 4922
rect 13882 4870 13892 4922
rect 13916 4870 13946 4922
rect 13946 4870 13958 4922
rect 13958 4870 13972 4922
rect 13996 4870 14010 4922
rect 14010 4870 14022 4922
rect 14022 4870 14052 4922
rect 14076 4870 14086 4922
rect 14086 4870 14132 4922
rect 13836 4868 13892 4870
rect 13916 4868 13972 4870
rect 13996 4868 14052 4870
rect 14076 4868 14132 4870
rect 14462 5616 14518 5672
rect 15198 9696 15254 9752
rect 13836 3834 13892 3836
rect 13916 3834 13972 3836
rect 13996 3834 14052 3836
rect 14076 3834 14132 3836
rect 13836 3782 13882 3834
rect 13882 3782 13892 3834
rect 13916 3782 13946 3834
rect 13946 3782 13958 3834
rect 13958 3782 13972 3834
rect 13996 3782 14010 3834
rect 14010 3782 14022 3834
rect 14022 3782 14052 3834
rect 14076 3782 14086 3834
rect 14086 3782 14132 3834
rect 13836 3780 13892 3782
rect 13916 3780 13972 3782
rect 13996 3780 14052 3782
rect 14076 3780 14132 3782
rect 13358 2896 13414 2952
rect 13836 2746 13892 2748
rect 13916 2746 13972 2748
rect 13996 2746 14052 2748
rect 14076 2746 14132 2748
rect 13836 2694 13882 2746
rect 13882 2694 13892 2746
rect 13916 2694 13946 2746
rect 13946 2694 13958 2746
rect 13958 2694 13972 2746
rect 13996 2694 14010 2746
rect 14010 2694 14022 2746
rect 14022 2694 14052 2746
rect 14076 2694 14086 2746
rect 14086 2694 14132 2746
rect 13836 2692 13892 2694
rect 13916 2692 13972 2694
rect 13996 2692 14052 2694
rect 14076 2692 14132 2694
rect 13450 2488 13506 2544
rect 14094 2508 14150 2544
rect 14094 2488 14096 2508
rect 14096 2488 14148 2508
rect 14148 2488 14150 2508
rect 14830 3440 14886 3496
rect 13836 1658 13892 1660
rect 13916 1658 13972 1660
rect 13996 1658 14052 1660
rect 14076 1658 14132 1660
rect 13836 1606 13882 1658
rect 13882 1606 13892 1658
rect 13916 1606 13946 1658
rect 13946 1606 13958 1658
rect 13958 1606 13972 1658
rect 13996 1606 14010 1658
rect 14010 1606 14022 1658
rect 14022 1606 14052 1658
rect 14076 1606 14086 1658
rect 14086 1606 14132 1658
rect 13836 1604 13892 1606
rect 13916 1604 13972 1606
rect 13996 1604 14052 1606
rect 14076 1604 14132 1606
rect 17038 16496 17094 16552
rect 17194 16346 17250 16348
rect 17274 16346 17330 16348
rect 17354 16346 17410 16348
rect 17434 16346 17490 16348
rect 17194 16294 17240 16346
rect 17240 16294 17250 16346
rect 17274 16294 17304 16346
rect 17304 16294 17316 16346
rect 17316 16294 17330 16346
rect 17354 16294 17368 16346
rect 17368 16294 17380 16346
rect 17380 16294 17410 16346
rect 17434 16294 17444 16346
rect 17444 16294 17490 16346
rect 17194 16292 17250 16294
rect 17274 16292 17330 16294
rect 17354 16292 17410 16294
rect 17434 16292 17490 16294
rect 16762 15408 16818 15464
rect 16394 15136 16450 15192
rect 17194 15258 17250 15260
rect 17274 15258 17330 15260
rect 17354 15258 17410 15260
rect 17434 15258 17490 15260
rect 17194 15206 17240 15258
rect 17240 15206 17250 15258
rect 17274 15206 17304 15258
rect 17304 15206 17316 15258
rect 17316 15206 17330 15258
rect 17354 15206 17368 15258
rect 17368 15206 17380 15258
rect 17380 15206 17410 15258
rect 17434 15206 17444 15258
rect 17444 15206 17490 15258
rect 17194 15204 17250 15206
rect 17274 15204 17330 15206
rect 17354 15204 17410 15206
rect 17434 15204 17490 15206
rect 15750 9444 15806 9480
rect 15750 9424 15752 9444
rect 15752 9424 15804 9444
rect 15804 9424 15806 9444
rect 17194 14170 17250 14172
rect 17274 14170 17330 14172
rect 17354 14170 17410 14172
rect 17434 14170 17490 14172
rect 17194 14118 17240 14170
rect 17240 14118 17250 14170
rect 17274 14118 17304 14170
rect 17304 14118 17316 14170
rect 17316 14118 17330 14170
rect 17354 14118 17368 14170
rect 17368 14118 17380 14170
rect 17380 14118 17410 14170
rect 17434 14118 17444 14170
rect 17444 14118 17490 14170
rect 17194 14116 17250 14118
rect 17274 14116 17330 14118
rect 17354 14116 17410 14118
rect 17434 14116 17490 14118
rect 17194 13082 17250 13084
rect 17274 13082 17330 13084
rect 17354 13082 17410 13084
rect 17434 13082 17490 13084
rect 17194 13030 17240 13082
rect 17240 13030 17250 13082
rect 17274 13030 17304 13082
rect 17304 13030 17316 13082
rect 17316 13030 17330 13082
rect 17354 13030 17368 13082
rect 17368 13030 17380 13082
rect 17380 13030 17410 13082
rect 17434 13030 17444 13082
rect 17444 13030 17490 13082
rect 17194 13028 17250 13030
rect 17274 13028 17330 13030
rect 17354 13028 17410 13030
rect 17434 13028 17490 13030
rect 18142 13368 18198 13424
rect 18142 12708 18198 12744
rect 18142 12688 18144 12708
rect 18144 12688 18196 12708
rect 18196 12688 18198 12708
rect 18050 12552 18106 12608
rect 17194 11994 17250 11996
rect 17274 11994 17330 11996
rect 17354 11994 17410 11996
rect 17434 11994 17490 11996
rect 17194 11942 17240 11994
rect 17240 11942 17250 11994
rect 17274 11942 17304 11994
rect 17304 11942 17316 11994
rect 17316 11942 17330 11994
rect 17354 11942 17368 11994
rect 17368 11942 17380 11994
rect 17380 11942 17410 11994
rect 17434 11942 17444 11994
rect 17444 11942 17490 11994
rect 17194 11940 17250 11942
rect 17274 11940 17330 11942
rect 17354 11940 17410 11942
rect 17434 11940 17490 11942
rect 17590 11872 17646 11928
rect 17590 11736 17646 11792
rect 17194 10906 17250 10908
rect 17274 10906 17330 10908
rect 17354 10906 17410 10908
rect 17434 10906 17490 10908
rect 17194 10854 17240 10906
rect 17240 10854 17250 10906
rect 17274 10854 17304 10906
rect 17304 10854 17316 10906
rect 17316 10854 17330 10906
rect 17354 10854 17368 10906
rect 17368 10854 17380 10906
rect 17380 10854 17410 10906
rect 17434 10854 17444 10906
rect 17444 10854 17490 10906
rect 17194 10852 17250 10854
rect 17274 10852 17330 10854
rect 17354 10852 17410 10854
rect 17434 10852 17490 10854
rect 16578 9288 16634 9344
rect 16854 9036 16910 9072
rect 16854 9016 16856 9036
rect 16856 9016 16908 9036
rect 16908 9016 16910 9036
rect 16670 7928 16726 7984
rect 17194 9818 17250 9820
rect 17274 9818 17330 9820
rect 17354 9818 17410 9820
rect 17434 9818 17490 9820
rect 17194 9766 17240 9818
rect 17240 9766 17250 9818
rect 17274 9766 17304 9818
rect 17304 9766 17316 9818
rect 17316 9766 17330 9818
rect 17354 9766 17368 9818
rect 17368 9766 17380 9818
rect 17380 9766 17410 9818
rect 17434 9766 17444 9818
rect 17444 9766 17490 9818
rect 17194 9764 17250 9766
rect 17274 9764 17330 9766
rect 17354 9764 17410 9766
rect 17434 9764 17490 9766
rect 17130 9288 17186 9344
rect 17194 8730 17250 8732
rect 17274 8730 17330 8732
rect 17354 8730 17410 8732
rect 17434 8730 17490 8732
rect 17194 8678 17240 8730
rect 17240 8678 17250 8730
rect 17274 8678 17304 8730
rect 17304 8678 17316 8730
rect 17316 8678 17330 8730
rect 17354 8678 17368 8730
rect 17368 8678 17380 8730
rect 17380 8678 17410 8730
rect 17434 8678 17444 8730
rect 17444 8678 17490 8730
rect 17194 8676 17250 8678
rect 17274 8676 17330 8678
rect 17354 8676 17410 8678
rect 17434 8676 17490 8678
rect 17774 9288 17830 9344
rect 17194 7642 17250 7644
rect 17274 7642 17330 7644
rect 17354 7642 17410 7644
rect 17434 7642 17490 7644
rect 17194 7590 17240 7642
rect 17240 7590 17250 7642
rect 17274 7590 17304 7642
rect 17304 7590 17316 7642
rect 17316 7590 17330 7642
rect 17354 7590 17368 7642
rect 17368 7590 17380 7642
rect 17380 7590 17410 7642
rect 17434 7590 17444 7642
rect 17444 7590 17490 7642
rect 17194 7588 17250 7590
rect 17274 7588 17330 7590
rect 17354 7588 17410 7590
rect 17434 7588 17490 7590
rect 17682 8472 17738 8528
rect 17194 6554 17250 6556
rect 17274 6554 17330 6556
rect 17354 6554 17410 6556
rect 17434 6554 17490 6556
rect 17194 6502 17240 6554
rect 17240 6502 17250 6554
rect 17274 6502 17304 6554
rect 17304 6502 17316 6554
rect 17316 6502 17330 6554
rect 17354 6502 17368 6554
rect 17368 6502 17380 6554
rect 17380 6502 17410 6554
rect 17434 6502 17444 6554
rect 17444 6502 17490 6554
rect 17194 6500 17250 6502
rect 17274 6500 17330 6502
rect 17354 6500 17410 6502
rect 17434 6500 17490 6502
rect 17194 5466 17250 5468
rect 17274 5466 17330 5468
rect 17354 5466 17410 5468
rect 17434 5466 17490 5468
rect 17194 5414 17240 5466
rect 17240 5414 17250 5466
rect 17274 5414 17304 5466
rect 17304 5414 17316 5466
rect 17316 5414 17330 5466
rect 17354 5414 17368 5466
rect 17368 5414 17380 5466
rect 17380 5414 17410 5466
rect 17434 5414 17444 5466
rect 17444 5414 17490 5466
rect 17194 5412 17250 5414
rect 17274 5412 17330 5414
rect 17354 5412 17410 5414
rect 17434 5412 17490 5414
rect 17222 4684 17278 4720
rect 17222 4664 17224 4684
rect 17224 4664 17276 4684
rect 17276 4664 17278 4684
rect 17194 4378 17250 4380
rect 17274 4378 17330 4380
rect 17354 4378 17410 4380
rect 17434 4378 17490 4380
rect 17194 4326 17240 4378
rect 17240 4326 17250 4378
rect 17274 4326 17304 4378
rect 17304 4326 17316 4378
rect 17316 4326 17330 4378
rect 17354 4326 17368 4378
rect 17368 4326 17380 4378
rect 17380 4326 17410 4378
rect 17434 4326 17444 4378
rect 17444 4326 17490 4378
rect 17194 4324 17250 4326
rect 17274 4324 17330 4326
rect 17354 4324 17410 4326
rect 17434 4324 17490 4326
rect 13836 570 13892 572
rect 13916 570 13972 572
rect 13996 570 14052 572
rect 14076 570 14132 572
rect 13836 518 13882 570
rect 13882 518 13892 570
rect 13916 518 13946 570
rect 13946 518 13958 570
rect 13958 518 13972 570
rect 13996 518 14010 570
rect 14010 518 14022 570
rect 14022 518 14052 570
rect 14076 518 14086 570
rect 14086 518 14132 570
rect 13836 516 13892 518
rect 13916 516 13972 518
rect 13996 516 14052 518
rect 14076 516 14132 518
rect 18142 4664 18198 4720
rect 17194 3290 17250 3292
rect 17274 3290 17330 3292
rect 17354 3290 17410 3292
rect 17434 3290 17490 3292
rect 17194 3238 17240 3290
rect 17240 3238 17250 3290
rect 17274 3238 17304 3290
rect 17304 3238 17316 3290
rect 17316 3238 17330 3290
rect 17354 3238 17368 3290
rect 17368 3238 17380 3290
rect 17380 3238 17410 3290
rect 17434 3238 17444 3290
rect 17444 3238 17490 3290
rect 17194 3236 17250 3238
rect 17274 3236 17330 3238
rect 17354 3236 17410 3238
rect 17434 3236 17490 3238
rect 17194 2202 17250 2204
rect 17274 2202 17330 2204
rect 17354 2202 17410 2204
rect 17434 2202 17490 2204
rect 17194 2150 17240 2202
rect 17240 2150 17250 2202
rect 17274 2150 17304 2202
rect 17304 2150 17316 2202
rect 17316 2150 17330 2202
rect 17354 2150 17368 2202
rect 17368 2150 17380 2202
rect 17380 2150 17410 2202
rect 17434 2150 17444 2202
rect 17444 2150 17490 2202
rect 17194 2148 17250 2150
rect 17274 2148 17330 2150
rect 17354 2148 17410 2150
rect 17434 2148 17490 2150
rect 18510 11600 18566 11656
rect 18694 11464 18750 11520
rect 18418 11056 18474 11112
rect 18602 10784 18658 10840
rect 19430 14320 19486 14376
rect 20552 16890 20608 16892
rect 20632 16890 20688 16892
rect 20712 16890 20768 16892
rect 20792 16890 20848 16892
rect 20552 16838 20598 16890
rect 20598 16838 20608 16890
rect 20632 16838 20662 16890
rect 20662 16838 20674 16890
rect 20674 16838 20688 16890
rect 20712 16838 20726 16890
rect 20726 16838 20738 16890
rect 20738 16838 20768 16890
rect 20792 16838 20802 16890
rect 20802 16838 20848 16890
rect 20552 16836 20608 16838
rect 20632 16836 20688 16838
rect 20712 16836 20768 16838
rect 20792 16836 20848 16838
rect 20552 15802 20608 15804
rect 20632 15802 20688 15804
rect 20712 15802 20768 15804
rect 20792 15802 20848 15804
rect 20552 15750 20598 15802
rect 20598 15750 20608 15802
rect 20632 15750 20662 15802
rect 20662 15750 20674 15802
rect 20674 15750 20688 15802
rect 20712 15750 20726 15802
rect 20726 15750 20738 15802
rect 20738 15750 20768 15802
rect 20792 15750 20802 15802
rect 20802 15750 20848 15802
rect 20552 15748 20608 15750
rect 20632 15748 20688 15750
rect 20712 15748 20768 15750
rect 20792 15748 20848 15750
rect 20552 14714 20608 14716
rect 20632 14714 20688 14716
rect 20712 14714 20768 14716
rect 20792 14714 20848 14716
rect 20552 14662 20598 14714
rect 20598 14662 20608 14714
rect 20632 14662 20662 14714
rect 20662 14662 20674 14714
rect 20674 14662 20688 14714
rect 20712 14662 20726 14714
rect 20726 14662 20738 14714
rect 20738 14662 20768 14714
rect 20792 14662 20802 14714
rect 20802 14662 20848 14714
rect 20552 14660 20608 14662
rect 20632 14660 20688 14662
rect 20712 14660 20768 14662
rect 20792 14660 20848 14662
rect 20552 13626 20608 13628
rect 20632 13626 20688 13628
rect 20712 13626 20768 13628
rect 20792 13626 20848 13628
rect 20552 13574 20598 13626
rect 20598 13574 20608 13626
rect 20632 13574 20662 13626
rect 20662 13574 20674 13626
rect 20674 13574 20688 13626
rect 20712 13574 20726 13626
rect 20726 13574 20738 13626
rect 20738 13574 20768 13626
rect 20792 13574 20802 13626
rect 20802 13574 20848 13626
rect 20552 13572 20608 13574
rect 20632 13572 20688 13574
rect 20712 13572 20768 13574
rect 20792 13572 20848 13574
rect 20552 12538 20608 12540
rect 20632 12538 20688 12540
rect 20712 12538 20768 12540
rect 20792 12538 20848 12540
rect 20552 12486 20598 12538
rect 20598 12486 20608 12538
rect 20632 12486 20662 12538
rect 20662 12486 20674 12538
rect 20674 12486 20688 12538
rect 20712 12486 20726 12538
rect 20726 12486 20738 12538
rect 20738 12486 20768 12538
rect 20792 12486 20802 12538
rect 20802 12486 20848 12538
rect 20552 12484 20608 12486
rect 20632 12484 20688 12486
rect 20712 12484 20768 12486
rect 20792 12484 20848 12486
rect 19430 6296 19486 6352
rect 21086 12280 21142 12336
rect 20552 11450 20608 11452
rect 20632 11450 20688 11452
rect 20712 11450 20768 11452
rect 20792 11450 20848 11452
rect 20552 11398 20598 11450
rect 20598 11398 20608 11450
rect 20632 11398 20662 11450
rect 20662 11398 20674 11450
rect 20674 11398 20688 11450
rect 20712 11398 20726 11450
rect 20726 11398 20738 11450
rect 20738 11398 20768 11450
rect 20792 11398 20802 11450
rect 20802 11398 20848 11450
rect 20552 11396 20608 11398
rect 20632 11396 20688 11398
rect 20712 11396 20768 11398
rect 20792 11396 20848 11398
rect 22374 13776 22430 13832
rect 21546 11600 21602 11656
rect 21362 11192 21418 11248
rect 20534 10648 20590 10704
rect 20552 10362 20608 10364
rect 20632 10362 20688 10364
rect 20712 10362 20768 10364
rect 20792 10362 20848 10364
rect 20552 10310 20598 10362
rect 20598 10310 20608 10362
rect 20632 10310 20662 10362
rect 20662 10310 20674 10362
rect 20674 10310 20688 10362
rect 20712 10310 20726 10362
rect 20726 10310 20738 10362
rect 20738 10310 20768 10362
rect 20792 10310 20802 10362
rect 20802 10310 20848 10362
rect 20552 10308 20608 10310
rect 20632 10308 20688 10310
rect 20712 10308 20768 10310
rect 20792 10308 20848 10310
rect 20902 9560 20958 9616
rect 20552 9274 20608 9276
rect 20632 9274 20688 9276
rect 20712 9274 20768 9276
rect 20792 9274 20848 9276
rect 20552 9222 20598 9274
rect 20598 9222 20608 9274
rect 20632 9222 20662 9274
rect 20662 9222 20674 9274
rect 20674 9222 20688 9274
rect 20712 9222 20726 9274
rect 20726 9222 20738 9274
rect 20738 9222 20768 9274
rect 20792 9222 20802 9274
rect 20802 9222 20848 9274
rect 20552 9220 20608 9222
rect 20632 9220 20688 9222
rect 20712 9220 20768 9222
rect 20792 9220 20848 9222
rect 20552 8186 20608 8188
rect 20632 8186 20688 8188
rect 20712 8186 20768 8188
rect 20792 8186 20848 8188
rect 20552 8134 20598 8186
rect 20598 8134 20608 8186
rect 20632 8134 20662 8186
rect 20662 8134 20674 8186
rect 20674 8134 20688 8186
rect 20712 8134 20726 8186
rect 20726 8134 20738 8186
rect 20738 8134 20768 8186
rect 20792 8134 20802 8186
rect 20802 8134 20848 8186
rect 20552 8132 20608 8134
rect 20632 8132 20688 8134
rect 20712 8132 20768 8134
rect 20792 8132 20848 8134
rect 21178 8880 21234 8936
rect 20552 7098 20608 7100
rect 20632 7098 20688 7100
rect 20712 7098 20768 7100
rect 20792 7098 20848 7100
rect 20552 7046 20598 7098
rect 20598 7046 20608 7098
rect 20632 7046 20662 7098
rect 20662 7046 20674 7098
rect 20674 7046 20688 7098
rect 20712 7046 20726 7098
rect 20726 7046 20738 7098
rect 20738 7046 20768 7098
rect 20792 7046 20802 7098
rect 20802 7046 20848 7098
rect 20552 7044 20608 7046
rect 20632 7044 20688 7046
rect 20712 7044 20768 7046
rect 20792 7044 20848 7046
rect 20552 6010 20608 6012
rect 20632 6010 20688 6012
rect 20712 6010 20768 6012
rect 20792 6010 20848 6012
rect 20552 5958 20598 6010
rect 20598 5958 20608 6010
rect 20632 5958 20662 6010
rect 20662 5958 20674 6010
rect 20674 5958 20688 6010
rect 20712 5958 20726 6010
rect 20726 5958 20738 6010
rect 20738 5958 20768 6010
rect 20792 5958 20802 6010
rect 20802 5958 20848 6010
rect 20552 5956 20608 5958
rect 20632 5956 20688 5958
rect 20712 5956 20768 5958
rect 20792 5956 20848 5958
rect 19430 5208 19486 5264
rect 18326 3984 18382 4040
rect 18234 2896 18290 2952
rect 17682 1808 17738 1864
rect 17194 1114 17250 1116
rect 17274 1114 17330 1116
rect 17354 1114 17410 1116
rect 17434 1114 17490 1116
rect 17194 1062 17240 1114
rect 17240 1062 17250 1114
rect 17274 1062 17304 1114
rect 17304 1062 17316 1114
rect 17316 1062 17330 1114
rect 17354 1062 17368 1114
rect 17368 1062 17380 1114
rect 17380 1062 17410 1114
rect 17434 1062 17444 1114
rect 17444 1062 17490 1114
rect 17194 1060 17250 1062
rect 17274 1060 17330 1062
rect 17354 1060 17410 1062
rect 17434 1060 17490 1062
rect 20074 4120 20130 4176
rect 18418 1980 18420 2000
rect 18420 1980 18472 2000
rect 18472 1980 18474 2000
rect 18418 1944 18474 1980
rect 21086 5208 21142 5264
rect 21546 5908 21602 5944
rect 21546 5888 21548 5908
rect 21548 5888 21600 5908
rect 21600 5888 21602 5908
rect 20552 4922 20608 4924
rect 20632 4922 20688 4924
rect 20712 4922 20768 4924
rect 20792 4922 20848 4924
rect 20552 4870 20598 4922
rect 20598 4870 20608 4922
rect 20632 4870 20662 4922
rect 20662 4870 20674 4922
rect 20674 4870 20688 4922
rect 20712 4870 20726 4922
rect 20726 4870 20738 4922
rect 20738 4870 20768 4922
rect 20792 4870 20802 4922
rect 20802 4870 20848 4922
rect 20552 4868 20608 4870
rect 20632 4868 20688 4870
rect 20712 4868 20768 4870
rect 20792 4868 20848 4870
rect 20552 3834 20608 3836
rect 20632 3834 20688 3836
rect 20712 3834 20768 3836
rect 20792 3834 20848 3836
rect 20552 3782 20598 3834
rect 20598 3782 20608 3834
rect 20632 3782 20662 3834
rect 20662 3782 20674 3834
rect 20674 3782 20688 3834
rect 20712 3782 20726 3834
rect 20726 3782 20738 3834
rect 20738 3782 20768 3834
rect 20792 3782 20802 3834
rect 20802 3782 20848 3834
rect 20552 3780 20608 3782
rect 20632 3780 20688 3782
rect 20712 3780 20768 3782
rect 20792 3780 20848 3782
rect 20552 2746 20608 2748
rect 20632 2746 20688 2748
rect 20712 2746 20768 2748
rect 20792 2746 20848 2748
rect 19062 1944 19118 2000
rect 20552 2694 20598 2746
rect 20598 2694 20608 2746
rect 20632 2694 20662 2746
rect 20662 2694 20674 2746
rect 20674 2694 20688 2746
rect 20712 2694 20726 2746
rect 20726 2694 20738 2746
rect 20738 2694 20768 2746
rect 20792 2694 20802 2746
rect 20802 2694 20848 2746
rect 20552 2692 20608 2694
rect 20632 2692 20688 2694
rect 20712 2692 20768 2694
rect 20792 2692 20848 2694
rect 20552 1658 20608 1660
rect 20632 1658 20688 1660
rect 20712 1658 20768 1660
rect 20792 1658 20848 1660
rect 20552 1606 20598 1658
rect 20598 1606 20608 1658
rect 20632 1606 20662 1658
rect 20662 1606 20674 1658
rect 20674 1606 20688 1658
rect 20712 1606 20726 1658
rect 20726 1606 20738 1658
rect 20738 1606 20768 1658
rect 20792 1606 20802 1658
rect 20802 1606 20848 1658
rect 20552 1604 20608 1606
rect 20632 1604 20688 1606
rect 20712 1604 20768 1606
rect 20792 1604 20848 1606
rect 23910 17434 23966 17436
rect 23990 17434 24046 17436
rect 24070 17434 24126 17436
rect 24150 17434 24206 17436
rect 23910 17382 23956 17434
rect 23956 17382 23966 17434
rect 23990 17382 24020 17434
rect 24020 17382 24032 17434
rect 24032 17382 24046 17434
rect 24070 17382 24084 17434
rect 24084 17382 24096 17434
rect 24096 17382 24126 17434
rect 24150 17382 24160 17434
rect 24160 17382 24206 17434
rect 23910 17380 23966 17382
rect 23990 17380 24046 17382
rect 24070 17380 24126 17382
rect 24150 17380 24206 17382
rect 23478 15000 23534 15056
rect 23478 14320 23534 14376
rect 23910 16346 23966 16348
rect 23990 16346 24046 16348
rect 24070 16346 24126 16348
rect 24150 16346 24206 16348
rect 23910 16294 23956 16346
rect 23956 16294 23966 16346
rect 23990 16294 24020 16346
rect 24020 16294 24032 16346
rect 24032 16294 24046 16346
rect 24070 16294 24084 16346
rect 24084 16294 24096 16346
rect 24096 16294 24126 16346
rect 24150 16294 24160 16346
rect 24160 16294 24206 16346
rect 23910 16292 23966 16294
rect 23990 16292 24046 16294
rect 24070 16292 24126 16294
rect 24150 16292 24206 16294
rect 23910 15258 23966 15260
rect 23990 15258 24046 15260
rect 24070 15258 24126 15260
rect 24150 15258 24206 15260
rect 23910 15206 23956 15258
rect 23956 15206 23966 15258
rect 23990 15206 24020 15258
rect 24020 15206 24032 15258
rect 24032 15206 24046 15258
rect 24070 15206 24084 15258
rect 24084 15206 24096 15258
rect 24096 15206 24126 15258
rect 24150 15206 24160 15258
rect 24160 15206 24206 15258
rect 23910 15204 23966 15206
rect 23990 15204 24046 15206
rect 24070 15204 24126 15206
rect 24150 15204 24206 15206
rect 23910 14170 23966 14172
rect 23990 14170 24046 14172
rect 24070 14170 24126 14172
rect 24150 14170 24206 14172
rect 23910 14118 23956 14170
rect 23956 14118 23966 14170
rect 23990 14118 24020 14170
rect 24020 14118 24032 14170
rect 24032 14118 24046 14170
rect 24070 14118 24084 14170
rect 24084 14118 24096 14170
rect 24096 14118 24126 14170
rect 24150 14118 24160 14170
rect 24160 14118 24206 14170
rect 23910 14116 23966 14118
rect 23990 14116 24046 14118
rect 24070 14116 24126 14118
rect 24150 14116 24206 14118
rect 23910 13082 23966 13084
rect 23990 13082 24046 13084
rect 24070 13082 24126 13084
rect 24150 13082 24206 13084
rect 23910 13030 23956 13082
rect 23956 13030 23966 13082
rect 23990 13030 24020 13082
rect 24020 13030 24032 13082
rect 24032 13030 24046 13082
rect 24070 13030 24084 13082
rect 24084 13030 24096 13082
rect 24096 13030 24126 13082
rect 24150 13030 24160 13082
rect 24160 13030 24206 13082
rect 23910 13028 23966 13030
rect 23990 13028 24046 13030
rect 24070 13028 24126 13030
rect 24150 13028 24206 13030
rect 22558 11600 22614 11656
rect 22558 11056 22614 11112
rect 22374 5888 22430 5944
rect 22558 3712 22614 3768
rect 23910 11994 23966 11996
rect 23990 11994 24046 11996
rect 24070 11994 24126 11996
rect 24150 11994 24206 11996
rect 23910 11942 23956 11994
rect 23956 11942 23966 11994
rect 23990 11942 24020 11994
rect 24020 11942 24032 11994
rect 24032 11942 24046 11994
rect 24070 11942 24084 11994
rect 24084 11942 24096 11994
rect 24096 11942 24126 11994
rect 24150 11942 24160 11994
rect 24160 11942 24206 11994
rect 23910 11940 23966 11942
rect 23990 11940 24046 11942
rect 24070 11940 24126 11942
rect 24150 11940 24206 11942
rect 24582 12144 24638 12200
rect 25318 12688 25374 12744
rect 27268 16890 27324 16892
rect 27348 16890 27404 16892
rect 27428 16890 27484 16892
rect 27508 16890 27564 16892
rect 27268 16838 27314 16890
rect 27314 16838 27324 16890
rect 27348 16838 27378 16890
rect 27378 16838 27390 16890
rect 27390 16838 27404 16890
rect 27428 16838 27442 16890
rect 27442 16838 27454 16890
rect 27454 16838 27484 16890
rect 27508 16838 27518 16890
rect 27518 16838 27564 16890
rect 27268 16836 27324 16838
rect 27348 16836 27404 16838
rect 27428 16836 27484 16838
rect 27508 16836 27564 16838
rect 27268 15802 27324 15804
rect 27348 15802 27404 15804
rect 27428 15802 27484 15804
rect 27508 15802 27564 15804
rect 27268 15750 27314 15802
rect 27314 15750 27324 15802
rect 27348 15750 27378 15802
rect 27378 15750 27390 15802
rect 27390 15750 27404 15802
rect 27428 15750 27442 15802
rect 27442 15750 27454 15802
rect 27454 15750 27484 15802
rect 27508 15750 27518 15802
rect 27518 15750 27564 15802
rect 27268 15748 27324 15750
rect 27348 15748 27404 15750
rect 27428 15748 27484 15750
rect 27508 15748 27564 15750
rect 27268 14714 27324 14716
rect 27348 14714 27404 14716
rect 27428 14714 27484 14716
rect 27508 14714 27564 14716
rect 27268 14662 27314 14714
rect 27314 14662 27324 14714
rect 27348 14662 27378 14714
rect 27378 14662 27390 14714
rect 27390 14662 27404 14714
rect 27428 14662 27442 14714
rect 27442 14662 27454 14714
rect 27454 14662 27484 14714
rect 27508 14662 27518 14714
rect 27518 14662 27564 14714
rect 27268 14660 27324 14662
rect 27348 14660 27404 14662
rect 27428 14660 27484 14662
rect 27508 14660 27564 14662
rect 25410 12416 25466 12472
rect 24122 11092 24124 11112
rect 24124 11092 24176 11112
rect 24176 11092 24178 11112
rect 24122 11056 24178 11092
rect 23910 10906 23966 10908
rect 23990 10906 24046 10908
rect 24070 10906 24126 10908
rect 24150 10906 24206 10908
rect 23910 10854 23956 10906
rect 23956 10854 23966 10906
rect 23990 10854 24020 10906
rect 24020 10854 24032 10906
rect 24032 10854 24046 10906
rect 24070 10854 24084 10906
rect 24084 10854 24096 10906
rect 24096 10854 24126 10906
rect 24150 10854 24160 10906
rect 24160 10854 24206 10906
rect 23910 10852 23966 10854
rect 23990 10852 24046 10854
rect 24070 10852 24126 10854
rect 24150 10852 24206 10854
rect 23754 10804 23810 10840
rect 23754 10784 23756 10804
rect 23756 10784 23808 10804
rect 23808 10784 23810 10804
rect 24122 10684 24124 10704
rect 24124 10684 24176 10704
rect 24176 10684 24178 10704
rect 24122 10648 24178 10684
rect 23910 9818 23966 9820
rect 23990 9818 24046 9820
rect 24070 9818 24126 9820
rect 24150 9818 24206 9820
rect 23910 9766 23956 9818
rect 23956 9766 23966 9818
rect 23990 9766 24020 9818
rect 24020 9766 24032 9818
rect 24032 9766 24046 9818
rect 24070 9766 24084 9818
rect 24084 9766 24096 9818
rect 24096 9766 24126 9818
rect 24150 9766 24160 9818
rect 24160 9766 24206 9818
rect 23910 9764 23966 9766
rect 23990 9764 24046 9766
rect 24070 9764 24126 9766
rect 24150 9764 24206 9766
rect 24858 9560 24914 9616
rect 23910 8730 23966 8732
rect 23990 8730 24046 8732
rect 24070 8730 24126 8732
rect 24150 8730 24206 8732
rect 23910 8678 23956 8730
rect 23956 8678 23966 8730
rect 23990 8678 24020 8730
rect 24020 8678 24032 8730
rect 24032 8678 24046 8730
rect 24070 8678 24084 8730
rect 24084 8678 24096 8730
rect 24096 8678 24126 8730
rect 24150 8678 24160 8730
rect 24160 8678 24206 8730
rect 23910 8676 23966 8678
rect 23990 8676 24046 8678
rect 24070 8676 24126 8678
rect 24150 8676 24206 8678
rect 23910 7642 23966 7644
rect 23990 7642 24046 7644
rect 24070 7642 24126 7644
rect 24150 7642 24206 7644
rect 23910 7590 23956 7642
rect 23956 7590 23966 7642
rect 23990 7590 24020 7642
rect 24020 7590 24032 7642
rect 24032 7590 24046 7642
rect 24070 7590 24084 7642
rect 24084 7590 24096 7642
rect 24096 7590 24126 7642
rect 24150 7590 24160 7642
rect 24160 7590 24206 7642
rect 23910 7588 23966 7590
rect 23990 7588 24046 7590
rect 24070 7588 24126 7590
rect 24150 7588 24206 7590
rect 26238 13776 26294 13832
rect 27158 13776 27214 13832
rect 27268 13626 27324 13628
rect 27348 13626 27404 13628
rect 27428 13626 27484 13628
rect 27508 13626 27564 13628
rect 27268 13574 27314 13626
rect 27314 13574 27324 13626
rect 27348 13574 27378 13626
rect 27378 13574 27390 13626
rect 27390 13574 27404 13626
rect 27428 13574 27442 13626
rect 27442 13574 27454 13626
rect 27454 13574 27484 13626
rect 27508 13574 27518 13626
rect 27518 13574 27564 13626
rect 27268 13572 27324 13574
rect 27348 13572 27404 13574
rect 27428 13572 27484 13574
rect 27508 13572 27564 13574
rect 26146 12280 26202 12336
rect 27268 12538 27324 12540
rect 27348 12538 27404 12540
rect 27428 12538 27484 12540
rect 27508 12538 27564 12540
rect 27268 12486 27314 12538
rect 27314 12486 27324 12538
rect 27348 12486 27378 12538
rect 27378 12486 27390 12538
rect 27390 12486 27404 12538
rect 27428 12486 27442 12538
rect 27442 12486 27454 12538
rect 27454 12486 27484 12538
rect 27508 12486 27518 12538
rect 27518 12486 27564 12538
rect 27268 12484 27324 12486
rect 27348 12484 27404 12486
rect 27428 12484 27484 12486
rect 27508 12484 27564 12486
rect 25318 9560 25374 9616
rect 23910 6554 23966 6556
rect 23990 6554 24046 6556
rect 24070 6554 24126 6556
rect 24150 6554 24206 6556
rect 23910 6502 23956 6554
rect 23956 6502 23966 6554
rect 23990 6502 24020 6554
rect 24020 6502 24032 6554
rect 24032 6502 24046 6554
rect 24070 6502 24084 6554
rect 24084 6502 24096 6554
rect 24096 6502 24126 6554
rect 24150 6502 24160 6554
rect 24160 6502 24206 6554
rect 23910 6500 23966 6502
rect 23990 6500 24046 6502
rect 24070 6500 24126 6502
rect 24150 6500 24206 6502
rect 23910 5466 23966 5468
rect 23990 5466 24046 5468
rect 24070 5466 24126 5468
rect 24150 5466 24206 5468
rect 23910 5414 23956 5466
rect 23956 5414 23966 5466
rect 23990 5414 24020 5466
rect 24020 5414 24032 5466
rect 24032 5414 24046 5466
rect 24070 5414 24084 5466
rect 24084 5414 24096 5466
rect 24096 5414 24126 5466
rect 24150 5414 24160 5466
rect 24160 5414 24206 5466
rect 23910 5412 23966 5414
rect 23990 5412 24046 5414
rect 24070 5412 24126 5414
rect 24150 5412 24206 5414
rect 23910 4378 23966 4380
rect 23990 4378 24046 4380
rect 24070 4378 24126 4380
rect 24150 4378 24206 4380
rect 23910 4326 23956 4378
rect 23956 4326 23966 4378
rect 23990 4326 24020 4378
rect 24020 4326 24032 4378
rect 24032 4326 24046 4378
rect 24070 4326 24084 4378
rect 24084 4326 24096 4378
rect 24096 4326 24126 4378
rect 24150 4326 24160 4378
rect 24160 4326 24206 4378
rect 23910 4324 23966 4326
rect 23990 4324 24046 4326
rect 24070 4324 24126 4326
rect 24150 4324 24206 4326
rect 24122 4120 24178 4176
rect 20552 570 20608 572
rect 20632 570 20688 572
rect 20712 570 20768 572
rect 20792 570 20848 572
rect 20552 518 20598 570
rect 20598 518 20608 570
rect 20632 518 20662 570
rect 20662 518 20674 570
rect 20674 518 20688 570
rect 20712 518 20726 570
rect 20726 518 20738 570
rect 20738 518 20768 570
rect 20792 518 20802 570
rect 20802 518 20848 570
rect 20552 516 20608 518
rect 20632 516 20688 518
rect 20712 516 20768 518
rect 20792 516 20848 518
rect 23910 3290 23966 3292
rect 23990 3290 24046 3292
rect 24070 3290 24126 3292
rect 24150 3290 24206 3292
rect 23910 3238 23956 3290
rect 23956 3238 23966 3290
rect 23990 3238 24020 3290
rect 24020 3238 24032 3290
rect 24032 3238 24046 3290
rect 24070 3238 24084 3290
rect 24084 3238 24096 3290
rect 24096 3238 24126 3290
rect 24150 3238 24160 3290
rect 24160 3238 24206 3290
rect 23910 3236 23966 3238
rect 23990 3236 24046 3238
rect 24070 3236 24126 3238
rect 24150 3236 24206 3238
rect 25318 3984 25374 4040
rect 23910 2202 23966 2204
rect 23990 2202 24046 2204
rect 24070 2202 24126 2204
rect 24150 2202 24206 2204
rect 23910 2150 23956 2202
rect 23956 2150 23966 2202
rect 23990 2150 24020 2202
rect 24020 2150 24032 2202
rect 24032 2150 24046 2202
rect 24070 2150 24084 2202
rect 24084 2150 24096 2202
rect 24096 2150 24126 2202
rect 24150 2150 24160 2202
rect 24160 2150 24206 2202
rect 23910 2148 23966 2150
rect 23990 2148 24046 2150
rect 24070 2148 24126 2150
rect 24150 2148 24206 2150
rect 24214 1828 24270 1864
rect 24214 1808 24216 1828
rect 24216 1808 24268 1828
rect 24268 1808 24270 1828
rect 23910 1114 23966 1116
rect 23990 1114 24046 1116
rect 24070 1114 24126 1116
rect 24150 1114 24206 1116
rect 23910 1062 23956 1114
rect 23956 1062 23966 1114
rect 23990 1062 24020 1114
rect 24020 1062 24032 1114
rect 24032 1062 24046 1114
rect 24070 1062 24084 1114
rect 24084 1062 24096 1114
rect 24096 1062 24126 1114
rect 24150 1062 24160 1114
rect 24160 1062 24206 1114
rect 23910 1060 23966 1062
rect 23990 1060 24046 1062
rect 24070 1060 24126 1062
rect 24150 1060 24206 1062
rect 25594 3732 25650 3768
rect 25594 3712 25596 3732
rect 25596 3712 25648 3732
rect 25648 3712 25650 3732
rect 27268 11450 27324 11452
rect 27348 11450 27404 11452
rect 27428 11450 27484 11452
rect 27508 11450 27564 11452
rect 27268 11398 27314 11450
rect 27314 11398 27324 11450
rect 27348 11398 27378 11450
rect 27378 11398 27390 11450
rect 27390 11398 27404 11450
rect 27428 11398 27442 11450
rect 27442 11398 27454 11450
rect 27454 11398 27484 11450
rect 27508 11398 27518 11450
rect 27518 11398 27564 11450
rect 27268 11396 27324 11398
rect 27348 11396 27404 11398
rect 27428 11396 27484 11398
rect 27508 11396 27564 11398
rect 27268 10362 27324 10364
rect 27348 10362 27404 10364
rect 27428 10362 27484 10364
rect 27508 10362 27564 10364
rect 27268 10310 27314 10362
rect 27314 10310 27324 10362
rect 27348 10310 27378 10362
rect 27378 10310 27390 10362
rect 27390 10310 27404 10362
rect 27428 10310 27442 10362
rect 27442 10310 27454 10362
rect 27454 10310 27484 10362
rect 27508 10310 27518 10362
rect 27518 10310 27564 10362
rect 27268 10308 27324 10310
rect 27348 10308 27404 10310
rect 27428 10308 27484 10310
rect 27508 10308 27564 10310
rect 27268 9274 27324 9276
rect 27348 9274 27404 9276
rect 27428 9274 27484 9276
rect 27508 9274 27564 9276
rect 27268 9222 27314 9274
rect 27314 9222 27324 9274
rect 27348 9222 27378 9274
rect 27378 9222 27390 9274
rect 27390 9222 27404 9274
rect 27428 9222 27442 9274
rect 27442 9222 27454 9274
rect 27454 9222 27484 9274
rect 27508 9222 27518 9274
rect 27518 9222 27564 9274
rect 27268 9220 27324 9222
rect 27348 9220 27404 9222
rect 27428 9220 27484 9222
rect 27508 9220 27564 9222
rect 27268 8186 27324 8188
rect 27348 8186 27404 8188
rect 27428 8186 27484 8188
rect 27508 8186 27564 8188
rect 27268 8134 27314 8186
rect 27314 8134 27324 8186
rect 27348 8134 27378 8186
rect 27378 8134 27390 8186
rect 27390 8134 27404 8186
rect 27428 8134 27442 8186
rect 27442 8134 27454 8186
rect 27454 8134 27484 8186
rect 27508 8134 27518 8186
rect 27518 8134 27564 8186
rect 27268 8132 27324 8134
rect 27348 8132 27404 8134
rect 27428 8132 27484 8134
rect 27508 8132 27564 8134
rect 27268 7098 27324 7100
rect 27348 7098 27404 7100
rect 27428 7098 27484 7100
rect 27508 7098 27564 7100
rect 27268 7046 27314 7098
rect 27314 7046 27324 7098
rect 27348 7046 27378 7098
rect 27378 7046 27390 7098
rect 27390 7046 27404 7098
rect 27428 7046 27442 7098
rect 27442 7046 27454 7098
rect 27454 7046 27484 7098
rect 27508 7046 27518 7098
rect 27518 7046 27564 7098
rect 27268 7044 27324 7046
rect 27348 7044 27404 7046
rect 27428 7044 27484 7046
rect 27508 7044 27564 7046
rect 27268 6010 27324 6012
rect 27348 6010 27404 6012
rect 27428 6010 27484 6012
rect 27508 6010 27564 6012
rect 27268 5958 27314 6010
rect 27314 5958 27324 6010
rect 27348 5958 27378 6010
rect 27378 5958 27390 6010
rect 27390 5958 27404 6010
rect 27428 5958 27442 6010
rect 27442 5958 27454 6010
rect 27454 5958 27484 6010
rect 27508 5958 27518 6010
rect 27518 5958 27564 6010
rect 27268 5956 27324 5958
rect 27348 5956 27404 5958
rect 27428 5956 27484 5958
rect 27508 5956 27564 5958
rect 27268 4922 27324 4924
rect 27348 4922 27404 4924
rect 27428 4922 27484 4924
rect 27508 4922 27564 4924
rect 27268 4870 27314 4922
rect 27314 4870 27324 4922
rect 27348 4870 27378 4922
rect 27378 4870 27390 4922
rect 27390 4870 27404 4922
rect 27428 4870 27442 4922
rect 27442 4870 27454 4922
rect 27454 4870 27484 4922
rect 27508 4870 27518 4922
rect 27518 4870 27564 4922
rect 27268 4868 27324 4870
rect 27348 4868 27404 4870
rect 27428 4868 27484 4870
rect 27508 4868 27564 4870
rect 27268 3834 27324 3836
rect 27348 3834 27404 3836
rect 27428 3834 27484 3836
rect 27508 3834 27564 3836
rect 27268 3782 27314 3834
rect 27314 3782 27324 3834
rect 27348 3782 27378 3834
rect 27378 3782 27390 3834
rect 27390 3782 27404 3834
rect 27428 3782 27442 3834
rect 27442 3782 27454 3834
rect 27454 3782 27484 3834
rect 27508 3782 27518 3834
rect 27518 3782 27564 3834
rect 27268 3780 27324 3782
rect 27348 3780 27404 3782
rect 27428 3780 27484 3782
rect 27508 3780 27564 3782
rect 27268 2746 27324 2748
rect 27348 2746 27404 2748
rect 27428 2746 27484 2748
rect 27508 2746 27564 2748
rect 27268 2694 27314 2746
rect 27314 2694 27324 2746
rect 27348 2694 27378 2746
rect 27378 2694 27390 2746
rect 27390 2694 27404 2746
rect 27428 2694 27442 2746
rect 27442 2694 27454 2746
rect 27454 2694 27484 2746
rect 27508 2694 27518 2746
rect 27518 2694 27564 2746
rect 27268 2692 27324 2694
rect 27348 2692 27404 2694
rect 27428 2692 27484 2694
rect 27508 2692 27564 2694
rect 27268 1658 27324 1660
rect 27348 1658 27404 1660
rect 27428 1658 27484 1660
rect 27508 1658 27564 1660
rect 27268 1606 27314 1658
rect 27314 1606 27324 1658
rect 27348 1606 27378 1658
rect 27378 1606 27390 1658
rect 27390 1606 27404 1658
rect 27428 1606 27442 1658
rect 27442 1606 27454 1658
rect 27454 1606 27484 1658
rect 27508 1606 27518 1658
rect 27518 1606 27564 1658
rect 27268 1604 27324 1606
rect 27348 1604 27404 1606
rect 27428 1604 27484 1606
rect 27508 1604 27564 1606
rect 27268 570 27324 572
rect 27348 570 27404 572
rect 27428 570 27484 572
rect 27508 570 27564 572
rect 27268 518 27314 570
rect 27314 518 27324 570
rect 27348 518 27378 570
rect 27378 518 27390 570
rect 27390 518 27404 570
rect 27428 518 27442 570
rect 27442 518 27454 570
rect 27454 518 27484 570
rect 27508 518 27518 570
rect 27518 518 27564 570
rect 27268 516 27324 518
rect 27348 516 27404 518
rect 27428 516 27484 518
rect 27508 516 27564 518
<< metal3 >>
rect 3752 17440 4068 17441
rect 3752 17376 3758 17440
rect 3822 17376 3838 17440
rect 3902 17376 3918 17440
rect 3982 17376 3998 17440
rect 4062 17376 4068 17440
rect 3752 17375 4068 17376
rect 10468 17440 10784 17441
rect 10468 17376 10474 17440
rect 10538 17376 10554 17440
rect 10618 17376 10634 17440
rect 10698 17376 10714 17440
rect 10778 17376 10784 17440
rect 10468 17375 10784 17376
rect 17184 17440 17500 17441
rect 17184 17376 17190 17440
rect 17254 17376 17270 17440
rect 17334 17376 17350 17440
rect 17414 17376 17430 17440
rect 17494 17376 17500 17440
rect 17184 17375 17500 17376
rect 23900 17440 24216 17441
rect 23900 17376 23906 17440
rect 23970 17376 23986 17440
rect 24050 17376 24066 17440
rect 24130 17376 24146 17440
rect 24210 17376 24216 17440
rect 23900 17375 24216 17376
rect 7110 16896 7426 16897
rect 7110 16832 7116 16896
rect 7180 16832 7196 16896
rect 7260 16832 7276 16896
rect 7340 16832 7356 16896
rect 7420 16832 7426 16896
rect 7110 16831 7426 16832
rect 13826 16896 14142 16897
rect 13826 16832 13832 16896
rect 13896 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14142 16896
rect 13826 16831 14142 16832
rect 20542 16896 20858 16897
rect 20542 16832 20548 16896
rect 20612 16832 20628 16896
rect 20692 16832 20708 16896
rect 20772 16832 20788 16896
rect 20852 16832 20858 16896
rect 20542 16831 20858 16832
rect 27258 16896 27574 16897
rect 27258 16832 27264 16896
rect 27328 16832 27344 16896
rect 27408 16832 27424 16896
rect 27488 16832 27504 16896
rect 27568 16832 27574 16896
rect 27258 16831 27574 16832
rect 11237 16554 11303 16557
rect 15101 16554 15167 16557
rect 17033 16554 17099 16557
rect 11237 16552 17099 16554
rect 11237 16496 11242 16552
rect 11298 16496 15106 16552
rect 15162 16496 17038 16552
rect 17094 16496 17099 16552
rect 11237 16494 17099 16496
rect 11237 16491 11303 16494
rect 15101 16491 15167 16494
rect 17033 16491 17099 16494
rect 3752 16352 4068 16353
rect 3752 16288 3758 16352
rect 3822 16288 3838 16352
rect 3902 16288 3918 16352
rect 3982 16288 3998 16352
rect 4062 16288 4068 16352
rect 3752 16287 4068 16288
rect 10468 16352 10784 16353
rect 10468 16288 10474 16352
rect 10538 16288 10554 16352
rect 10618 16288 10634 16352
rect 10698 16288 10714 16352
rect 10778 16288 10784 16352
rect 10468 16287 10784 16288
rect 17184 16352 17500 16353
rect 17184 16288 17190 16352
rect 17254 16288 17270 16352
rect 17334 16288 17350 16352
rect 17414 16288 17430 16352
rect 17494 16288 17500 16352
rect 17184 16287 17500 16288
rect 23900 16352 24216 16353
rect 23900 16288 23906 16352
rect 23970 16288 23986 16352
rect 24050 16288 24066 16352
rect 24130 16288 24146 16352
rect 24210 16288 24216 16352
rect 23900 16287 24216 16288
rect 7110 15808 7426 15809
rect 7110 15744 7116 15808
rect 7180 15744 7196 15808
rect 7260 15744 7276 15808
rect 7340 15744 7356 15808
rect 7420 15744 7426 15808
rect 7110 15743 7426 15744
rect 13826 15808 14142 15809
rect 13826 15744 13832 15808
rect 13896 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14142 15808
rect 13826 15743 14142 15744
rect 20542 15808 20858 15809
rect 20542 15744 20548 15808
rect 20612 15744 20628 15808
rect 20692 15744 20708 15808
rect 20772 15744 20788 15808
rect 20852 15744 20858 15808
rect 20542 15743 20858 15744
rect 27258 15808 27574 15809
rect 27258 15744 27264 15808
rect 27328 15744 27344 15808
rect 27408 15744 27424 15808
rect 27488 15744 27504 15808
rect 27568 15744 27574 15808
rect 27258 15743 27574 15744
rect 16757 15466 16823 15469
rect 17718 15466 17724 15468
rect 16757 15464 17724 15466
rect 16757 15408 16762 15464
rect 16818 15408 17724 15464
rect 16757 15406 17724 15408
rect 16757 15403 16823 15406
rect 17718 15404 17724 15406
rect 17788 15404 17794 15468
rect 3752 15264 4068 15265
rect 3752 15200 3758 15264
rect 3822 15200 3838 15264
rect 3902 15200 3918 15264
rect 3982 15200 3998 15264
rect 4062 15200 4068 15264
rect 3752 15199 4068 15200
rect 10468 15264 10784 15265
rect 10468 15200 10474 15264
rect 10538 15200 10554 15264
rect 10618 15200 10634 15264
rect 10698 15200 10714 15264
rect 10778 15200 10784 15264
rect 10468 15199 10784 15200
rect 17184 15264 17500 15265
rect 17184 15200 17190 15264
rect 17254 15200 17270 15264
rect 17334 15200 17350 15264
rect 17414 15200 17430 15264
rect 17494 15200 17500 15264
rect 17184 15199 17500 15200
rect 23900 15264 24216 15265
rect 23900 15200 23906 15264
rect 23970 15200 23986 15264
rect 24050 15200 24066 15264
rect 24130 15200 24146 15264
rect 24210 15200 24216 15264
rect 23900 15199 24216 15200
rect 11881 15194 11947 15197
rect 16389 15194 16455 15197
rect 11881 15192 16455 15194
rect 11881 15136 11886 15192
rect 11942 15136 16394 15192
rect 16450 15136 16455 15192
rect 11881 15134 16455 15136
rect 11881 15131 11947 15134
rect 16389 15131 16455 15134
rect 8477 15058 8543 15061
rect 23473 15058 23539 15061
rect 8477 15056 23539 15058
rect 8477 15000 8482 15056
rect 8538 15000 23478 15056
rect 23534 15000 23539 15056
rect 8477 14998 23539 15000
rect 8477 14995 8543 14998
rect 23473 14995 23539 14998
rect 4889 14922 4955 14925
rect 8477 14922 8543 14925
rect 13905 14922 13971 14925
rect 4889 14920 13971 14922
rect 4889 14864 4894 14920
rect 4950 14864 8482 14920
rect 8538 14864 13910 14920
rect 13966 14864 13971 14920
rect 4889 14862 13971 14864
rect 4889 14859 4955 14862
rect 8477 14859 8543 14862
rect 13905 14859 13971 14862
rect 7110 14720 7426 14721
rect 7110 14656 7116 14720
rect 7180 14656 7196 14720
rect 7260 14656 7276 14720
rect 7340 14656 7356 14720
rect 7420 14656 7426 14720
rect 7110 14655 7426 14656
rect 13826 14720 14142 14721
rect 13826 14656 13832 14720
rect 13896 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14142 14720
rect 13826 14655 14142 14656
rect 20542 14720 20858 14721
rect 20542 14656 20548 14720
rect 20612 14656 20628 14720
rect 20692 14656 20708 14720
rect 20772 14656 20788 14720
rect 20852 14656 20858 14720
rect 20542 14655 20858 14656
rect 27258 14720 27574 14721
rect 27258 14656 27264 14720
rect 27328 14656 27344 14720
rect 27408 14656 27424 14720
rect 27488 14656 27504 14720
rect 27568 14656 27574 14720
rect 27258 14655 27574 14656
rect 19425 14378 19491 14381
rect 23473 14378 23539 14381
rect 19425 14376 23539 14378
rect 19425 14320 19430 14376
rect 19486 14320 23478 14376
rect 23534 14320 23539 14376
rect 19425 14318 23539 14320
rect 19425 14315 19491 14318
rect 23473 14315 23539 14318
rect 3752 14176 4068 14177
rect 3752 14112 3758 14176
rect 3822 14112 3838 14176
rect 3902 14112 3918 14176
rect 3982 14112 3998 14176
rect 4062 14112 4068 14176
rect 3752 14111 4068 14112
rect 10468 14176 10784 14177
rect 10468 14112 10474 14176
rect 10538 14112 10554 14176
rect 10618 14112 10634 14176
rect 10698 14112 10714 14176
rect 10778 14112 10784 14176
rect 10468 14111 10784 14112
rect 17184 14176 17500 14177
rect 17184 14112 17190 14176
rect 17254 14112 17270 14176
rect 17334 14112 17350 14176
rect 17414 14112 17430 14176
rect 17494 14112 17500 14176
rect 17184 14111 17500 14112
rect 23900 14176 24216 14177
rect 23900 14112 23906 14176
rect 23970 14112 23986 14176
rect 24050 14112 24066 14176
rect 24130 14112 24146 14176
rect 24210 14112 24216 14176
rect 23900 14111 24216 14112
rect 5809 13970 5875 13973
rect 9581 13970 9647 13973
rect 5809 13968 9647 13970
rect 5809 13912 5814 13968
rect 5870 13912 9586 13968
rect 9642 13912 9647 13968
rect 5809 13910 9647 13912
rect 5809 13907 5875 13910
rect 9581 13907 9647 13910
rect 8017 13834 8083 13837
rect 9121 13834 9187 13837
rect 22369 13836 22435 13837
rect 22318 13834 22324 13836
rect 8017 13832 9187 13834
rect 8017 13776 8022 13832
rect 8078 13776 9126 13832
rect 9182 13776 9187 13832
rect 8017 13774 9187 13776
rect 22278 13774 22324 13834
rect 22388 13832 22435 13836
rect 22430 13776 22435 13832
rect 8017 13771 8083 13774
rect 9121 13771 9187 13774
rect 22318 13772 22324 13774
rect 22388 13772 22435 13776
rect 22369 13771 22435 13772
rect 26233 13834 26299 13837
rect 27153 13834 27219 13837
rect 26233 13832 27219 13834
rect 26233 13776 26238 13832
rect 26294 13776 27158 13832
rect 27214 13776 27219 13832
rect 26233 13774 27219 13776
rect 26233 13771 26299 13774
rect 27153 13771 27219 13774
rect 7110 13632 7426 13633
rect 7110 13568 7116 13632
rect 7180 13568 7196 13632
rect 7260 13568 7276 13632
rect 7340 13568 7356 13632
rect 7420 13568 7426 13632
rect 7110 13567 7426 13568
rect 13826 13632 14142 13633
rect 13826 13568 13832 13632
rect 13896 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14142 13632
rect 13826 13567 14142 13568
rect 20542 13632 20858 13633
rect 20542 13568 20548 13632
rect 20612 13568 20628 13632
rect 20692 13568 20708 13632
rect 20772 13568 20788 13632
rect 20852 13568 20858 13632
rect 20542 13567 20858 13568
rect 27258 13632 27574 13633
rect 27258 13568 27264 13632
rect 27328 13568 27344 13632
rect 27408 13568 27424 13632
rect 27488 13568 27504 13632
rect 27568 13568 27574 13632
rect 27258 13567 27574 13568
rect 12617 13426 12683 13429
rect 18137 13426 18203 13429
rect 12617 13424 18203 13426
rect 12617 13368 12622 13424
rect 12678 13368 18142 13424
rect 18198 13368 18203 13424
rect 12617 13366 18203 13368
rect 12617 13363 12683 13366
rect 18137 13363 18203 13366
rect 3752 13088 4068 13089
rect 3752 13024 3758 13088
rect 3822 13024 3838 13088
rect 3902 13024 3918 13088
rect 3982 13024 3998 13088
rect 4062 13024 4068 13088
rect 3752 13023 4068 13024
rect 10468 13088 10784 13089
rect 10468 13024 10474 13088
rect 10538 13024 10554 13088
rect 10618 13024 10634 13088
rect 10698 13024 10714 13088
rect 10778 13024 10784 13088
rect 10468 13023 10784 13024
rect 17184 13088 17500 13089
rect 17184 13024 17190 13088
rect 17254 13024 17270 13088
rect 17334 13024 17350 13088
rect 17414 13024 17430 13088
rect 17494 13024 17500 13088
rect 17184 13023 17500 13024
rect 23900 13088 24216 13089
rect 23900 13024 23906 13088
rect 23970 13024 23986 13088
rect 24050 13024 24066 13088
rect 24130 13024 24146 13088
rect 24210 13024 24216 13088
rect 23900 13023 24216 13024
rect 10501 12882 10567 12885
rect 12525 12882 12591 12885
rect 10501 12880 12591 12882
rect 10501 12824 10506 12880
rect 10562 12824 12530 12880
rect 12586 12824 12591 12880
rect 10501 12822 12591 12824
rect 10501 12819 10567 12822
rect 12525 12819 12591 12822
rect 12249 12746 12315 12749
rect 18137 12746 18203 12749
rect 12249 12744 18203 12746
rect 12249 12688 12254 12744
rect 12310 12688 18142 12744
rect 18198 12688 18203 12744
rect 12249 12686 18203 12688
rect 12249 12683 12315 12686
rect 18137 12683 18203 12686
rect 25313 12746 25379 12749
rect 25313 12744 25514 12746
rect 25313 12688 25318 12744
rect 25374 12688 25514 12744
rect 25313 12686 25514 12688
rect 25313 12683 25379 12686
rect 17718 12548 17724 12612
rect 17788 12610 17794 12612
rect 18045 12610 18111 12613
rect 17788 12608 18111 12610
rect 17788 12552 18050 12608
rect 18106 12552 18111 12608
rect 17788 12550 18111 12552
rect 17788 12548 17794 12550
rect 18045 12547 18111 12550
rect 7110 12544 7426 12545
rect 7110 12480 7116 12544
rect 7180 12480 7196 12544
rect 7260 12480 7276 12544
rect 7340 12480 7356 12544
rect 7420 12480 7426 12544
rect 7110 12479 7426 12480
rect 13826 12544 14142 12545
rect 13826 12480 13832 12544
rect 13896 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14142 12544
rect 13826 12479 14142 12480
rect 20542 12544 20858 12545
rect 20542 12480 20548 12544
rect 20612 12480 20628 12544
rect 20692 12480 20708 12544
rect 20772 12480 20788 12544
rect 20852 12480 20858 12544
rect 20542 12479 20858 12480
rect 25454 12477 25514 12686
rect 27258 12544 27574 12545
rect 27258 12480 27264 12544
rect 27328 12480 27344 12544
rect 27408 12480 27424 12544
rect 27488 12480 27504 12544
rect 27568 12480 27574 12544
rect 27258 12479 27574 12480
rect 8201 12474 8267 12477
rect 10869 12474 10935 12477
rect 8201 12472 10935 12474
rect 8201 12416 8206 12472
rect 8262 12416 10874 12472
rect 10930 12416 10935 12472
rect 8201 12414 10935 12416
rect 8201 12411 8267 12414
rect 10869 12411 10935 12414
rect 25405 12472 25514 12477
rect 25405 12416 25410 12472
rect 25466 12416 25514 12472
rect 25405 12414 25514 12416
rect 25405 12411 25471 12414
rect 7833 12338 7899 12341
rect 21081 12338 21147 12341
rect 7833 12336 21147 12338
rect 7833 12280 7838 12336
rect 7894 12280 21086 12336
rect 21142 12280 21147 12336
rect 7833 12278 21147 12280
rect 7833 12275 7899 12278
rect 21081 12275 21147 12278
rect 26141 12340 26207 12341
rect 26141 12336 26188 12340
rect 26252 12338 26258 12340
rect 26141 12280 26146 12336
rect 26141 12276 26188 12280
rect 26252 12278 26298 12338
rect 26252 12276 26258 12278
rect 26141 12275 26207 12276
rect 10174 12140 10180 12204
rect 10244 12202 10250 12204
rect 10869 12202 10935 12205
rect 24577 12202 24643 12205
rect 10244 12200 10935 12202
rect 10244 12144 10874 12200
rect 10930 12144 10935 12200
rect 10244 12142 10935 12144
rect 10244 12140 10250 12142
rect 10869 12139 10935 12142
rect 22050 12200 24643 12202
rect 22050 12144 24582 12200
rect 24638 12144 24643 12200
rect 22050 12142 24643 12144
rect 3752 12000 4068 12001
rect 3752 11936 3758 12000
rect 3822 11936 3838 12000
rect 3902 11936 3918 12000
rect 3982 11936 3998 12000
rect 4062 11936 4068 12000
rect 3752 11935 4068 11936
rect 10468 12000 10784 12001
rect 10468 11936 10474 12000
rect 10538 11936 10554 12000
rect 10618 11936 10634 12000
rect 10698 11936 10714 12000
rect 10778 11936 10784 12000
rect 10468 11935 10784 11936
rect 17184 12000 17500 12001
rect 17184 11936 17190 12000
rect 17254 11936 17270 12000
rect 17334 11936 17350 12000
rect 17414 11936 17430 12000
rect 17494 11936 17500 12000
rect 17184 11935 17500 11936
rect 17585 11930 17651 11933
rect 22050 11930 22110 12142
rect 24577 12139 24643 12142
rect 23900 12000 24216 12001
rect 23900 11936 23906 12000
rect 23970 11936 23986 12000
rect 24050 11936 24066 12000
rect 24130 11936 24146 12000
rect 24210 11936 24216 12000
rect 23900 11935 24216 11936
rect 17585 11928 22110 11930
rect 17585 11872 17590 11928
rect 17646 11872 22110 11928
rect 17585 11870 22110 11872
rect 17585 11867 17651 11870
rect 11697 11794 11763 11797
rect 17585 11794 17651 11797
rect 11697 11792 17651 11794
rect 11697 11736 11702 11792
rect 11758 11736 17590 11792
rect 17646 11736 17651 11792
rect 11697 11734 17651 11736
rect 11697 11731 11763 11734
rect 17585 11731 17651 11734
rect 20118 11734 21834 11794
rect 7465 11658 7531 11661
rect 18505 11658 18571 11661
rect 20118 11658 20178 11734
rect 21541 11658 21607 11661
rect 7465 11656 20178 11658
rect 7465 11600 7470 11656
rect 7526 11600 18510 11656
rect 18566 11600 20178 11656
rect 7465 11598 20178 11600
rect 20302 11656 21607 11658
rect 20302 11600 21546 11656
rect 21602 11600 21607 11656
rect 20302 11598 21607 11600
rect 21774 11658 21834 11734
rect 22553 11658 22619 11661
rect 21774 11656 22619 11658
rect 21774 11600 22558 11656
rect 22614 11600 22619 11656
rect 21774 11598 22619 11600
rect 7465 11595 7531 11598
rect 18505 11595 18571 11598
rect 11053 11522 11119 11525
rect 11605 11522 11671 11525
rect 18689 11524 18755 11525
rect 11053 11520 11671 11522
rect 11053 11464 11058 11520
rect 11114 11464 11610 11520
rect 11666 11464 11671 11520
rect 11053 11462 11671 11464
rect 11053 11459 11119 11462
rect 11605 11459 11671 11462
rect 18638 11460 18644 11524
rect 18708 11522 18755 11524
rect 20302 11522 20362 11598
rect 21541 11595 21607 11598
rect 22553 11595 22619 11598
rect 18708 11520 20362 11522
rect 18750 11464 20362 11520
rect 18708 11462 20362 11464
rect 18708 11460 18755 11462
rect 18689 11459 18755 11460
rect 7110 11456 7426 11457
rect 7110 11392 7116 11456
rect 7180 11392 7196 11456
rect 7260 11392 7276 11456
rect 7340 11392 7356 11456
rect 7420 11392 7426 11456
rect 7110 11391 7426 11392
rect 13826 11456 14142 11457
rect 13826 11392 13832 11456
rect 13896 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14142 11456
rect 13826 11391 14142 11392
rect 20542 11456 20858 11457
rect 20542 11392 20548 11456
rect 20612 11392 20628 11456
rect 20692 11392 20708 11456
rect 20772 11392 20788 11456
rect 20852 11392 20858 11456
rect 20542 11391 20858 11392
rect 27258 11456 27574 11457
rect 27258 11392 27264 11456
rect 27328 11392 27344 11456
rect 27408 11392 27424 11456
rect 27488 11392 27504 11456
rect 27568 11392 27574 11456
rect 27258 11391 27574 11392
rect 9673 11386 9739 11389
rect 13629 11386 13695 11389
rect 9673 11384 13695 11386
rect 9673 11328 9678 11384
rect 9734 11328 13634 11384
rect 13690 11328 13695 11384
rect 9673 11326 13695 11328
rect 9673 11323 9739 11326
rect 13629 11323 13695 11326
rect 11605 11250 11671 11253
rect 21357 11250 21423 11253
rect 11605 11248 21423 11250
rect 11605 11192 11610 11248
rect 11666 11192 21362 11248
rect 21418 11192 21423 11248
rect 11605 11190 21423 11192
rect 11605 11187 11671 11190
rect 21357 11187 21423 11190
rect 18270 11052 18276 11116
rect 18340 11114 18346 11116
rect 18413 11114 18479 11117
rect 18340 11112 18479 11114
rect 18340 11056 18418 11112
rect 18474 11056 18479 11112
rect 18340 11054 18479 11056
rect 18340 11052 18346 11054
rect 18413 11051 18479 11054
rect 22553 11114 22619 11117
rect 24117 11114 24183 11117
rect 22553 11112 24183 11114
rect 22553 11056 22558 11112
rect 22614 11056 24122 11112
rect 24178 11056 24183 11112
rect 22553 11054 24183 11056
rect 22553 11051 22619 11054
rect 24117 11051 24183 11054
rect 3752 10912 4068 10913
rect 3752 10848 3758 10912
rect 3822 10848 3838 10912
rect 3902 10848 3918 10912
rect 3982 10848 3998 10912
rect 4062 10848 4068 10912
rect 3752 10847 4068 10848
rect 10468 10912 10784 10913
rect 10468 10848 10474 10912
rect 10538 10848 10554 10912
rect 10618 10848 10634 10912
rect 10698 10848 10714 10912
rect 10778 10848 10784 10912
rect 10468 10847 10784 10848
rect 17184 10912 17500 10913
rect 17184 10848 17190 10912
rect 17254 10848 17270 10912
rect 17334 10848 17350 10912
rect 17414 10848 17430 10912
rect 17494 10848 17500 10912
rect 17184 10847 17500 10848
rect 23900 10912 24216 10913
rect 23900 10848 23906 10912
rect 23970 10848 23986 10912
rect 24050 10848 24066 10912
rect 24130 10848 24146 10912
rect 24210 10848 24216 10912
rect 23900 10847 24216 10848
rect 18597 10842 18663 10845
rect 23749 10842 23815 10845
rect 18597 10840 23815 10842
rect 18597 10784 18602 10840
rect 18658 10784 23754 10840
rect 23810 10784 23815 10840
rect 18597 10782 23815 10784
rect 18597 10779 18663 10782
rect 23749 10779 23815 10782
rect 20529 10706 20595 10709
rect 24117 10706 24183 10709
rect 20529 10704 24183 10706
rect 20529 10648 20534 10704
rect 20590 10648 24122 10704
rect 24178 10648 24183 10704
rect 20529 10646 24183 10648
rect 20529 10643 20595 10646
rect 24117 10643 24183 10646
rect 11973 10570 12039 10573
rect 12709 10570 12775 10573
rect 11973 10568 12775 10570
rect 11973 10512 11978 10568
rect 12034 10512 12714 10568
rect 12770 10512 12775 10568
rect 11973 10510 12775 10512
rect 11973 10507 12039 10510
rect 12709 10507 12775 10510
rect 7110 10368 7426 10369
rect 7110 10304 7116 10368
rect 7180 10304 7196 10368
rect 7260 10304 7276 10368
rect 7340 10304 7356 10368
rect 7420 10304 7426 10368
rect 7110 10303 7426 10304
rect 13826 10368 14142 10369
rect 13826 10304 13832 10368
rect 13896 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14142 10368
rect 13826 10303 14142 10304
rect 20542 10368 20858 10369
rect 20542 10304 20548 10368
rect 20612 10304 20628 10368
rect 20692 10304 20708 10368
rect 20772 10304 20788 10368
rect 20852 10304 20858 10368
rect 20542 10303 20858 10304
rect 27258 10368 27574 10369
rect 27258 10304 27264 10368
rect 27328 10304 27344 10368
rect 27408 10304 27424 10368
rect 27488 10304 27504 10368
rect 27568 10304 27574 10368
rect 27258 10303 27574 10304
rect 3752 9824 4068 9825
rect 3752 9760 3758 9824
rect 3822 9760 3838 9824
rect 3902 9760 3918 9824
rect 3982 9760 3998 9824
rect 4062 9760 4068 9824
rect 3752 9759 4068 9760
rect 10468 9824 10784 9825
rect 10468 9760 10474 9824
rect 10538 9760 10554 9824
rect 10618 9760 10634 9824
rect 10698 9760 10714 9824
rect 10778 9760 10784 9824
rect 10468 9759 10784 9760
rect 17184 9824 17500 9825
rect 17184 9760 17190 9824
rect 17254 9760 17270 9824
rect 17334 9760 17350 9824
rect 17414 9760 17430 9824
rect 17494 9760 17500 9824
rect 17184 9759 17500 9760
rect 23900 9824 24216 9825
rect 23900 9760 23906 9824
rect 23970 9760 23986 9824
rect 24050 9760 24066 9824
rect 24130 9760 24146 9824
rect 24210 9760 24216 9824
rect 23900 9759 24216 9760
rect 12065 9754 12131 9757
rect 15193 9754 15259 9757
rect 12065 9752 15259 9754
rect 12065 9696 12070 9752
rect 12126 9696 15198 9752
rect 15254 9696 15259 9752
rect 12065 9694 15259 9696
rect 12065 9691 12131 9694
rect 15193 9691 15259 9694
rect 10174 9556 10180 9620
rect 10244 9618 10250 9620
rect 13997 9618 14063 9621
rect 18638 9618 18644 9620
rect 10244 9616 18644 9618
rect 10244 9560 14002 9616
rect 14058 9560 18644 9616
rect 10244 9558 18644 9560
rect 10244 9556 10250 9558
rect 13997 9555 14063 9558
rect 18638 9556 18644 9558
rect 18708 9618 18714 9620
rect 20294 9618 20300 9620
rect 18708 9558 20300 9618
rect 18708 9556 18714 9558
rect 20294 9556 20300 9558
rect 20364 9556 20370 9620
rect 20897 9618 20963 9621
rect 24853 9618 24919 9621
rect 25313 9618 25379 9621
rect 20897 9616 25379 9618
rect 20897 9560 20902 9616
rect 20958 9560 24858 9616
rect 24914 9560 25318 9616
rect 25374 9560 25379 9616
rect 20897 9558 25379 9560
rect 20897 9555 20963 9558
rect 24853 9555 24919 9558
rect 25313 9555 25379 9558
rect 7833 9482 7899 9485
rect 11605 9482 11671 9485
rect 7833 9480 11671 9482
rect 7833 9424 7838 9480
rect 7894 9424 11610 9480
rect 11666 9424 11671 9480
rect 7833 9422 11671 9424
rect 7833 9419 7899 9422
rect 11605 9419 11671 9422
rect 15745 9482 15811 9485
rect 26182 9482 26188 9484
rect 15745 9480 26188 9482
rect 15745 9424 15750 9480
rect 15806 9424 26188 9480
rect 15745 9422 26188 9424
rect 15745 9419 15811 9422
rect 26182 9420 26188 9422
rect 26252 9420 26258 9484
rect 16573 9346 16639 9349
rect 17125 9346 17191 9349
rect 17769 9346 17835 9349
rect 16573 9344 17835 9346
rect 16573 9288 16578 9344
rect 16634 9288 17130 9344
rect 17186 9288 17774 9344
rect 17830 9288 17835 9344
rect 16573 9286 17835 9288
rect 16573 9283 16639 9286
rect 17125 9283 17191 9286
rect 17769 9283 17835 9286
rect 7110 9280 7426 9281
rect 7110 9216 7116 9280
rect 7180 9216 7196 9280
rect 7260 9216 7276 9280
rect 7340 9216 7356 9280
rect 7420 9216 7426 9280
rect 7110 9215 7426 9216
rect 13826 9280 14142 9281
rect 13826 9216 13832 9280
rect 13896 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14142 9280
rect 13826 9215 14142 9216
rect 20542 9280 20858 9281
rect 20542 9216 20548 9280
rect 20612 9216 20628 9280
rect 20692 9216 20708 9280
rect 20772 9216 20788 9280
rect 20852 9216 20858 9280
rect 20542 9215 20858 9216
rect 27258 9280 27574 9281
rect 27258 9216 27264 9280
rect 27328 9216 27344 9280
rect 27408 9216 27424 9280
rect 27488 9216 27504 9280
rect 27568 9216 27574 9280
rect 27258 9215 27574 9216
rect 12249 9074 12315 9077
rect 13721 9074 13787 9077
rect 16849 9074 16915 9077
rect 12249 9072 16915 9074
rect 12249 9016 12254 9072
rect 12310 9016 13726 9072
rect 13782 9016 16854 9072
rect 16910 9016 16915 9072
rect 12249 9014 16915 9016
rect 12249 9011 12315 9014
rect 13721 9011 13787 9014
rect 16849 9011 16915 9014
rect 10501 8938 10567 8941
rect 21173 8938 21239 8941
rect 10501 8936 21239 8938
rect 10501 8880 10506 8936
rect 10562 8880 21178 8936
rect 21234 8880 21239 8936
rect 10501 8878 21239 8880
rect 10501 8875 10567 8878
rect 21173 8875 21239 8878
rect 3752 8736 4068 8737
rect 3752 8672 3758 8736
rect 3822 8672 3838 8736
rect 3902 8672 3918 8736
rect 3982 8672 3998 8736
rect 4062 8672 4068 8736
rect 3752 8671 4068 8672
rect 10468 8736 10784 8737
rect 10468 8672 10474 8736
rect 10538 8672 10554 8736
rect 10618 8672 10634 8736
rect 10698 8672 10714 8736
rect 10778 8672 10784 8736
rect 10468 8671 10784 8672
rect 17184 8736 17500 8737
rect 17184 8672 17190 8736
rect 17254 8672 17270 8736
rect 17334 8672 17350 8736
rect 17414 8672 17430 8736
rect 17494 8672 17500 8736
rect 17184 8671 17500 8672
rect 23900 8736 24216 8737
rect 23900 8672 23906 8736
rect 23970 8672 23986 8736
rect 24050 8672 24066 8736
rect 24130 8672 24146 8736
rect 24210 8672 24216 8736
rect 23900 8671 24216 8672
rect 12341 8666 12407 8669
rect 12801 8666 12867 8669
rect 13813 8666 13879 8669
rect 12341 8664 13879 8666
rect 12341 8608 12346 8664
rect 12402 8608 12806 8664
rect 12862 8608 13818 8664
rect 13874 8608 13879 8664
rect 12341 8606 13879 8608
rect 12341 8603 12407 8606
rect 12801 8603 12867 8606
rect 13813 8603 13879 8606
rect 10041 8530 10107 8533
rect 13905 8530 13971 8533
rect 17677 8530 17743 8533
rect 10041 8528 17743 8530
rect 10041 8472 10046 8528
rect 10102 8472 13910 8528
rect 13966 8472 17682 8528
rect 17738 8472 17743 8528
rect 10041 8470 17743 8472
rect 10041 8467 10107 8470
rect 13905 8467 13971 8470
rect 17677 8467 17743 8470
rect 5809 8394 5875 8397
rect 17718 8394 17724 8396
rect 5809 8392 17724 8394
rect 5809 8336 5814 8392
rect 5870 8336 17724 8392
rect 5809 8334 17724 8336
rect 5809 8331 5875 8334
rect 17718 8332 17724 8334
rect 17788 8332 17794 8396
rect 7110 8192 7426 8193
rect 7110 8128 7116 8192
rect 7180 8128 7196 8192
rect 7260 8128 7276 8192
rect 7340 8128 7356 8192
rect 7420 8128 7426 8192
rect 7110 8127 7426 8128
rect 13826 8192 14142 8193
rect 13826 8128 13832 8192
rect 13896 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14142 8192
rect 13826 8127 14142 8128
rect 20542 8192 20858 8193
rect 20542 8128 20548 8192
rect 20612 8128 20628 8192
rect 20692 8128 20708 8192
rect 20772 8128 20788 8192
rect 20852 8128 20858 8192
rect 20542 8127 20858 8128
rect 27258 8192 27574 8193
rect 27258 8128 27264 8192
rect 27328 8128 27344 8192
rect 27408 8128 27424 8192
rect 27488 8128 27504 8192
rect 27568 8128 27574 8192
rect 27258 8127 27574 8128
rect 11513 8122 11579 8125
rect 13445 8122 13511 8125
rect 13629 8122 13695 8125
rect 11513 8120 13695 8122
rect 11513 8064 11518 8120
rect 11574 8064 13450 8120
rect 13506 8064 13634 8120
rect 13690 8064 13695 8120
rect 11513 8062 13695 8064
rect 11513 8059 11579 8062
rect 13445 8059 13511 8062
rect 13629 8059 13695 8062
rect 8845 7986 8911 7989
rect 16665 7986 16731 7989
rect 8845 7984 16731 7986
rect 8845 7928 8850 7984
rect 8906 7928 16670 7984
rect 16726 7928 16731 7984
rect 8845 7926 16731 7928
rect 8845 7923 8911 7926
rect 16665 7923 16731 7926
rect 3752 7648 4068 7649
rect 3752 7584 3758 7648
rect 3822 7584 3838 7648
rect 3902 7584 3918 7648
rect 3982 7584 3998 7648
rect 4062 7584 4068 7648
rect 3752 7583 4068 7584
rect 10468 7648 10784 7649
rect 10468 7584 10474 7648
rect 10538 7584 10554 7648
rect 10618 7584 10634 7648
rect 10698 7584 10714 7648
rect 10778 7584 10784 7648
rect 10468 7583 10784 7584
rect 17184 7648 17500 7649
rect 17184 7584 17190 7648
rect 17254 7584 17270 7648
rect 17334 7584 17350 7648
rect 17414 7584 17430 7648
rect 17494 7584 17500 7648
rect 17184 7583 17500 7584
rect 23900 7648 24216 7649
rect 23900 7584 23906 7648
rect 23970 7584 23986 7648
rect 24050 7584 24066 7648
rect 24130 7584 24146 7648
rect 24210 7584 24216 7648
rect 23900 7583 24216 7584
rect 7110 7104 7426 7105
rect 7110 7040 7116 7104
rect 7180 7040 7196 7104
rect 7260 7040 7276 7104
rect 7340 7040 7356 7104
rect 7420 7040 7426 7104
rect 7110 7039 7426 7040
rect 13826 7104 14142 7105
rect 13826 7040 13832 7104
rect 13896 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14142 7104
rect 13826 7039 14142 7040
rect 20542 7104 20858 7105
rect 20542 7040 20548 7104
rect 20612 7040 20628 7104
rect 20692 7040 20708 7104
rect 20772 7040 20788 7104
rect 20852 7040 20858 7104
rect 20542 7039 20858 7040
rect 27258 7104 27574 7105
rect 27258 7040 27264 7104
rect 27328 7040 27344 7104
rect 27408 7040 27424 7104
rect 27488 7040 27504 7104
rect 27568 7040 27574 7104
rect 27258 7039 27574 7040
rect 3752 6560 4068 6561
rect 3752 6496 3758 6560
rect 3822 6496 3838 6560
rect 3902 6496 3918 6560
rect 3982 6496 3998 6560
rect 4062 6496 4068 6560
rect 3752 6495 4068 6496
rect 10468 6560 10784 6561
rect 10468 6496 10474 6560
rect 10538 6496 10554 6560
rect 10618 6496 10634 6560
rect 10698 6496 10714 6560
rect 10778 6496 10784 6560
rect 10468 6495 10784 6496
rect 17184 6560 17500 6561
rect 17184 6496 17190 6560
rect 17254 6496 17270 6560
rect 17334 6496 17350 6560
rect 17414 6496 17430 6560
rect 17494 6496 17500 6560
rect 17184 6495 17500 6496
rect 23900 6560 24216 6561
rect 23900 6496 23906 6560
rect 23970 6496 23986 6560
rect 24050 6496 24066 6560
rect 24130 6496 24146 6560
rect 24210 6496 24216 6560
rect 23900 6495 24216 6496
rect 8109 6354 8175 6357
rect 9857 6354 9923 6357
rect 10174 6354 10180 6356
rect 8109 6352 10180 6354
rect 8109 6296 8114 6352
rect 8170 6296 9862 6352
rect 9918 6296 10180 6352
rect 8109 6294 10180 6296
rect 8109 6291 8175 6294
rect 9857 6291 9923 6294
rect 10174 6292 10180 6294
rect 10244 6292 10250 6356
rect 19425 6354 19491 6357
rect 12390 6352 19491 6354
rect 12390 6296 19430 6352
rect 19486 6296 19491 6352
rect 12390 6294 19491 6296
rect 12249 6218 12315 6221
rect 12390 6218 12450 6294
rect 19425 6291 19491 6294
rect 12249 6216 12450 6218
rect 12249 6160 12254 6216
rect 12310 6160 12450 6216
rect 12249 6158 12450 6160
rect 12249 6155 12315 6158
rect 7110 6016 7426 6017
rect 7110 5952 7116 6016
rect 7180 5952 7196 6016
rect 7260 5952 7276 6016
rect 7340 5952 7356 6016
rect 7420 5952 7426 6016
rect 7110 5951 7426 5952
rect 13826 6016 14142 6017
rect 13826 5952 13832 6016
rect 13896 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14142 6016
rect 13826 5951 14142 5952
rect 20542 6016 20858 6017
rect 20542 5952 20548 6016
rect 20612 5952 20628 6016
rect 20692 5952 20708 6016
rect 20772 5952 20788 6016
rect 20852 5952 20858 6016
rect 20542 5951 20858 5952
rect 27258 6016 27574 6017
rect 27258 5952 27264 6016
rect 27328 5952 27344 6016
rect 27408 5952 27424 6016
rect 27488 5952 27504 6016
rect 27568 5952 27574 6016
rect 27258 5951 27574 5952
rect 21541 5946 21607 5949
rect 22369 5946 22435 5949
rect 21541 5944 22435 5946
rect 21541 5888 21546 5944
rect 21602 5888 22374 5944
rect 22430 5888 22435 5944
rect 21541 5886 22435 5888
rect 21541 5883 21607 5886
rect 22369 5883 22435 5886
rect 6637 5674 6703 5677
rect 14457 5674 14523 5677
rect 6637 5672 14523 5674
rect 6637 5616 6642 5672
rect 6698 5616 14462 5672
rect 14518 5616 14523 5672
rect 6637 5614 14523 5616
rect 6637 5611 6703 5614
rect 14457 5611 14523 5614
rect 3752 5472 4068 5473
rect 3752 5408 3758 5472
rect 3822 5408 3838 5472
rect 3902 5408 3918 5472
rect 3982 5408 3998 5472
rect 4062 5408 4068 5472
rect 3752 5407 4068 5408
rect 10468 5472 10784 5473
rect 10468 5408 10474 5472
rect 10538 5408 10554 5472
rect 10618 5408 10634 5472
rect 10698 5408 10714 5472
rect 10778 5408 10784 5472
rect 10468 5407 10784 5408
rect 17184 5472 17500 5473
rect 17184 5408 17190 5472
rect 17254 5408 17270 5472
rect 17334 5408 17350 5472
rect 17414 5408 17430 5472
rect 17494 5408 17500 5472
rect 17184 5407 17500 5408
rect 23900 5472 24216 5473
rect 23900 5408 23906 5472
rect 23970 5408 23986 5472
rect 24050 5408 24066 5472
rect 24130 5408 24146 5472
rect 24210 5408 24216 5472
rect 23900 5407 24216 5408
rect 19425 5266 19491 5269
rect 20294 5266 20300 5268
rect 19425 5264 20300 5266
rect 19425 5208 19430 5264
rect 19486 5208 20300 5264
rect 19425 5206 20300 5208
rect 19425 5203 19491 5206
rect 20294 5204 20300 5206
rect 20364 5266 20370 5268
rect 21081 5266 21147 5269
rect 20364 5264 21147 5266
rect 20364 5208 21086 5264
rect 21142 5208 21147 5264
rect 20364 5206 21147 5208
rect 20364 5204 20370 5206
rect 21081 5203 21147 5206
rect 7110 4928 7426 4929
rect 7110 4864 7116 4928
rect 7180 4864 7196 4928
rect 7260 4864 7276 4928
rect 7340 4864 7356 4928
rect 7420 4864 7426 4928
rect 7110 4863 7426 4864
rect 13826 4928 14142 4929
rect 13826 4864 13832 4928
rect 13896 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14142 4928
rect 13826 4863 14142 4864
rect 20542 4928 20858 4929
rect 20542 4864 20548 4928
rect 20612 4864 20628 4928
rect 20692 4864 20708 4928
rect 20772 4864 20788 4928
rect 20852 4864 20858 4928
rect 20542 4863 20858 4864
rect 27258 4928 27574 4929
rect 27258 4864 27264 4928
rect 27328 4864 27344 4928
rect 27408 4864 27424 4928
rect 27488 4864 27504 4928
rect 27568 4864 27574 4928
rect 27258 4863 27574 4864
rect 17217 4722 17283 4725
rect 18137 4722 18203 4725
rect 17217 4720 18203 4722
rect 17217 4664 17222 4720
rect 17278 4664 18142 4720
rect 18198 4664 18203 4720
rect 17217 4662 18203 4664
rect 17217 4659 17283 4662
rect 18137 4659 18203 4662
rect 3752 4384 4068 4385
rect 3752 4320 3758 4384
rect 3822 4320 3838 4384
rect 3902 4320 3918 4384
rect 3982 4320 3998 4384
rect 4062 4320 4068 4384
rect 3752 4319 4068 4320
rect 10468 4384 10784 4385
rect 10468 4320 10474 4384
rect 10538 4320 10554 4384
rect 10618 4320 10634 4384
rect 10698 4320 10714 4384
rect 10778 4320 10784 4384
rect 10468 4319 10784 4320
rect 17184 4384 17500 4385
rect 17184 4320 17190 4384
rect 17254 4320 17270 4384
rect 17334 4320 17350 4384
rect 17414 4320 17430 4384
rect 17494 4320 17500 4384
rect 17184 4319 17500 4320
rect 23900 4384 24216 4385
rect 23900 4320 23906 4384
rect 23970 4320 23986 4384
rect 24050 4320 24066 4384
rect 24130 4320 24146 4384
rect 24210 4320 24216 4384
rect 23900 4319 24216 4320
rect 20069 4178 20135 4181
rect 24117 4178 24183 4181
rect 20069 4176 24183 4178
rect 20069 4120 20074 4176
rect 20130 4120 24122 4176
rect 24178 4120 24183 4176
rect 20069 4118 24183 4120
rect 20069 4115 20135 4118
rect 24117 4115 24183 4118
rect 18321 4044 18387 4045
rect 18270 3980 18276 4044
rect 18340 4042 18387 4044
rect 18340 4040 18432 4042
rect 18382 3984 18432 4040
rect 18340 3982 18432 3984
rect 18340 3980 18387 3982
rect 22318 3980 22324 4044
rect 22388 4042 22394 4044
rect 25313 4042 25379 4045
rect 22388 4040 25379 4042
rect 22388 3984 25318 4040
rect 25374 3984 25379 4040
rect 22388 3982 25379 3984
rect 22388 3980 22394 3982
rect 18321 3979 18387 3980
rect 25313 3979 25379 3982
rect 7110 3840 7426 3841
rect 7110 3776 7116 3840
rect 7180 3776 7196 3840
rect 7260 3776 7276 3840
rect 7340 3776 7356 3840
rect 7420 3776 7426 3840
rect 7110 3775 7426 3776
rect 13826 3840 14142 3841
rect 13826 3776 13832 3840
rect 13896 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14142 3840
rect 13826 3775 14142 3776
rect 20542 3840 20858 3841
rect 20542 3776 20548 3840
rect 20612 3776 20628 3840
rect 20692 3776 20708 3840
rect 20772 3776 20788 3840
rect 20852 3776 20858 3840
rect 20542 3775 20858 3776
rect 27258 3840 27574 3841
rect 27258 3776 27264 3840
rect 27328 3776 27344 3840
rect 27408 3776 27424 3840
rect 27488 3776 27504 3840
rect 27568 3776 27574 3840
rect 27258 3775 27574 3776
rect 22553 3770 22619 3773
rect 25589 3770 25655 3773
rect 22553 3768 25655 3770
rect 22553 3712 22558 3768
rect 22614 3712 25594 3768
rect 25650 3712 25655 3768
rect 22553 3710 25655 3712
rect 22553 3707 22619 3710
rect 25589 3707 25655 3710
rect 841 3498 907 3501
rect 14825 3498 14891 3501
rect 841 3496 14891 3498
rect 841 3440 846 3496
rect 902 3440 14830 3496
rect 14886 3440 14891 3496
rect 841 3438 14891 3440
rect 841 3435 907 3438
rect 14825 3435 14891 3438
rect 3752 3296 4068 3297
rect 3752 3232 3758 3296
rect 3822 3232 3838 3296
rect 3902 3232 3918 3296
rect 3982 3232 3998 3296
rect 4062 3232 4068 3296
rect 3752 3231 4068 3232
rect 10468 3296 10784 3297
rect 10468 3232 10474 3296
rect 10538 3232 10554 3296
rect 10618 3232 10634 3296
rect 10698 3232 10714 3296
rect 10778 3232 10784 3296
rect 10468 3231 10784 3232
rect 17184 3296 17500 3297
rect 17184 3232 17190 3296
rect 17254 3232 17270 3296
rect 17334 3232 17350 3296
rect 17414 3232 17430 3296
rect 17494 3232 17500 3296
rect 17184 3231 17500 3232
rect 23900 3296 24216 3297
rect 23900 3232 23906 3296
rect 23970 3232 23986 3296
rect 24050 3232 24066 3296
rect 24130 3232 24146 3296
rect 24210 3232 24216 3296
rect 23900 3231 24216 3232
rect 9857 2954 9923 2957
rect 13353 2954 13419 2957
rect 18229 2954 18295 2957
rect 9857 2952 18295 2954
rect 9857 2896 9862 2952
rect 9918 2896 13358 2952
rect 13414 2896 18234 2952
rect 18290 2896 18295 2952
rect 9857 2894 18295 2896
rect 9857 2891 9923 2894
rect 13353 2891 13419 2894
rect 18229 2891 18295 2894
rect 7110 2752 7426 2753
rect 7110 2688 7116 2752
rect 7180 2688 7196 2752
rect 7260 2688 7276 2752
rect 7340 2688 7356 2752
rect 7420 2688 7426 2752
rect 7110 2687 7426 2688
rect 13826 2752 14142 2753
rect 13826 2688 13832 2752
rect 13896 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14142 2752
rect 13826 2687 14142 2688
rect 20542 2752 20858 2753
rect 20542 2688 20548 2752
rect 20612 2688 20628 2752
rect 20692 2688 20708 2752
rect 20772 2688 20788 2752
rect 20852 2688 20858 2752
rect 20542 2687 20858 2688
rect 27258 2752 27574 2753
rect 27258 2688 27264 2752
rect 27328 2688 27344 2752
rect 27408 2688 27424 2752
rect 27488 2688 27504 2752
rect 27568 2688 27574 2752
rect 27258 2687 27574 2688
rect 13445 2546 13511 2549
rect 14089 2546 14155 2549
rect 13445 2544 14155 2546
rect 13445 2488 13450 2544
rect 13506 2488 14094 2544
rect 14150 2488 14155 2544
rect 13445 2486 14155 2488
rect 13445 2483 13511 2486
rect 14089 2483 14155 2486
rect 3752 2208 4068 2209
rect 3752 2144 3758 2208
rect 3822 2144 3838 2208
rect 3902 2144 3918 2208
rect 3982 2144 3998 2208
rect 4062 2144 4068 2208
rect 3752 2143 4068 2144
rect 10468 2208 10784 2209
rect 10468 2144 10474 2208
rect 10538 2144 10554 2208
rect 10618 2144 10634 2208
rect 10698 2144 10714 2208
rect 10778 2144 10784 2208
rect 10468 2143 10784 2144
rect 17184 2208 17500 2209
rect 17184 2144 17190 2208
rect 17254 2144 17270 2208
rect 17334 2144 17350 2208
rect 17414 2144 17430 2208
rect 17494 2144 17500 2208
rect 17184 2143 17500 2144
rect 23900 2208 24216 2209
rect 23900 2144 23906 2208
rect 23970 2144 23986 2208
rect 24050 2144 24066 2208
rect 24130 2144 24146 2208
rect 24210 2144 24216 2208
rect 23900 2143 24216 2144
rect 18413 2002 18479 2005
rect 19057 2002 19123 2005
rect 18413 2000 19123 2002
rect 18413 1944 18418 2000
rect 18474 1944 19062 2000
rect 19118 1944 19123 2000
rect 18413 1942 19123 1944
rect 18413 1939 18479 1942
rect 19057 1939 19123 1942
rect 17677 1866 17743 1869
rect 24209 1866 24275 1869
rect 17677 1864 24275 1866
rect 17677 1808 17682 1864
rect 17738 1808 24214 1864
rect 24270 1808 24275 1864
rect 17677 1806 24275 1808
rect 17677 1803 17743 1806
rect 24209 1803 24275 1806
rect 7110 1664 7426 1665
rect 7110 1600 7116 1664
rect 7180 1600 7196 1664
rect 7260 1600 7276 1664
rect 7340 1600 7356 1664
rect 7420 1600 7426 1664
rect 7110 1599 7426 1600
rect 13826 1664 14142 1665
rect 13826 1600 13832 1664
rect 13896 1600 13912 1664
rect 13976 1600 13992 1664
rect 14056 1600 14072 1664
rect 14136 1600 14142 1664
rect 13826 1599 14142 1600
rect 20542 1664 20858 1665
rect 20542 1600 20548 1664
rect 20612 1600 20628 1664
rect 20692 1600 20708 1664
rect 20772 1600 20788 1664
rect 20852 1600 20858 1664
rect 20542 1599 20858 1600
rect 27258 1664 27574 1665
rect 27258 1600 27264 1664
rect 27328 1600 27344 1664
rect 27408 1600 27424 1664
rect 27488 1600 27504 1664
rect 27568 1600 27574 1664
rect 27258 1599 27574 1600
rect 3752 1120 4068 1121
rect 3752 1056 3758 1120
rect 3822 1056 3838 1120
rect 3902 1056 3918 1120
rect 3982 1056 3998 1120
rect 4062 1056 4068 1120
rect 3752 1055 4068 1056
rect 10468 1120 10784 1121
rect 10468 1056 10474 1120
rect 10538 1056 10554 1120
rect 10618 1056 10634 1120
rect 10698 1056 10714 1120
rect 10778 1056 10784 1120
rect 10468 1055 10784 1056
rect 17184 1120 17500 1121
rect 17184 1056 17190 1120
rect 17254 1056 17270 1120
rect 17334 1056 17350 1120
rect 17414 1056 17430 1120
rect 17494 1056 17500 1120
rect 17184 1055 17500 1056
rect 23900 1120 24216 1121
rect 23900 1056 23906 1120
rect 23970 1056 23986 1120
rect 24050 1056 24066 1120
rect 24130 1056 24146 1120
rect 24210 1056 24216 1120
rect 23900 1055 24216 1056
rect 7110 576 7426 577
rect 7110 512 7116 576
rect 7180 512 7196 576
rect 7260 512 7276 576
rect 7340 512 7356 576
rect 7420 512 7426 576
rect 7110 511 7426 512
rect 13826 576 14142 577
rect 13826 512 13832 576
rect 13896 512 13912 576
rect 13976 512 13992 576
rect 14056 512 14072 576
rect 14136 512 14142 576
rect 13826 511 14142 512
rect 20542 576 20858 577
rect 20542 512 20548 576
rect 20612 512 20628 576
rect 20692 512 20708 576
rect 20772 512 20788 576
rect 20852 512 20858 576
rect 20542 511 20858 512
rect 27258 576 27574 577
rect 27258 512 27264 576
rect 27328 512 27344 576
rect 27408 512 27424 576
rect 27488 512 27504 576
rect 27568 512 27574 576
rect 27258 511 27574 512
<< via3 >>
rect 3758 17436 3822 17440
rect 3758 17380 3762 17436
rect 3762 17380 3818 17436
rect 3818 17380 3822 17436
rect 3758 17376 3822 17380
rect 3838 17436 3902 17440
rect 3838 17380 3842 17436
rect 3842 17380 3898 17436
rect 3898 17380 3902 17436
rect 3838 17376 3902 17380
rect 3918 17436 3982 17440
rect 3918 17380 3922 17436
rect 3922 17380 3978 17436
rect 3978 17380 3982 17436
rect 3918 17376 3982 17380
rect 3998 17436 4062 17440
rect 3998 17380 4002 17436
rect 4002 17380 4058 17436
rect 4058 17380 4062 17436
rect 3998 17376 4062 17380
rect 10474 17436 10538 17440
rect 10474 17380 10478 17436
rect 10478 17380 10534 17436
rect 10534 17380 10538 17436
rect 10474 17376 10538 17380
rect 10554 17436 10618 17440
rect 10554 17380 10558 17436
rect 10558 17380 10614 17436
rect 10614 17380 10618 17436
rect 10554 17376 10618 17380
rect 10634 17436 10698 17440
rect 10634 17380 10638 17436
rect 10638 17380 10694 17436
rect 10694 17380 10698 17436
rect 10634 17376 10698 17380
rect 10714 17436 10778 17440
rect 10714 17380 10718 17436
rect 10718 17380 10774 17436
rect 10774 17380 10778 17436
rect 10714 17376 10778 17380
rect 17190 17436 17254 17440
rect 17190 17380 17194 17436
rect 17194 17380 17250 17436
rect 17250 17380 17254 17436
rect 17190 17376 17254 17380
rect 17270 17436 17334 17440
rect 17270 17380 17274 17436
rect 17274 17380 17330 17436
rect 17330 17380 17334 17436
rect 17270 17376 17334 17380
rect 17350 17436 17414 17440
rect 17350 17380 17354 17436
rect 17354 17380 17410 17436
rect 17410 17380 17414 17436
rect 17350 17376 17414 17380
rect 17430 17436 17494 17440
rect 17430 17380 17434 17436
rect 17434 17380 17490 17436
rect 17490 17380 17494 17436
rect 17430 17376 17494 17380
rect 23906 17436 23970 17440
rect 23906 17380 23910 17436
rect 23910 17380 23966 17436
rect 23966 17380 23970 17436
rect 23906 17376 23970 17380
rect 23986 17436 24050 17440
rect 23986 17380 23990 17436
rect 23990 17380 24046 17436
rect 24046 17380 24050 17436
rect 23986 17376 24050 17380
rect 24066 17436 24130 17440
rect 24066 17380 24070 17436
rect 24070 17380 24126 17436
rect 24126 17380 24130 17436
rect 24066 17376 24130 17380
rect 24146 17436 24210 17440
rect 24146 17380 24150 17436
rect 24150 17380 24206 17436
rect 24206 17380 24210 17436
rect 24146 17376 24210 17380
rect 7116 16892 7180 16896
rect 7116 16836 7120 16892
rect 7120 16836 7176 16892
rect 7176 16836 7180 16892
rect 7116 16832 7180 16836
rect 7196 16892 7260 16896
rect 7196 16836 7200 16892
rect 7200 16836 7256 16892
rect 7256 16836 7260 16892
rect 7196 16832 7260 16836
rect 7276 16892 7340 16896
rect 7276 16836 7280 16892
rect 7280 16836 7336 16892
rect 7336 16836 7340 16892
rect 7276 16832 7340 16836
rect 7356 16892 7420 16896
rect 7356 16836 7360 16892
rect 7360 16836 7416 16892
rect 7416 16836 7420 16892
rect 7356 16832 7420 16836
rect 13832 16892 13896 16896
rect 13832 16836 13836 16892
rect 13836 16836 13892 16892
rect 13892 16836 13896 16892
rect 13832 16832 13896 16836
rect 13912 16892 13976 16896
rect 13912 16836 13916 16892
rect 13916 16836 13972 16892
rect 13972 16836 13976 16892
rect 13912 16832 13976 16836
rect 13992 16892 14056 16896
rect 13992 16836 13996 16892
rect 13996 16836 14052 16892
rect 14052 16836 14056 16892
rect 13992 16832 14056 16836
rect 14072 16892 14136 16896
rect 14072 16836 14076 16892
rect 14076 16836 14132 16892
rect 14132 16836 14136 16892
rect 14072 16832 14136 16836
rect 20548 16892 20612 16896
rect 20548 16836 20552 16892
rect 20552 16836 20608 16892
rect 20608 16836 20612 16892
rect 20548 16832 20612 16836
rect 20628 16892 20692 16896
rect 20628 16836 20632 16892
rect 20632 16836 20688 16892
rect 20688 16836 20692 16892
rect 20628 16832 20692 16836
rect 20708 16892 20772 16896
rect 20708 16836 20712 16892
rect 20712 16836 20768 16892
rect 20768 16836 20772 16892
rect 20708 16832 20772 16836
rect 20788 16892 20852 16896
rect 20788 16836 20792 16892
rect 20792 16836 20848 16892
rect 20848 16836 20852 16892
rect 20788 16832 20852 16836
rect 27264 16892 27328 16896
rect 27264 16836 27268 16892
rect 27268 16836 27324 16892
rect 27324 16836 27328 16892
rect 27264 16832 27328 16836
rect 27344 16892 27408 16896
rect 27344 16836 27348 16892
rect 27348 16836 27404 16892
rect 27404 16836 27408 16892
rect 27344 16832 27408 16836
rect 27424 16892 27488 16896
rect 27424 16836 27428 16892
rect 27428 16836 27484 16892
rect 27484 16836 27488 16892
rect 27424 16832 27488 16836
rect 27504 16892 27568 16896
rect 27504 16836 27508 16892
rect 27508 16836 27564 16892
rect 27564 16836 27568 16892
rect 27504 16832 27568 16836
rect 3758 16348 3822 16352
rect 3758 16292 3762 16348
rect 3762 16292 3818 16348
rect 3818 16292 3822 16348
rect 3758 16288 3822 16292
rect 3838 16348 3902 16352
rect 3838 16292 3842 16348
rect 3842 16292 3898 16348
rect 3898 16292 3902 16348
rect 3838 16288 3902 16292
rect 3918 16348 3982 16352
rect 3918 16292 3922 16348
rect 3922 16292 3978 16348
rect 3978 16292 3982 16348
rect 3918 16288 3982 16292
rect 3998 16348 4062 16352
rect 3998 16292 4002 16348
rect 4002 16292 4058 16348
rect 4058 16292 4062 16348
rect 3998 16288 4062 16292
rect 10474 16348 10538 16352
rect 10474 16292 10478 16348
rect 10478 16292 10534 16348
rect 10534 16292 10538 16348
rect 10474 16288 10538 16292
rect 10554 16348 10618 16352
rect 10554 16292 10558 16348
rect 10558 16292 10614 16348
rect 10614 16292 10618 16348
rect 10554 16288 10618 16292
rect 10634 16348 10698 16352
rect 10634 16292 10638 16348
rect 10638 16292 10694 16348
rect 10694 16292 10698 16348
rect 10634 16288 10698 16292
rect 10714 16348 10778 16352
rect 10714 16292 10718 16348
rect 10718 16292 10774 16348
rect 10774 16292 10778 16348
rect 10714 16288 10778 16292
rect 17190 16348 17254 16352
rect 17190 16292 17194 16348
rect 17194 16292 17250 16348
rect 17250 16292 17254 16348
rect 17190 16288 17254 16292
rect 17270 16348 17334 16352
rect 17270 16292 17274 16348
rect 17274 16292 17330 16348
rect 17330 16292 17334 16348
rect 17270 16288 17334 16292
rect 17350 16348 17414 16352
rect 17350 16292 17354 16348
rect 17354 16292 17410 16348
rect 17410 16292 17414 16348
rect 17350 16288 17414 16292
rect 17430 16348 17494 16352
rect 17430 16292 17434 16348
rect 17434 16292 17490 16348
rect 17490 16292 17494 16348
rect 17430 16288 17494 16292
rect 23906 16348 23970 16352
rect 23906 16292 23910 16348
rect 23910 16292 23966 16348
rect 23966 16292 23970 16348
rect 23906 16288 23970 16292
rect 23986 16348 24050 16352
rect 23986 16292 23990 16348
rect 23990 16292 24046 16348
rect 24046 16292 24050 16348
rect 23986 16288 24050 16292
rect 24066 16348 24130 16352
rect 24066 16292 24070 16348
rect 24070 16292 24126 16348
rect 24126 16292 24130 16348
rect 24066 16288 24130 16292
rect 24146 16348 24210 16352
rect 24146 16292 24150 16348
rect 24150 16292 24206 16348
rect 24206 16292 24210 16348
rect 24146 16288 24210 16292
rect 7116 15804 7180 15808
rect 7116 15748 7120 15804
rect 7120 15748 7176 15804
rect 7176 15748 7180 15804
rect 7116 15744 7180 15748
rect 7196 15804 7260 15808
rect 7196 15748 7200 15804
rect 7200 15748 7256 15804
rect 7256 15748 7260 15804
rect 7196 15744 7260 15748
rect 7276 15804 7340 15808
rect 7276 15748 7280 15804
rect 7280 15748 7336 15804
rect 7336 15748 7340 15804
rect 7276 15744 7340 15748
rect 7356 15804 7420 15808
rect 7356 15748 7360 15804
rect 7360 15748 7416 15804
rect 7416 15748 7420 15804
rect 7356 15744 7420 15748
rect 13832 15804 13896 15808
rect 13832 15748 13836 15804
rect 13836 15748 13892 15804
rect 13892 15748 13896 15804
rect 13832 15744 13896 15748
rect 13912 15804 13976 15808
rect 13912 15748 13916 15804
rect 13916 15748 13972 15804
rect 13972 15748 13976 15804
rect 13912 15744 13976 15748
rect 13992 15804 14056 15808
rect 13992 15748 13996 15804
rect 13996 15748 14052 15804
rect 14052 15748 14056 15804
rect 13992 15744 14056 15748
rect 14072 15804 14136 15808
rect 14072 15748 14076 15804
rect 14076 15748 14132 15804
rect 14132 15748 14136 15804
rect 14072 15744 14136 15748
rect 20548 15804 20612 15808
rect 20548 15748 20552 15804
rect 20552 15748 20608 15804
rect 20608 15748 20612 15804
rect 20548 15744 20612 15748
rect 20628 15804 20692 15808
rect 20628 15748 20632 15804
rect 20632 15748 20688 15804
rect 20688 15748 20692 15804
rect 20628 15744 20692 15748
rect 20708 15804 20772 15808
rect 20708 15748 20712 15804
rect 20712 15748 20768 15804
rect 20768 15748 20772 15804
rect 20708 15744 20772 15748
rect 20788 15804 20852 15808
rect 20788 15748 20792 15804
rect 20792 15748 20848 15804
rect 20848 15748 20852 15804
rect 20788 15744 20852 15748
rect 27264 15804 27328 15808
rect 27264 15748 27268 15804
rect 27268 15748 27324 15804
rect 27324 15748 27328 15804
rect 27264 15744 27328 15748
rect 27344 15804 27408 15808
rect 27344 15748 27348 15804
rect 27348 15748 27404 15804
rect 27404 15748 27408 15804
rect 27344 15744 27408 15748
rect 27424 15804 27488 15808
rect 27424 15748 27428 15804
rect 27428 15748 27484 15804
rect 27484 15748 27488 15804
rect 27424 15744 27488 15748
rect 27504 15804 27568 15808
rect 27504 15748 27508 15804
rect 27508 15748 27564 15804
rect 27564 15748 27568 15804
rect 27504 15744 27568 15748
rect 17724 15404 17788 15468
rect 3758 15260 3822 15264
rect 3758 15204 3762 15260
rect 3762 15204 3818 15260
rect 3818 15204 3822 15260
rect 3758 15200 3822 15204
rect 3838 15260 3902 15264
rect 3838 15204 3842 15260
rect 3842 15204 3898 15260
rect 3898 15204 3902 15260
rect 3838 15200 3902 15204
rect 3918 15260 3982 15264
rect 3918 15204 3922 15260
rect 3922 15204 3978 15260
rect 3978 15204 3982 15260
rect 3918 15200 3982 15204
rect 3998 15260 4062 15264
rect 3998 15204 4002 15260
rect 4002 15204 4058 15260
rect 4058 15204 4062 15260
rect 3998 15200 4062 15204
rect 10474 15260 10538 15264
rect 10474 15204 10478 15260
rect 10478 15204 10534 15260
rect 10534 15204 10538 15260
rect 10474 15200 10538 15204
rect 10554 15260 10618 15264
rect 10554 15204 10558 15260
rect 10558 15204 10614 15260
rect 10614 15204 10618 15260
rect 10554 15200 10618 15204
rect 10634 15260 10698 15264
rect 10634 15204 10638 15260
rect 10638 15204 10694 15260
rect 10694 15204 10698 15260
rect 10634 15200 10698 15204
rect 10714 15260 10778 15264
rect 10714 15204 10718 15260
rect 10718 15204 10774 15260
rect 10774 15204 10778 15260
rect 10714 15200 10778 15204
rect 17190 15260 17254 15264
rect 17190 15204 17194 15260
rect 17194 15204 17250 15260
rect 17250 15204 17254 15260
rect 17190 15200 17254 15204
rect 17270 15260 17334 15264
rect 17270 15204 17274 15260
rect 17274 15204 17330 15260
rect 17330 15204 17334 15260
rect 17270 15200 17334 15204
rect 17350 15260 17414 15264
rect 17350 15204 17354 15260
rect 17354 15204 17410 15260
rect 17410 15204 17414 15260
rect 17350 15200 17414 15204
rect 17430 15260 17494 15264
rect 17430 15204 17434 15260
rect 17434 15204 17490 15260
rect 17490 15204 17494 15260
rect 17430 15200 17494 15204
rect 23906 15260 23970 15264
rect 23906 15204 23910 15260
rect 23910 15204 23966 15260
rect 23966 15204 23970 15260
rect 23906 15200 23970 15204
rect 23986 15260 24050 15264
rect 23986 15204 23990 15260
rect 23990 15204 24046 15260
rect 24046 15204 24050 15260
rect 23986 15200 24050 15204
rect 24066 15260 24130 15264
rect 24066 15204 24070 15260
rect 24070 15204 24126 15260
rect 24126 15204 24130 15260
rect 24066 15200 24130 15204
rect 24146 15260 24210 15264
rect 24146 15204 24150 15260
rect 24150 15204 24206 15260
rect 24206 15204 24210 15260
rect 24146 15200 24210 15204
rect 7116 14716 7180 14720
rect 7116 14660 7120 14716
rect 7120 14660 7176 14716
rect 7176 14660 7180 14716
rect 7116 14656 7180 14660
rect 7196 14716 7260 14720
rect 7196 14660 7200 14716
rect 7200 14660 7256 14716
rect 7256 14660 7260 14716
rect 7196 14656 7260 14660
rect 7276 14716 7340 14720
rect 7276 14660 7280 14716
rect 7280 14660 7336 14716
rect 7336 14660 7340 14716
rect 7276 14656 7340 14660
rect 7356 14716 7420 14720
rect 7356 14660 7360 14716
rect 7360 14660 7416 14716
rect 7416 14660 7420 14716
rect 7356 14656 7420 14660
rect 13832 14716 13896 14720
rect 13832 14660 13836 14716
rect 13836 14660 13892 14716
rect 13892 14660 13896 14716
rect 13832 14656 13896 14660
rect 13912 14716 13976 14720
rect 13912 14660 13916 14716
rect 13916 14660 13972 14716
rect 13972 14660 13976 14716
rect 13912 14656 13976 14660
rect 13992 14716 14056 14720
rect 13992 14660 13996 14716
rect 13996 14660 14052 14716
rect 14052 14660 14056 14716
rect 13992 14656 14056 14660
rect 14072 14716 14136 14720
rect 14072 14660 14076 14716
rect 14076 14660 14132 14716
rect 14132 14660 14136 14716
rect 14072 14656 14136 14660
rect 20548 14716 20612 14720
rect 20548 14660 20552 14716
rect 20552 14660 20608 14716
rect 20608 14660 20612 14716
rect 20548 14656 20612 14660
rect 20628 14716 20692 14720
rect 20628 14660 20632 14716
rect 20632 14660 20688 14716
rect 20688 14660 20692 14716
rect 20628 14656 20692 14660
rect 20708 14716 20772 14720
rect 20708 14660 20712 14716
rect 20712 14660 20768 14716
rect 20768 14660 20772 14716
rect 20708 14656 20772 14660
rect 20788 14716 20852 14720
rect 20788 14660 20792 14716
rect 20792 14660 20848 14716
rect 20848 14660 20852 14716
rect 20788 14656 20852 14660
rect 27264 14716 27328 14720
rect 27264 14660 27268 14716
rect 27268 14660 27324 14716
rect 27324 14660 27328 14716
rect 27264 14656 27328 14660
rect 27344 14716 27408 14720
rect 27344 14660 27348 14716
rect 27348 14660 27404 14716
rect 27404 14660 27408 14716
rect 27344 14656 27408 14660
rect 27424 14716 27488 14720
rect 27424 14660 27428 14716
rect 27428 14660 27484 14716
rect 27484 14660 27488 14716
rect 27424 14656 27488 14660
rect 27504 14716 27568 14720
rect 27504 14660 27508 14716
rect 27508 14660 27564 14716
rect 27564 14660 27568 14716
rect 27504 14656 27568 14660
rect 3758 14172 3822 14176
rect 3758 14116 3762 14172
rect 3762 14116 3818 14172
rect 3818 14116 3822 14172
rect 3758 14112 3822 14116
rect 3838 14172 3902 14176
rect 3838 14116 3842 14172
rect 3842 14116 3898 14172
rect 3898 14116 3902 14172
rect 3838 14112 3902 14116
rect 3918 14172 3982 14176
rect 3918 14116 3922 14172
rect 3922 14116 3978 14172
rect 3978 14116 3982 14172
rect 3918 14112 3982 14116
rect 3998 14172 4062 14176
rect 3998 14116 4002 14172
rect 4002 14116 4058 14172
rect 4058 14116 4062 14172
rect 3998 14112 4062 14116
rect 10474 14172 10538 14176
rect 10474 14116 10478 14172
rect 10478 14116 10534 14172
rect 10534 14116 10538 14172
rect 10474 14112 10538 14116
rect 10554 14172 10618 14176
rect 10554 14116 10558 14172
rect 10558 14116 10614 14172
rect 10614 14116 10618 14172
rect 10554 14112 10618 14116
rect 10634 14172 10698 14176
rect 10634 14116 10638 14172
rect 10638 14116 10694 14172
rect 10694 14116 10698 14172
rect 10634 14112 10698 14116
rect 10714 14172 10778 14176
rect 10714 14116 10718 14172
rect 10718 14116 10774 14172
rect 10774 14116 10778 14172
rect 10714 14112 10778 14116
rect 17190 14172 17254 14176
rect 17190 14116 17194 14172
rect 17194 14116 17250 14172
rect 17250 14116 17254 14172
rect 17190 14112 17254 14116
rect 17270 14172 17334 14176
rect 17270 14116 17274 14172
rect 17274 14116 17330 14172
rect 17330 14116 17334 14172
rect 17270 14112 17334 14116
rect 17350 14172 17414 14176
rect 17350 14116 17354 14172
rect 17354 14116 17410 14172
rect 17410 14116 17414 14172
rect 17350 14112 17414 14116
rect 17430 14172 17494 14176
rect 17430 14116 17434 14172
rect 17434 14116 17490 14172
rect 17490 14116 17494 14172
rect 17430 14112 17494 14116
rect 23906 14172 23970 14176
rect 23906 14116 23910 14172
rect 23910 14116 23966 14172
rect 23966 14116 23970 14172
rect 23906 14112 23970 14116
rect 23986 14172 24050 14176
rect 23986 14116 23990 14172
rect 23990 14116 24046 14172
rect 24046 14116 24050 14172
rect 23986 14112 24050 14116
rect 24066 14172 24130 14176
rect 24066 14116 24070 14172
rect 24070 14116 24126 14172
rect 24126 14116 24130 14172
rect 24066 14112 24130 14116
rect 24146 14172 24210 14176
rect 24146 14116 24150 14172
rect 24150 14116 24206 14172
rect 24206 14116 24210 14172
rect 24146 14112 24210 14116
rect 22324 13832 22388 13836
rect 22324 13776 22374 13832
rect 22374 13776 22388 13832
rect 22324 13772 22388 13776
rect 7116 13628 7180 13632
rect 7116 13572 7120 13628
rect 7120 13572 7176 13628
rect 7176 13572 7180 13628
rect 7116 13568 7180 13572
rect 7196 13628 7260 13632
rect 7196 13572 7200 13628
rect 7200 13572 7256 13628
rect 7256 13572 7260 13628
rect 7196 13568 7260 13572
rect 7276 13628 7340 13632
rect 7276 13572 7280 13628
rect 7280 13572 7336 13628
rect 7336 13572 7340 13628
rect 7276 13568 7340 13572
rect 7356 13628 7420 13632
rect 7356 13572 7360 13628
rect 7360 13572 7416 13628
rect 7416 13572 7420 13628
rect 7356 13568 7420 13572
rect 13832 13628 13896 13632
rect 13832 13572 13836 13628
rect 13836 13572 13892 13628
rect 13892 13572 13896 13628
rect 13832 13568 13896 13572
rect 13912 13628 13976 13632
rect 13912 13572 13916 13628
rect 13916 13572 13972 13628
rect 13972 13572 13976 13628
rect 13912 13568 13976 13572
rect 13992 13628 14056 13632
rect 13992 13572 13996 13628
rect 13996 13572 14052 13628
rect 14052 13572 14056 13628
rect 13992 13568 14056 13572
rect 14072 13628 14136 13632
rect 14072 13572 14076 13628
rect 14076 13572 14132 13628
rect 14132 13572 14136 13628
rect 14072 13568 14136 13572
rect 20548 13628 20612 13632
rect 20548 13572 20552 13628
rect 20552 13572 20608 13628
rect 20608 13572 20612 13628
rect 20548 13568 20612 13572
rect 20628 13628 20692 13632
rect 20628 13572 20632 13628
rect 20632 13572 20688 13628
rect 20688 13572 20692 13628
rect 20628 13568 20692 13572
rect 20708 13628 20772 13632
rect 20708 13572 20712 13628
rect 20712 13572 20768 13628
rect 20768 13572 20772 13628
rect 20708 13568 20772 13572
rect 20788 13628 20852 13632
rect 20788 13572 20792 13628
rect 20792 13572 20848 13628
rect 20848 13572 20852 13628
rect 20788 13568 20852 13572
rect 27264 13628 27328 13632
rect 27264 13572 27268 13628
rect 27268 13572 27324 13628
rect 27324 13572 27328 13628
rect 27264 13568 27328 13572
rect 27344 13628 27408 13632
rect 27344 13572 27348 13628
rect 27348 13572 27404 13628
rect 27404 13572 27408 13628
rect 27344 13568 27408 13572
rect 27424 13628 27488 13632
rect 27424 13572 27428 13628
rect 27428 13572 27484 13628
rect 27484 13572 27488 13628
rect 27424 13568 27488 13572
rect 27504 13628 27568 13632
rect 27504 13572 27508 13628
rect 27508 13572 27564 13628
rect 27564 13572 27568 13628
rect 27504 13568 27568 13572
rect 3758 13084 3822 13088
rect 3758 13028 3762 13084
rect 3762 13028 3818 13084
rect 3818 13028 3822 13084
rect 3758 13024 3822 13028
rect 3838 13084 3902 13088
rect 3838 13028 3842 13084
rect 3842 13028 3898 13084
rect 3898 13028 3902 13084
rect 3838 13024 3902 13028
rect 3918 13084 3982 13088
rect 3918 13028 3922 13084
rect 3922 13028 3978 13084
rect 3978 13028 3982 13084
rect 3918 13024 3982 13028
rect 3998 13084 4062 13088
rect 3998 13028 4002 13084
rect 4002 13028 4058 13084
rect 4058 13028 4062 13084
rect 3998 13024 4062 13028
rect 10474 13084 10538 13088
rect 10474 13028 10478 13084
rect 10478 13028 10534 13084
rect 10534 13028 10538 13084
rect 10474 13024 10538 13028
rect 10554 13084 10618 13088
rect 10554 13028 10558 13084
rect 10558 13028 10614 13084
rect 10614 13028 10618 13084
rect 10554 13024 10618 13028
rect 10634 13084 10698 13088
rect 10634 13028 10638 13084
rect 10638 13028 10694 13084
rect 10694 13028 10698 13084
rect 10634 13024 10698 13028
rect 10714 13084 10778 13088
rect 10714 13028 10718 13084
rect 10718 13028 10774 13084
rect 10774 13028 10778 13084
rect 10714 13024 10778 13028
rect 17190 13084 17254 13088
rect 17190 13028 17194 13084
rect 17194 13028 17250 13084
rect 17250 13028 17254 13084
rect 17190 13024 17254 13028
rect 17270 13084 17334 13088
rect 17270 13028 17274 13084
rect 17274 13028 17330 13084
rect 17330 13028 17334 13084
rect 17270 13024 17334 13028
rect 17350 13084 17414 13088
rect 17350 13028 17354 13084
rect 17354 13028 17410 13084
rect 17410 13028 17414 13084
rect 17350 13024 17414 13028
rect 17430 13084 17494 13088
rect 17430 13028 17434 13084
rect 17434 13028 17490 13084
rect 17490 13028 17494 13084
rect 17430 13024 17494 13028
rect 23906 13084 23970 13088
rect 23906 13028 23910 13084
rect 23910 13028 23966 13084
rect 23966 13028 23970 13084
rect 23906 13024 23970 13028
rect 23986 13084 24050 13088
rect 23986 13028 23990 13084
rect 23990 13028 24046 13084
rect 24046 13028 24050 13084
rect 23986 13024 24050 13028
rect 24066 13084 24130 13088
rect 24066 13028 24070 13084
rect 24070 13028 24126 13084
rect 24126 13028 24130 13084
rect 24066 13024 24130 13028
rect 24146 13084 24210 13088
rect 24146 13028 24150 13084
rect 24150 13028 24206 13084
rect 24206 13028 24210 13084
rect 24146 13024 24210 13028
rect 17724 12548 17788 12612
rect 7116 12540 7180 12544
rect 7116 12484 7120 12540
rect 7120 12484 7176 12540
rect 7176 12484 7180 12540
rect 7116 12480 7180 12484
rect 7196 12540 7260 12544
rect 7196 12484 7200 12540
rect 7200 12484 7256 12540
rect 7256 12484 7260 12540
rect 7196 12480 7260 12484
rect 7276 12540 7340 12544
rect 7276 12484 7280 12540
rect 7280 12484 7336 12540
rect 7336 12484 7340 12540
rect 7276 12480 7340 12484
rect 7356 12540 7420 12544
rect 7356 12484 7360 12540
rect 7360 12484 7416 12540
rect 7416 12484 7420 12540
rect 7356 12480 7420 12484
rect 13832 12540 13896 12544
rect 13832 12484 13836 12540
rect 13836 12484 13892 12540
rect 13892 12484 13896 12540
rect 13832 12480 13896 12484
rect 13912 12540 13976 12544
rect 13912 12484 13916 12540
rect 13916 12484 13972 12540
rect 13972 12484 13976 12540
rect 13912 12480 13976 12484
rect 13992 12540 14056 12544
rect 13992 12484 13996 12540
rect 13996 12484 14052 12540
rect 14052 12484 14056 12540
rect 13992 12480 14056 12484
rect 14072 12540 14136 12544
rect 14072 12484 14076 12540
rect 14076 12484 14132 12540
rect 14132 12484 14136 12540
rect 14072 12480 14136 12484
rect 20548 12540 20612 12544
rect 20548 12484 20552 12540
rect 20552 12484 20608 12540
rect 20608 12484 20612 12540
rect 20548 12480 20612 12484
rect 20628 12540 20692 12544
rect 20628 12484 20632 12540
rect 20632 12484 20688 12540
rect 20688 12484 20692 12540
rect 20628 12480 20692 12484
rect 20708 12540 20772 12544
rect 20708 12484 20712 12540
rect 20712 12484 20768 12540
rect 20768 12484 20772 12540
rect 20708 12480 20772 12484
rect 20788 12540 20852 12544
rect 20788 12484 20792 12540
rect 20792 12484 20848 12540
rect 20848 12484 20852 12540
rect 20788 12480 20852 12484
rect 27264 12540 27328 12544
rect 27264 12484 27268 12540
rect 27268 12484 27324 12540
rect 27324 12484 27328 12540
rect 27264 12480 27328 12484
rect 27344 12540 27408 12544
rect 27344 12484 27348 12540
rect 27348 12484 27404 12540
rect 27404 12484 27408 12540
rect 27344 12480 27408 12484
rect 27424 12540 27488 12544
rect 27424 12484 27428 12540
rect 27428 12484 27484 12540
rect 27484 12484 27488 12540
rect 27424 12480 27488 12484
rect 27504 12540 27568 12544
rect 27504 12484 27508 12540
rect 27508 12484 27564 12540
rect 27564 12484 27568 12540
rect 27504 12480 27568 12484
rect 26188 12336 26252 12340
rect 26188 12280 26202 12336
rect 26202 12280 26252 12336
rect 26188 12276 26252 12280
rect 10180 12140 10244 12204
rect 3758 11996 3822 12000
rect 3758 11940 3762 11996
rect 3762 11940 3818 11996
rect 3818 11940 3822 11996
rect 3758 11936 3822 11940
rect 3838 11996 3902 12000
rect 3838 11940 3842 11996
rect 3842 11940 3898 11996
rect 3898 11940 3902 11996
rect 3838 11936 3902 11940
rect 3918 11996 3982 12000
rect 3918 11940 3922 11996
rect 3922 11940 3978 11996
rect 3978 11940 3982 11996
rect 3918 11936 3982 11940
rect 3998 11996 4062 12000
rect 3998 11940 4002 11996
rect 4002 11940 4058 11996
rect 4058 11940 4062 11996
rect 3998 11936 4062 11940
rect 10474 11996 10538 12000
rect 10474 11940 10478 11996
rect 10478 11940 10534 11996
rect 10534 11940 10538 11996
rect 10474 11936 10538 11940
rect 10554 11996 10618 12000
rect 10554 11940 10558 11996
rect 10558 11940 10614 11996
rect 10614 11940 10618 11996
rect 10554 11936 10618 11940
rect 10634 11996 10698 12000
rect 10634 11940 10638 11996
rect 10638 11940 10694 11996
rect 10694 11940 10698 11996
rect 10634 11936 10698 11940
rect 10714 11996 10778 12000
rect 10714 11940 10718 11996
rect 10718 11940 10774 11996
rect 10774 11940 10778 11996
rect 10714 11936 10778 11940
rect 17190 11996 17254 12000
rect 17190 11940 17194 11996
rect 17194 11940 17250 11996
rect 17250 11940 17254 11996
rect 17190 11936 17254 11940
rect 17270 11996 17334 12000
rect 17270 11940 17274 11996
rect 17274 11940 17330 11996
rect 17330 11940 17334 11996
rect 17270 11936 17334 11940
rect 17350 11996 17414 12000
rect 17350 11940 17354 11996
rect 17354 11940 17410 11996
rect 17410 11940 17414 11996
rect 17350 11936 17414 11940
rect 17430 11996 17494 12000
rect 17430 11940 17434 11996
rect 17434 11940 17490 11996
rect 17490 11940 17494 11996
rect 17430 11936 17494 11940
rect 23906 11996 23970 12000
rect 23906 11940 23910 11996
rect 23910 11940 23966 11996
rect 23966 11940 23970 11996
rect 23906 11936 23970 11940
rect 23986 11996 24050 12000
rect 23986 11940 23990 11996
rect 23990 11940 24046 11996
rect 24046 11940 24050 11996
rect 23986 11936 24050 11940
rect 24066 11996 24130 12000
rect 24066 11940 24070 11996
rect 24070 11940 24126 11996
rect 24126 11940 24130 11996
rect 24066 11936 24130 11940
rect 24146 11996 24210 12000
rect 24146 11940 24150 11996
rect 24150 11940 24206 11996
rect 24206 11940 24210 11996
rect 24146 11936 24210 11940
rect 18644 11520 18708 11524
rect 18644 11464 18694 11520
rect 18694 11464 18708 11520
rect 18644 11460 18708 11464
rect 7116 11452 7180 11456
rect 7116 11396 7120 11452
rect 7120 11396 7176 11452
rect 7176 11396 7180 11452
rect 7116 11392 7180 11396
rect 7196 11452 7260 11456
rect 7196 11396 7200 11452
rect 7200 11396 7256 11452
rect 7256 11396 7260 11452
rect 7196 11392 7260 11396
rect 7276 11452 7340 11456
rect 7276 11396 7280 11452
rect 7280 11396 7336 11452
rect 7336 11396 7340 11452
rect 7276 11392 7340 11396
rect 7356 11452 7420 11456
rect 7356 11396 7360 11452
rect 7360 11396 7416 11452
rect 7416 11396 7420 11452
rect 7356 11392 7420 11396
rect 13832 11452 13896 11456
rect 13832 11396 13836 11452
rect 13836 11396 13892 11452
rect 13892 11396 13896 11452
rect 13832 11392 13896 11396
rect 13912 11452 13976 11456
rect 13912 11396 13916 11452
rect 13916 11396 13972 11452
rect 13972 11396 13976 11452
rect 13912 11392 13976 11396
rect 13992 11452 14056 11456
rect 13992 11396 13996 11452
rect 13996 11396 14052 11452
rect 14052 11396 14056 11452
rect 13992 11392 14056 11396
rect 14072 11452 14136 11456
rect 14072 11396 14076 11452
rect 14076 11396 14132 11452
rect 14132 11396 14136 11452
rect 14072 11392 14136 11396
rect 20548 11452 20612 11456
rect 20548 11396 20552 11452
rect 20552 11396 20608 11452
rect 20608 11396 20612 11452
rect 20548 11392 20612 11396
rect 20628 11452 20692 11456
rect 20628 11396 20632 11452
rect 20632 11396 20688 11452
rect 20688 11396 20692 11452
rect 20628 11392 20692 11396
rect 20708 11452 20772 11456
rect 20708 11396 20712 11452
rect 20712 11396 20768 11452
rect 20768 11396 20772 11452
rect 20708 11392 20772 11396
rect 20788 11452 20852 11456
rect 20788 11396 20792 11452
rect 20792 11396 20848 11452
rect 20848 11396 20852 11452
rect 20788 11392 20852 11396
rect 27264 11452 27328 11456
rect 27264 11396 27268 11452
rect 27268 11396 27324 11452
rect 27324 11396 27328 11452
rect 27264 11392 27328 11396
rect 27344 11452 27408 11456
rect 27344 11396 27348 11452
rect 27348 11396 27404 11452
rect 27404 11396 27408 11452
rect 27344 11392 27408 11396
rect 27424 11452 27488 11456
rect 27424 11396 27428 11452
rect 27428 11396 27484 11452
rect 27484 11396 27488 11452
rect 27424 11392 27488 11396
rect 27504 11452 27568 11456
rect 27504 11396 27508 11452
rect 27508 11396 27564 11452
rect 27564 11396 27568 11452
rect 27504 11392 27568 11396
rect 18276 11052 18340 11116
rect 3758 10908 3822 10912
rect 3758 10852 3762 10908
rect 3762 10852 3818 10908
rect 3818 10852 3822 10908
rect 3758 10848 3822 10852
rect 3838 10908 3902 10912
rect 3838 10852 3842 10908
rect 3842 10852 3898 10908
rect 3898 10852 3902 10908
rect 3838 10848 3902 10852
rect 3918 10908 3982 10912
rect 3918 10852 3922 10908
rect 3922 10852 3978 10908
rect 3978 10852 3982 10908
rect 3918 10848 3982 10852
rect 3998 10908 4062 10912
rect 3998 10852 4002 10908
rect 4002 10852 4058 10908
rect 4058 10852 4062 10908
rect 3998 10848 4062 10852
rect 10474 10908 10538 10912
rect 10474 10852 10478 10908
rect 10478 10852 10534 10908
rect 10534 10852 10538 10908
rect 10474 10848 10538 10852
rect 10554 10908 10618 10912
rect 10554 10852 10558 10908
rect 10558 10852 10614 10908
rect 10614 10852 10618 10908
rect 10554 10848 10618 10852
rect 10634 10908 10698 10912
rect 10634 10852 10638 10908
rect 10638 10852 10694 10908
rect 10694 10852 10698 10908
rect 10634 10848 10698 10852
rect 10714 10908 10778 10912
rect 10714 10852 10718 10908
rect 10718 10852 10774 10908
rect 10774 10852 10778 10908
rect 10714 10848 10778 10852
rect 17190 10908 17254 10912
rect 17190 10852 17194 10908
rect 17194 10852 17250 10908
rect 17250 10852 17254 10908
rect 17190 10848 17254 10852
rect 17270 10908 17334 10912
rect 17270 10852 17274 10908
rect 17274 10852 17330 10908
rect 17330 10852 17334 10908
rect 17270 10848 17334 10852
rect 17350 10908 17414 10912
rect 17350 10852 17354 10908
rect 17354 10852 17410 10908
rect 17410 10852 17414 10908
rect 17350 10848 17414 10852
rect 17430 10908 17494 10912
rect 17430 10852 17434 10908
rect 17434 10852 17490 10908
rect 17490 10852 17494 10908
rect 17430 10848 17494 10852
rect 23906 10908 23970 10912
rect 23906 10852 23910 10908
rect 23910 10852 23966 10908
rect 23966 10852 23970 10908
rect 23906 10848 23970 10852
rect 23986 10908 24050 10912
rect 23986 10852 23990 10908
rect 23990 10852 24046 10908
rect 24046 10852 24050 10908
rect 23986 10848 24050 10852
rect 24066 10908 24130 10912
rect 24066 10852 24070 10908
rect 24070 10852 24126 10908
rect 24126 10852 24130 10908
rect 24066 10848 24130 10852
rect 24146 10908 24210 10912
rect 24146 10852 24150 10908
rect 24150 10852 24206 10908
rect 24206 10852 24210 10908
rect 24146 10848 24210 10852
rect 7116 10364 7180 10368
rect 7116 10308 7120 10364
rect 7120 10308 7176 10364
rect 7176 10308 7180 10364
rect 7116 10304 7180 10308
rect 7196 10364 7260 10368
rect 7196 10308 7200 10364
rect 7200 10308 7256 10364
rect 7256 10308 7260 10364
rect 7196 10304 7260 10308
rect 7276 10364 7340 10368
rect 7276 10308 7280 10364
rect 7280 10308 7336 10364
rect 7336 10308 7340 10364
rect 7276 10304 7340 10308
rect 7356 10364 7420 10368
rect 7356 10308 7360 10364
rect 7360 10308 7416 10364
rect 7416 10308 7420 10364
rect 7356 10304 7420 10308
rect 13832 10364 13896 10368
rect 13832 10308 13836 10364
rect 13836 10308 13892 10364
rect 13892 10308 13896 10364
rect 13832 10304 13896 10308
rect 13912 10364 13976 10368
rect 13912 10308 13916 10364
rect 13916 10308 13972 10364
rect 13972 10308 13976 10364
rect 13912 10304 13976 10308
rect 13992 10364 14056 10368
rect 13992 10308 13996 10364
rect 13996 10308 14052 10364
rect 14052 10308 14056 10364
rect 13992 10304 14056 10308
rect 14072 10364 14136 10368
rect 14072 10308 14076 10364
rect 14076 10308 14132 10364
rect 14132 10308 14136 10364
rect 14072 10304 14136 10308
rect 20548 10364 20612 10368
rect 20548 10308 20552 10364
rect 20552 10308 20608 10364
rect 20608 10308 20612 10364
rect 20548 10304 20612 10308
rect 20628 10364 20692 10368
rect 20628 10308 20632 10364
rect 20632 10308 20688 10364
rect 20688 10308 20692 10364
rect 20628 10304 20692 10308
rect 20708 10364 20772 10368
rect 20708 10308 20712 10364
rect 20712 10308 20768 10364
rect 20768 10308 20772 10364
rect 20708 10304 20772 10308
rect 20788 10364 20852 10368
rect 20788 10308 20792 10364
rect 20792 10308 20848 10364
rect 20848 10308 20852 10364
rect 20788 10304 20852 10308
rect 27264 10364 27328 10368
rect 27264 10308 27268 10364
rect 27268 10308 27324 10364
rect 27324 10308 27328 10364
rect 27264 10304 27328 10308
rect 27344 10364 27408 10368
rect 27344 10308 27348 10364
rect 27348 10308 27404 10364
rect 27404 10308 27408 10364
rect 27344 10304 27408 10308
rect 27424 10364 27488 10368
rect 27424 10308 27428 10364
rect 27428 10308 27484 10364
rect 27484 10308 27488 10364
rect 27424 10304 27488 10308
rect 27504 10364 27568 10368
rect 27504 10308 27508 10364
rect 27508 10308 27564 10364
rect 27564 10308 27568 10364
rect 27504 10304 27568 10308
rect 3758 9820 3822 9824
rect 3758 9764 3762 9820
rect 3762 9764 3818 9820
rect 3818 9764 3822 9820
rect 3758 9760 3822 9764
rect 3838 9820 3902 9824
rect 3838 9764 3842 9820
rect 3842 9764 3898 9820
rect 3898 9764 3902 9820
rect 3838 9760 3902 9764
rect 3918 9820 3982 9824
rect 3918 9764 3922 9820
rect 3922 9764 3978 9820
rect 3978 9764 3982 9820
rect 3918 9760 3982 9764
rect 3998 9820 4062 9824
rect 3998 9764 4002 9820
rect 4002 9764 4058 9820
rect 4058 9764 4062 9820
rect 3998 9760 4062 9764
rect 10474 9820 10538 9824
rect 10474 9764 10478 9820
rect 10478 9764 10534 9820
rect 10534 9764 10538 9820
rect 10474 9760 10538 9764
rect 10554 9820 10618 9824
rect 10554 9764 10558 9820
rect 10558 9764 10614 9820
rect 10614 9764 10618 9820
rect 10554 9760 10618 9764
rect 10634 9820 10698 9824
rect 10634 9764 10638 9820
rect 10638 9764 10694 9820
rect 10694 9764 10698 9820
rect 10634 9760 10698 9764
rect 10714 9820 10778 9824
rect 10714 9764 10718 9820
rect 10718 9764 10774 9820
rect 10774 9764 10778 9820
rect 10714 9760 10778 9764
rect 17190 9820 17254 9824
rect 17190 9764 17194 9820
rect 17194 9764 17250 9820
rect 17250 9764 17254 9820
rect 17190 9760 17254 9764
rect 17270 9820 17334 9824
rect 17270 9764 17274 9820
rect 17274 9764 17330 9820
rect 17330 9764 17334 9820
rect 17270 9760 17334 9764
rect 17350 9820 17414 9824
rect 17350 9764 17354 9820
rect 17354 9764 17410 9820
rect 17410 9764 17414 9820
rect 17350 9760 17414 9764
rect 17430 9820 17494 9824
rect 17430 9764 17434 9820
rect 17434 9764 17490 9820
rect 17490 9764 17494 9820
rect 17430 9760 17494 9764
rect 23906 9820 23970 9824
rect 23906 9764 23910 9820
rect 23910 9764 23966 9820
rect 23966 9764 23970 9820
rect 23906 9760 23970 9764
rect 23986 9820 24050 9824
rect 23986 9764 23990 9820
rect 23990 9764 24046 9820
rect 24046 9764 24050 9820
rect 23986 9760 24050 9764
rect 24066 9820 24130 9824
rect 24066 9764 24070 9820
rect 24070 9764 24126 9820
rect 24126 9764 24130 9820
rect 24066 9760 24130 9764
rect 24146 9820 24210 9824
rect 24146 9764 24150 9820
rect 24150 9764 24206 9820
rect 24206 9764 24210 9820
rect 24146 9760 24210 9764
rect 10180 9556 10244 9620
rect 18644 9556 18708 9620
rect 20300 9556 20364 9620
rect 26188 9420 26252 9484
rect 7116 9276 7180 9280
rect 7116 9220 7120 9276
rect 7120 9220 7176 9276
rect 7176 9220 7180 9276
rect 7116 9216 7180 9220
rect 7196 9276 7260 9280
rect 7196 9220 7200 9276
rect 7200 9220 7256 9276
rect 7256 9220 7260 9276
rect 7196 9216 7260 9220
rect 7276 9276 7340 9280
rect 7276 9220 7280 9276
rect 7280 9220 7336 9276
rect 7336 9220 7340 9276
rect 7276 9216 7340 9220
rect 7356 9276 7420 9280
rect 7356 9220 7360 9276
rect 7360 9220 7416 9276
rect 7416 9220 7420 9276
rect 7356 9216 7420 9220
rect 13832 9276 13896 9280
rect 13832 9220 13836 9276
rect 13836 9220 13892 9276
rect 13892 9220 13896 9276
rect 13832 9216 13896 9220
rect 13912 9276 13976 9280
rect 13912 9220 13916 9276
rect 13916 9220 13972 9276
rect 13972 9220 13976 9276
rect 13912 9216 13976 9220
rect 13992 9276 14056 9280
rect 13992 9220 13996 9276
rect 13996 9220 14052 9276
rect 14052 9220 14056 9276
rect 13992 9216 14056 9220
rect 14072 9276 14136 9280
rect 14072 9220 14076 9276
rect 14076 9220 14132 9276
rect 14132 9220 14136 9276
rect 14072 9216 14136 9220
rect 20548 9276 20612 9280
rect 20548 9220 20552 9276
rect 20552 9220 20608 9276
rect 20608 9220 20612 9276
rect 20548 9216 20612 9220
rect 20628 9276 20692 9280
rect 20628 9220 20632 9276
rect 20632 9220 20688 9276
rect 20688 9220 20692 9276
rect 20628 9216 20692 9220
rect 20708 9276 20772 9280
rect 20708 9220 20712 9276
rect 20712 9220 20768 9276
rect 20768 9220 20772 9276
rect 20708 9216 20772 9220
rect 20788 9276 20852 9280
rect 20788 9220 20792 9276
rect 20792 9220 20848 9276
rect 20848 9220 20852 9276
rect 20788 9216 20852 9220
rect 27264 9276 27328 9280
rect 27264 9220 27268 9276
rect 27268 9220 27324 9276
rect 27324 9220 27328 9276
rect 27264 9216 27328 9220
rect 27344 9276 27408 9280
rect 27344 9220 27348 9276
rect 27348 9220 27404 9276
rect 27404 9220 27408 9276
rect 27344 9216 27408 9220
rect 27424 9276 27488 9280
rect 27424 9220 27428 9276
rect 27428 9220 27484 9276
rect 27484 9220 27488 9276
rect 27424 9216 27488 9220
rect 27504 9276 27568 9280
rect 27504 9220 27508 9276
rect 27508 9220 27564 9276
rect 27564 9220 27568 9276
rect 27504 9216 27568 9220
rect 3758 8732 3822 8736
rect 3758 8676 3762 8732
rect 3762 8676 3818 8732
rect 3818 8676 3822 8732
rect 3758 8672 3822 8676
rect 3838 8732 3902 8736
rect 3838 8676 3842 8732
rect 3842 8676 3898 8732
rect 3898 8676 3902 8732
rect 3838 8672 3902 8676
rect 3918 8732 3982 8736
rect 3918 8676 3922 8732
rect 3922 8676 3978 8732
rect 3978 8676 3982 8732
rect 3918 8672 3982 8676
rect 3998 8732 4062 8736
rect 3998 8676 4002 8732
rect 4002 8676 4058 8732
rect 4058 8676 4062 8732
rect 3998 8672 4062 8676
rect 10474 8732 10538 8736
rect 10474 8676 10478 8732
rect 10478 8676 10534 8732
rect 10534 8676 10538 8732
rect 10474 8672 10538 8676
rect 10554 8732 10618 8736
rect 10554 8676 10558 8732
rect 10558 8676 10614 8732
rect 10614 8676 10618 8732
rect 10554 8672 10618 8676
rect 10634 8732 10698 8736
rect 10634 8676 10638 8732
rect 10638 8676 10694 8732
rect 10694 8676 10698 8732
rect 10634 8672 10698 8676
rect 10714 8732 10778 8736
rect 10714 8676 10718 8732
rect 10718 8676 10774 8732
rect 10774 8676 10778 8732
rect 10714 8672 10778 8676
rect 17190 8732 17254 8736
rect 17190 8676 17194 8732
rect 17194 8676 17250 8732
rect 17250 8676 17254 8732
rect 17190 8672 17254 8676
rect 17270 8732 17334 8736
rect 17270 8676 17274 8732
rect 17274 8676 17330 8732
rect 17330 8676 17334 8732
rect 17270 8672 17334 8676
rect 17350 8732 17414 8736
rect 17350 8676 17354 8732
rect 17354 8676 17410 8732
rect 17410 8676 17414 8732
rect 17350 8672 17414 8676
rect 17430 8732 17494 8736
rect 17430 8676 17434 8732
rect 17434 8676 17490 8732
rect 17490 8676 17494 8732
rect 17430 8672 17494 8676
rect 23906 8732 23970 8736
rect 23906 8676 23910 8732
rect 23910 8676 23966 8732
rect 23966 8676 23970 8732
rect 23906 8672 23970 8676
rect 23986 8732 24050 8736
rect 23986 8676 23990 8732
rect 23990 8676 24046 8732
rect 24046 8676 24050 8732
rect 23986 8672 24050 8676
rect 24066 8732 24130 8736
rect 24066 8676 24070 8732
rect 24070 8676 24126 8732
rect 24126 8676 24130 8732
rect 24066 8672 24130 8676
rect 24146 8732 24210 8736
rect 24146 8676 24150 8732
rect 24150 8676 24206 8732
rect 24206 8676 24210 8732
rect 24146 8672 24210 8676
rect 17724 8332 17788 8396
rect 7116 8188 7180 8192
rect 7116 8132 7120 8188
rect 7120 8132 7176 8188
rect 7176 8132 7180 8188
rect 7116 8128 7180 8132
rect 7196 8188 7260 8192
rect 7196 8132 7200 8188
rect 7200 8132 7256 8188
rect 7256 8132 7260 8188
rect 7196 8128 7260 8132
rect 7276 8188 7340 8192
rect 7276 8132 7280 8188
rect 7280 8132 7336 8188
rect 7336 8132 7340 8188
rect 7276 8128 7340 8132
rect 7356 8188 7420 8192
rect 7356 8132 7360 8188
rect 7360 8132 7416 8188
rect 7416 8132 7420 8188
rect 7356 8128 7420 8132
rect 13832 8188 13896 8192
rect 13832 8132 13836 8188
rect 13836 8132 13892 8188
rect 13892 8132 13896 8188
rect 13832 8128 13896 8132
rect 13912 8188 13976 8192
rect 13912 8132 13916 8188
rect 13916 8132 13972 8188
rect 13972 8132 13976 8188
rect 13912 8128 13976 8132
rect 13992 8188 14056 8192
rect 13992 8132 13996 8188
rect 13996 8132 14052 8188
rect 14052 8132 14056 8188
rect 13992 8128 14056 8132
rect 14072 8188 14136 8192
rect 14072 8132 14076 8188
rect 14076 8132 14132 8188
rect 14132 8132 14136 8188
rect 14072 8128 14136 8132
rect 20548 8188 20612 8192
rect 20548 8132 20552 8188
rect 20552 8132 20608 8188
rect 20608 8132 20612 8188
rect 20548 8128 20612 8132
rect 20628 8188 20692 8192
rect 20628 8132 20632 8188
rect 20632 8132 20688 8188
rect 20688 8132 20692 8188
rect 20628 8128 20692 8132
rect 20708 8188 20772 8192
rect 20708 8132 20712 8188
rect 20712 8132 20768 8188
rect 20768 8132 20772 8188
rect 20708 8128 20772 8132
rect 20788 8188 20852 8192
rect 20788 8132 20792 8188
rect 20792 8132 20848 8188
rect 20848 8132 20852 8188
rect 20788 8128 20852 8132
rect 27264 8188 27328 8192
rect 27264 8132 27268 8188
rect 27268 8132 27324 8188
rect 27324 8132 27328 8188
rect 27264 8128 27328 8132
rect 27344 8188 27408 8192
rect 27344 8132 27348 8188
rect 27348 8132 27404 8188
rect 27404 8132 27408 8188
rect 27344 8128 27408 8132
rect 27424 8188 27488 8192
rect 27424 8132 27428 8188
rect 27428 8132 27484 8188
rect 27484 8132 27488 8188
rect 27424 8128 27488 8132
rect 27504 8188 27568 8192
rect 27504 8132 27508 8188
rect 27508 8132 27564 8188
rect 27564 8132 27568 8188
rect 27504 8128 27568 8132
rect 3758 7644 3822 7648
rect 3758 7588 3762 7644
rect 3762 7588 3818 7644
rect 3818 7588 3822 7644
rect 3758 7584 3822 7588
rect 3838 7644 3902 7648
rect 3838 7588 3842 7644
rect 3842 7588 3898 7644
rect 3898 7588 3902 7644
rect 3838 7584 3902 7588
rect 3918 7644 3982 7648
rect 3918 7588 3922 7644
rect 3922 7588 3978 7644
rect 3978 7588 3982 7644
rect 3918 7584 3982 7588
rect 3998 7644 4062 7648
rect 3998 7588 4002 7644
rect 4002 7588 4058 7644
rect 4058 7588 4062 7644
rect 3998 7584 4062 7588
rect 10474 7644 10538 7648
rect 10474 7588 10478 7644
rect 10478 7588 10534 7644
rect 10534 7588 10538 7644
rect 10474 7584 10538 7588
rect 10554 7644 10618 7648
rect 10554 7588 10558 7644
rect 10558 7588 10614 7644
rect 10614 7588 10618 7644
rect 10554 7584 10618 7588
rect 10634 7644 10698 7648
rect 10634 7588 10638 7644
rect 10638 7588 10694 7644
rect 10694 7588 10698 7644
rect 10634 7584 10698 7588
rect 10714 7644 10778 7648
rect 10714 7588 10718 7644
rect 10718 7588 10774 7644
rect 10774 7588 10778 7644
rect 10714 7584 10778 7588
rect 17190 7644 17254 7648
rect 17190 7588 17194 7644
rect 17194 7588 17250 7644
rect 17250 7588 17254 7644
rect 17190 7584 17254 7588
rect 17270 7644 17334 7648
rect 17270 7588 17274 7644
rect 17274 7588 17330 7644
rect 17330 7588 17334 7644
rect 17270 7584 17334 7588
rect 17350 7644 17414 7648
rect 17350 7588 17354 7644
rect 17354 7588 17410 7644
rect 17410 7588 17414 7644
rect 17350 7584 17414 7588
rect 17430 7644 17494 7648
rect 17430 7588 17434 7644
rect 17434 7588 17490 7644
rect 17490 7588 17494 7644
rect 17430 7584 17494 7588
rect 23906 7644 23970 7648
rect 23906 7588 23910 7644
rect 23910 7588 23966 7644
rect 23966 7588 23970 7644
rect 23906 7584 23970 7588
rect 23986 7644 24050 7648
rect 23986 7588 23990 7644
rect 23990 7588 24046 7644
rect 24046 7588 24050 7644
rect 23986 7584 24050 7588
rect 24066 7644 24130 7648
rect 24066 7588 24070 7644
rect 24070 7588 24126 7644
rect 24126 7588 24130 7644
rect 24066 7584 24130 7588
rect 24146 7644 24210 7648
rect 24146 7588 24150 7644
rect 24150 7588 24206 7644
rect 24206 7588 24210 7644
rect 24146 7584 24210 7588
rect 7116 7100 7180 7104
rect 7116 7044 7120 7100
rect 7120 7044 7176 7100
rect 7176 7044 7180 7100
rect 7116 7040 7180 7044
rect 7196 7100 7260 7104
rect 7196 7044 7200 7100
rect 7200 7044 7256 7100
rect 7256 7044 7260 7100
rect 7196 7040 7260 7044
rect 7276 7100 7340 7104
rect 7276 7044 7280 7100
rect 7280 7044 7336 7100
rect 7336 7044 7340 7100
rect 7276 7040 7340 7044
rect 7356 7100 7420 7104
rect 7356 7044 7360 7100
rect 7360 7044 7416 7100
rect 7416 7044 7420 7100
rect 7356 7040 7420 7044
rect 13832 7100 13896 7104
rect 13832 7044 13836 7100
rect 13836 7044 13892 7100
rect 13892 7044 13896 7100
rect 13832 7040 13896 7044
rect 13912 7100 13976 7104
rect 13912 7044 13916 7100
rect 13916 7044 13972 7100
rect 13972 7044 13976 7100
rect 13912 7040 13976 7044
rect 13992 7100 14056 7104
rect 13992 7044 13996 7100
rect 13996 7044 14052 7100
rect 14052 7044 14056 7100
rect 13992 7040 14056 7044
rect 14072 7100 14136 7104
rect 14072 7044 14076 7100
rect 14076 7044 14132 7100
rect 14132 7044 14136 7100
rect 14072 7040 14136 7044
rect 20548 7100 20612 7104
rect 20548 7044 20552 7100
rect 20552 7044 20608 7100
rect 20608 7044 20612 7100
rect 20548 7040 20612 7044
rect 20628 7100 20692 7104
rect 20628 7044 20632 7100
rect 20632 7044 20688 7100
rect 20688 7044 20692 7100
rect 20628 7040 20692 7044
rect 20708 7100 20772 7104
rect 20708 7044 20712 7100
rect 20712 7044 20768 7100
rect 20768 7044 20772 7100
rect 20708 7040 20772 7044
rect 20788 7100 20852 7104
rect 20788 7044 20792 7100
rect 20792 7044 20848 7100
rect 20848 7044 20852 7100
rect 20788 7040 20852 7044
rect 27264 7100 27328 7104
rect 27264 7044 27268 7100
rect 27268 7044 27324 7100
rect 27324 7044 27328 7100
rect 27264 7040 27328 7044
rect 27344 7100 27408 7104
rect 27344 7044 27348 7100
rect 27348 7044 27404 7100
rect 27404 7044 27408 7100
rect 27344 7040 27408 7044
rect 27424 7100 27488 7104
rect 27424 7044 27428 7100
rect 27428 7044 27484 7100
rect 27484 7044 27488 7100
rect 27424 7040 27488 7044
rect 27504 7100 27568 7104
rect 27504 7044 27508 7100
rect 27508 7044 27564 7100
rect 27564 7044 27568 7100
rect 27504 7040 27568 7044
rect 3758 6556 3822 6560
rect 3758 6500 3762 6556
rect 3762 6500 3818 6556
rect 3818 6500 3822 6556
rect 3758 6496 3822 6500
rect 3838 6556 3902 6560
rect 3838 6500 3842 6556
rect 3842 6500 3898 6556
rect 3898 6500 3902 6556
rect 3838 6496 3902 6500
rect 3918 6556 3982 6560
rect 3918 6500 3922 6556
rect 3922 6500 3978 6556
rect 3978 6500 3982 6556
rect 3918 6496 3982 6500
rect 3998 6556 4062 6560
rect 3998 6500 4002 6556
rect 4002 6500 4058 6556
rect 4058 6500 4062 6556
rect 3998 6496 4062 6500
rect 10474 6556 10538 6560
rect 10474 6500 10478 6556
rect 10478 6500 10534 6556
rect 10534 6500 10538 6556
rect 10474 6496 10538 6500
rect 10554 6556 10618 6560
rect 10554 6500 10558 6556
rect 10558 6500 10614 6556
rect 10614 6500 10618 6556
rect 10554 6496 10618 6500
rect 10634 6556 10698 6560
rect 10634 6500 10638 6556
rect 10638 6500 10694 6556
rect 10694 6500 10698 6556
rect 10634 6496 10698 6500
rect 10714 6556 10778 6560
rect 10714 6500 10718 6556
rect 10718 6500 10774 6556
rect 10774 6500 10778 6556
rect 10714 6496 10778 6500
rect 17190 6556 17254 6560
rect 17190 6500 17194 6556
rect 17194 6500 17250 6556
rect 17250 6500 17254 6556
rect 17190 6496 17254 6500
rect 17270 6556 17334 6560
rect 17270 6500 17274 6556
rect 17274 6500 17330 6556
rect 17330 6500 17334 6556
rect 17270 6496 17334 6500
rect 17350 6556 17414 6560
rect 17350 6500 17354 6556
rect 17354 6500 17410 6556
rect 17410 6500 17414 6556
rect 17350 6496 17414 6500
rect 17430 6556 17494 6560
rect 17430 6500 17434 6556
rect 17434 6500 17490 6556
rect 17490 6500 17494 6556
rect 17430 6496 17494 6500
rect 23906 6556 23970 6560
rect 23906 6500 23910 6556
rect 23910 6500 23966 6556
rect 23966 6500 23970 6556
rect 23906 6496 23970 6500
rect 23986 6556 24050 6560
rect 23986 6500 23990 6556
rect 23990 6500 24046 6556
rect 24046 6500 24050 6556
rect 23986 6496 24050 6500
rect 24066 6556 24130 6560
rect 24066 6500 24070 6556
rect 24070 6500 24126 6556
rect 24126 6500 24130 6556
rect 24066 6496 24130 6500
rect 24146 6556 24210 6560
rect 24146 6500 24150 6556
rect 24150 6500 24206 6556
rect 24206 6500 24210 6556
rect 24146 6496 24210 6500
rect 10180 6292 10244 6356
rect 7116 6012 7180 6016
rect 7116 5956 7120 6012
rect 7120 5956 7176 6012
rect 7176 5956 7180 6012
rect 7116 5952 7180 5956
rect 7196 6012 7260 6016
rect 7196 5956 7200 6012
rect 7200 5956 7256 6012
rect 7256 5956 7260 6012
rect 7196 5952 7260 5956
rect 7276 6012 7340 6016
rect 7276 5956 7280 6012
rect 7280 5956 7336 6012
rect 7336 5956 7340 6012
rect 7276 5952 7340 5956
rect 7356 6012 7420 6016
rect 7356 5956 7360 6012
rect 7360 5956 7416 6012
rect 7416 5956 7420 6012
rect 7356 5952 7420 5956
rect 13832 6012 13896 6016
rect 13832 5956 13836 6012
rect 13836 5956 13892 6012
rect 13892 5956 13896 6012
rect 13832 5952 13896 5956
rect 13912 6012 13976 6016
rect 13912 5956 13916 6012
rect 13916 5956 13972 6012
rect 13972 5956 13976 6012
rect 13912 5952 13976 5956
rect 13992 6012 14056 6016
rect 13992 5956 13996 6012
rect 13996 5956 14052 6012
rect 14052 5956 14056 6012
rect 13992 5952 14056 5956
rect 14072 6012 14136 6016
rect 14072 5956 14076 6012
rect 14076 5956 14132 6012
rect 14132 5956 14136 6012
rect 14072 5952 14136 5956
rect 20548 6012 20612 6016
rect 20548 5956 20552 6012
rect 20552 5956 20608 6012
rect 20608 5956 20612 6012
rect 20548 5952 20612 5956
rect 20628 6012 20692 6016
rect 20628 5956 20632 6012
rect 20632 5956 20688 6012
rect 20688 5956 20692 6012
rect 20628 5952 20692 5956
rect 20708 6012 20772 6016
rect 20708 5956 20712 6012
rect 20712 5956 20768 6012
rect 20768 5956 20772 6012
rect 20708 5952 20772 5956
rect 20788 6012 20852 6016
rect 20788 5956 20792 6012
rect 20792 5956 20848 6012
rect 20848 5956 20852 6012
rect 20788 5952 20852 5956
rect 27264 6012 27328 6016
rect 27264 5956 27268 6012
rect 27268 5956 27324 6012
rect 27324 5956 27328 6012
rect 27264 5952 27328 5956
rect 27344 6012 27408 6016
rect 27344 5956 27348 6012
rect 27348 5956 27404 6012
rect 27404 5956 27408 6012
rect 27344 5952 27408 5956
rect 27424 6012 27488 6016
rect 27424 5956 27428 6012
rect 27428 5956 27484 6012
rect 27484 5956 27488 6012
rect 27424 5952 27488 5956
rect 27504 6012 27568 6016
rect 27504 5956 27508 6012
rect 27508 5956 27564 6012
rect 27564 5956 27568 6012
rect 27504 5952 27568 5956
rect 3758 5468 3822 5472
rect 3758 5412 3762 5468
rect 3762 5412 3818 5468
rect 3818 5412 3822 5468
rect 3758 5408 3822 5412
rect 3838 5468 3902 5472
rect 3838 5412 3842 5468
rect 3842 5412 3898 5468
rect 3898 5412 3902 5468
rect 3838 5408 3902 5412
rect 3918 5468 3982 5472
rect 3918 5412 3922 5468
rect 3922 5412 3978 5468
rect 3978 5412 3982 5468
rect 3918 5408 3982 5412
rect 3998 5468 4062 5472
rect 3998 5412 4002 5468
rect 4002 5412 4058 5468
rect 4058 5412 4062 5468
rect 3998 5408 4062 5412
rect 10474 5468 10538 5472
rect 10474 5412 10478 5468
rect 10478 5412 10534 5468
rect 10534 5412 10538 5468
rect 10474 5408 10538 5412
rect 10554 5468 10618 5472
rect 10554 5412 10558 5468
rect 10558 5412 10614 5468
rect 10614 5412 10618 5468
rect 10554 5408 10618 5412
rect 10634 5468 10698 5472
rect 10634 5412 10638 5468
rect 10638 5412 10694 5468
rect 10694 5412 10698 5468
rect 10634 5408 10698 5412
rect 10714 5468 10778 5472
rect 10714 5412 10718 5468
rect 10718 5412 10774 5468
rect 10774 5412 10778 5468
rect 10714 5408 10778 5412
rect 17190 5468 17254 5472
rect 17190 5412 17194 5468
rect 17194 5412 17250 5468
rect 17250 5412 17254 5468
rect 17190 5408 17254 5412
rect 17270 5468 17334 5472
rect 17270 5412 17274 5468
rect 17274 5412 17330 5468
rect 17330 5412 17334 5468
rect 17270 5408 17334 5412
rect 17350 5468 17414 5472
rect 17350 5412 17354 5468
rect 17354 5412 17410 5468
rect 17410 5412 17414 5468
rect 17350 5408 17414 5412
rect 17430 5468 17494 5472
rect 17430 5412 17434 5468
rect 17434 5412 17490 5468
rect 17490 5412 17494 5468
rect 17430 5408 17494 5412
rect 23906 5468 23970 5472
rect 23906 5412 23910 5468
rect 23910 5412 23966 5468
rect 23966 5412 23970 5468
rect 23906 5408 23970 5412
rect 23986 5468 24050 5472
rect 23986 5412 23990 5468
rect 23990 5412 24046 5468
rect 24046 5412 24050 5468
rect 23986 5408 24050 5412
rect 24066 5468 24130 5472
rect 24066 5412 24070 5468
rect 24070 5412 24126 5468
rect 24126 5412 24130 5468
rect 24066 5408 24130 5412
rect 24146 5468 24210 5472
rect 24146 5412 24150 5468
rect 24150 5412 24206 5468
rect 24206 5412 24210 5468
rect 24146 5408 24210 5412
rect 20300 5204 20364 5268
rect 7116 4924 7180 4928
rect 7116 4868 7120 4924
rect 7120 4868 7176 4924
rect 7176 4868 7180 4924
rect 7116 4864 7180 4868
rect 7196 4924 7260 4928
rect 7196 4868 7200 4924
rect 7200 4868 7256 4924
rect 7256 4868 7260 4924
rect 7196 4864 7260 4868
rect 7276 4924 7340 4928
rect 7276 4868 7280 4924
rect 7280 4868 7336 4924
rect 7336 4868 7340 4924
rect 7276 4864 7340 4868
rect 7356 4924 7420 4928
rect 7356 4868 7360 4924
rect 7360 4868 7416 4924
rect 7416 4868 7420 4924
rect 7356 4864 7420 4868
rect 13832 4924 13896 4928
rect 13832 4868 13836 4924
rect 13836 4868 13892 4924
rect 13892 4868 13896 4924
rect 13832 4864 13896 4868
rect 13912 4924 13976 4928
rect 13912 4868 13916 4924
rect 13916 4868 13972 4924
rect 13972 4868 13976 4924
rect 13912 4864 13976 4868
rect 13992 4924 14056 4928
rect 13992 4868 13996 4924
rect 13996 4868 14052 4924
rect 14052 4868 14056 4924
rect 13992 4864 14056 4868
rect 14072 4924 14136 4928
rect 14072 4868 14076 4924
rect 14076 4868 14132 4924
rect 14132 4868 14136 4924
rect 14072 4864 14136 4868
rect 20548 4924 20612 4928
rect 20548 4868 20552 4924
rect 20552 4868 20608 4924
rect 20608 4868 20612 4924
rect 20548 4864 20612 4868
rect 20628 4924 20692 4928
rect 20628 4868 20632 4924
rect 20632 4868 20688 4924
rect 20688 4868 20692 4924
rect 20628 4864 20692 4868
rect 20708 4924 20772 4928
rect 20708 4868 20712 4924
rect 20712 4868 20768 4924
rect 20768 4868 20772 4924
rect 20708 4864 20772 4868
rect 20788 4924 20852 4928
rect 20788 4868 20792 4924
rect 20792 4868 20848 4924
rect 20848 4868 20852 4924
rect 20788 4864 20852 4868
rect 27264 4924 27328 4928
rect 27264 4868 27268 4924
rect 27268 4868 27324 4924
rect 27324 4868 27328 4924
rect 27264 4864 27328 4868
rect 27344 4924 27408 4928
rect 27344 4868 27348 4924
rect 27348 4868 27404 4924
rect 27404 4868 27408 4924
rect 27344 4864 27408 4868
rect 27424 4924 27488 4928
rect 27424 4868 27428 4924
rect 27428 4868 27484 4924
rect 27484 4868 27488 4924
rect 27424 4864 27488 4868
rect 27504 4924 27568 4928
rect 27504 4868 27508 4924
rect 27508 4868 27564 4924
rect 27564 4868 27568 4924
rect 27504 4864 27568 4868
rect 3758 4380 3822 4384
rect 3758 4324 3762 4380
rect 3762 4324 3818 4380
rect 3818 4324 3822 4380
rect 3758 4320 3822 4324
rect 3838 4380 3902 4384
rect 3838 4324 3842 4380
rect 3842 4324 3898 4380
rect 3898 4324 3902 4380
rect 3838 4320 3902 4324
rect 3918 4380 3982 4384
rect 3918 4324 3922 4380
rect 3922 4324 3978 4380
rect 3978 4324 3982 4380
rect 3918 4320 3982 4324
rect 3998 4380 4062 4384
rect 3998 4324 4002 4380
rect 4002 4324 4058 4380
rect 4058 4324 4062 4380
rect 3998 4320 4062 4324
rect 10474 4380 10538 4384
rect 10474 4324 10478 4380
rect 10478 4324 10534 4380
rect 10534 4324 10538 4380
rect 10474 4320 10538 4324
rect 10554 4380 10618 4384
rect 10554 4324 10558 4380
rect 10558 4324 10614 4380
rect 10614 4324 10618 4380
rect 10554 4320 10618 4324
rect 10634 4380 10698 4384
rect 10634 4324 10638 4380
rect 10638 4324 10694 4380
rect 10694 4324 10698 4380
rect 10634 4320 10698 4324
rect 10714 4380 10778 4384
rect 10714 4324 10718 4380
rect 10718 4324 10774 4380
rect 10774 4324 10778 4380
rect 10714 4320 10778 4324
rect 17190 4380 17254 4384
rect 17190 4324 17194 4380
rect 17194 4324 17250 4380
rect 17250 4324 17254 4380
rect 17190 4320 17254 4324
rect 17270 4380 17334 4384
rect 17270 4324 17274 4380
rect 17274 4324 17330 4380
rect 17330 4324 17334 4380
rect 17270 4320 17334 4324
rect 17350 4380 17414 4384
rect 17350 4324 17354 4380
rect 17354 4324 17410 4380
rect 17410 4324 17414 4380
rect 17350 4320 17414 4324
rect 17430 4380 17494 4384
rect 17430 4324 17434 4380
rect 17434 4324 17490 4380
rect 17490 4324 17494 4380
rect 17430 4320 17494 4324
rect 23906 4380 23970 4384
rect 23906 4324 23910 4380
rect 23910 4324 23966 4380
rect 23966 4324 23970 4380
rect 23906 4320 23970 4324
rect 23986 4380 24050 4384
rect 23986 4324 23990 4380
rect 23990 4324 24046 4380
rect 24046 4324 24050 4380
rect 23986 4320 24050 4324
rect 24066 4380 24130 4384
rect 24066 4324 24070 4380
rect 24070 4324 24126 4380
rect 24126 4324 24130 4380
rect 24066 4320 24130 4324
rect 24146 4380 24210 4384
rect 24146 4324 24150 4380
rect 24150 4324 24206 4380
rect 24206 4324 24210 4380
rect 24146 4320 24210 4324
rect 18276 4040 18340 4044
rect 18276 3984 18326 4040
rect 18326 3984 18340 4040
rect 18276 3980 18340 3984
rect 22324 3980 22388 4044
rect 7116 3836 7180 3840
rect 7116 3780 7120 3836
rect 7120 3780 7176 3836
rect 7176 3780 7180 3836
rect 7116 3776 7180 3780
rect 7196 3836 7260 3840
rect 7196 3780 7200 3836
rect 7200 3780 7256 3836
rect 7256 3780 7260 3836
rect 7196 3776 7260 3780
rect 7276 3836 7340 3840
rect 7276 3780 7280 3836
rect 7280 3780 7336 3836
rect 7336 3780 7340 3836
rect 7276 3776 7340 3780
rect 7356 3836 7420 3840
rect 7356 3780 7360 3836
rect 7360 3780 7416 3836
rect 7416 3780 7420 3836
rect 7356 3776 7420 3780
rect 13832 3836 13896 3840
rect 13832 3780 13836 3836
rect 13836 3780 13892 3836
rect 13892 3780 13896 3836
rect 13832 3776 13896 3780
rect 13912 3836 13976 3840
rect 13912 3780 13916 3836
rect 13916 3780 13972 3836
rect 13972 3780 13976 3836
rect 13912 3776 13976 3780
rect 13992 3836 14056 3840
rect 13992 3780 13996 3836
rect 13996 3780 14052 3836
rect 14052 3780 14056 3836
rect 13992 3776 14056 3780
rect 14072 3836 14136 3840
rect 14072 3780 14076 3836
rect 14076 3780 14132 3836
rect 14132 3780 14136 3836
rect 14072 3776 14136 3780
rect 20548 3836 20612 3840
rect 20548 3780 20552 3836
rect 20552 3780 20608 3836
rect 20608 3780 20612 3836
rect 20548 3776 20612 3780
rect 20628 3836 20692 3840
rect 20628 3780 20632 3836
rect 20632 3780 20688 3836
rect 20688 3780 20692 3836
rect 20628 3776 20692 3780
rect 20708 3836 20772 3840
rect 20708 3780 20712 3836
rect 20712 3780 20768 3836
rect 20768 3780 20772 3836
rect 20708 3776 20772 3780
rect 20788 3836 20852 3840
rect 20788 3780 20792 3836
rect 20792 3780 20848 3836
rect 20848 3780 20852 3836
rect 20788 3776 20852 3780
rect 27264 3836 27328 3840
rect 27264 3780 27268 3836
rect 27268 3780 27324 3836
rect 27324 3780 27328 3836
rect 27264 3776 27328 3780
rect 27344 3836 27408 3840
rect 27344 3780 27348 3836
rect 27348 3780 27404 3836
rect 27404 3780 27408 3836
rect 27344 3776 27408 3780
rect 27424 3836 27488 3840
rect 27424 3780 27428 3836
rect 27428 3780 27484 3836
rect 27484 3780 27488 3836
rect 27424 3776 27488 3780
rect 27504 3836 27568 3840
rect 27504 3780 27508 3836
rect 27508 3780 27564 3836
rect 27564 3780 27568 3836
rect 27504 3776 27568 3780
rect 3758 3292 3822 3296
rect 3758 3236 3762 3292
rect 3762 3236 3818 3292
rect 3818 3236 3822 3292
rect 3758 3232 3822 3236
rect 3838 3292 3902 3296
rect 3838 3236 3842 3292
rect 3842 3236 3898 3292
rect 3898 3236 3902 3292
rect 3838 3232 3902 3236
rect 3918 3292 3982 3296
rect 3918 3236 3922 3292
rect 3922 3236 3978 3292
rect 3978 3236 3982 3292
rect 3918 3232 3982 3236
rect 3998 3292 4062 3296
rect 3998 3236 4002 3292
rect 4002 3236 4058 3292
rect 4058 3236 4062 3292
rect 3998 3232 4062 3236
rect 10474 3292 10538 3296
rect 10474 3236 10478 3292
rect 10478 3236 10534 3292
rect 10534 3236 10538 3292
rect 10474 3232 10538 3236
rect 10554 3292 10618 3296
rect 10554 3236 10558 3292
rect 10558 3236 10614 3292
rect 10614 3236 10618 3292
rect 10554 3232 10618 3236
rect 10634 3292 10698 3296
rect 10634 3236 10638 3292
rect 10638 3236 10694 3292
rect 10694 3236 10698 3292
rect 10634 3232 10698 3236
rect 10714 3292 10778 3296
rect 10714 3236 10718 3292
rect 10718 3236 10774 3292
rect 10774 3236 10778 3292
rect 10714 3232 10778 3236
rect 17190 3292 17254 3296
rect 17190 3236 17194 3292
rect 17194 3236 17250 3292
rect 17250 3236 17254 3292
rect 17190 3232 17254 3236
rect 17270 3292 17334 3296
rect 17270 3236 17274 3292
rect 17274 3236 17330 3292
rect 17330 3236 17334 3292
rect 17270 3232 17334 3236
rect 17350 3292 17414 3296
rect 17350 3236 17354 3292
rect 17354 3236 17410 3292
rect 17410 3236 17414 3292
rect 17350 3232 17414 3236
rect 17430 3292 17494 3296
rect 17430 3236 17434 3292
rect 17434 3236 17490 3292
rect 17490 3236 17494 3292
rect 17430 3232 17494 3236
rect 23906 3292 23970 3296
rect 23906 3236 23910 3292
rect 23910 3236 23966 3292
rect 23966 3236 23970 3292
rect 23906 3232 23970 3236
rect 23986 3292 24050 3296
rect 23986 3236 23990 3292
rect 23990 3236 24046 3292
rect 24046 3236 24050 3292
rect 23986 3232 24050 3236
rect 24066 3292 24130 3296
rect 24066 3236 24070 3292
rect 24070 3236 24126 3292
rect 24126 3236 24130 3292
rect 24066 3232 24130 3236
rect 24146 3292 24210 3296
rect 24146 3236 24150 3292
rect 24150 3236 24206 3292
rect 24206 3236 24210 3292
rect 24146 3232 24210 3236
rect 7116 2748 7180 2752
rect 7116 2692 7120 2748
rect 7120 2692 7176 2748
rect 7176 2692 7180 2748
rect 7116 2688 7180 2692
rect 7196 2748 7260 2752
rect 7196 2692 7200 2748
rect 7200 2692 7256 2748
rect 7256 2692 7260 2748
rect 7196 2688 7260 2692
rect 7276 2748 7340 2752
rect 7276 2692 7280 2748
rect 7280 2692 7336 2748
rect 7336 2692 7340 2748
rect 7276 2688 7340 2692
rect 7356 2748 7420 2752
rect 7356 2692 7360 2748
rect 7360 2692 7416 2748
rect 7416 2692 7420 2748
rect 7356 2688 7420 2692
rect 13832 2748 13896 2752
rect 13832 2692 13836 2748
rect 13836 2692 13892 2748
rect 13892 2692 13896 2748
rect 13832 2688 13896 2692
rect 13912 2748 13976 2752
rect 13912 2692 13916 2748
rect 13916 2692 13972 2748
rect 13972 2692 13976 2748
rect 13912 2688 13976 2692
rect 13992 2748 14056 2752
rect 13992 2692 13996 2748
rect 13996 2692 14052 2748
rect 14052 2692 14056 2748
rect 13992 2688 14056 2692
rect 14072 2748 14136 2752
rect 14072 2692 14076 2748
rect 14076 2692 14132 2748
rect 14132 2692 14136 2748
rect 14072 2688 14136 2692
rect 20548 2748 20612 2752
rect 20548 2692 20552 2748
rect 20552 2692 20608 2748
rect 20608 2692 20612 2748
rect 20548 2688 20612 2692
rect 20628 2748 20692 2752
rect 20628 2692 20632 2748
rect 20632 2692 20688 2748
rect 20688 2692 20692 2748
rect 20628 2688 20692 2692
rect 20708 2748 20772 2752
rect 20708 2692 20712 2748
rect 20712 2692 20768 2748
rect 20768 2692 20772 2748
rect 20708 2688 20772 2692
rect 20788 2748 20852 2752
rect 20788 2692 20792 2748
rect 20792 2692 20848 2748
rect 20848 2692 20852 2748
rect 20788 2688 20852 2692
rect 27264 2748 27328 2752
rect 27264 2692 27268 2748
rect 27268 2692 27324 2748
rect 27324 2692 27328 2748
rect 27264 2688 27328 2692
rect 27344 2748 27408 2752
rect 27344 2692 27348 2748
rect 27348 2692 27404 2748
rect 27404 2692 27408 2748
rect 27344 2688 27408 2692
rect 27424 2748 27488 2752
rect 27424 2692 27428 2748
rect 27428 2692 27484 2748
rect 27484 2692 27488 2748
rect 27424 2688 27488 2692
rect 27504 2748 27568 2752
rect 27504 2692 27508 2748
rect 27508 2692 27564 2748
rect 27564 2692 27568 2748
rect 27504 2688 27568 2692
rect 3758 2204 3822 2208
rect 3758 2148 3762 2204
rect 3762 2148 3818 2204
rect 3818 2148 3822 2204
rect 3758 2144 3822 2148
rect 3838 2204 3902 2208
rect 3838 2148 3842 2204
rect 3842 2148 3898 2204
rect 3898 2148 3902 2204
rect 3838 2144 3902 2148
rect 3918 2204 3982 2208
rect 3918 2148 3922 2204
rect 3922 2148 3978 2204
rect 3978 2148 3982 2204
rect 3918 2144 3982 2148
rect 3998 2204 4062 2208
rect 3998 2148 4002 2204
rect 4002 2148 4058 2204
rect 4058 2148 4062 2204
rect 3998 2144 4062 2148
rect 10474 2204 10538 2208
rect 10474 2148 10478 2204
rect 10478 2148 10534 2204
rect 10534 2148 10538 2204
rect 10474 2144 10538 2148
rect 10554 2204 10618 2208
rect 10554 2148 10558 2204
rect 10558 2148 10614 2204
rect 10614 2148 10618 2204
rect 10554 2144 10618 2148
rect 10634 2204 10698 2208
rect 10634 2148 10638 2204
rect 10638 2148 10694 2204
rect 10694 2148 10698 2204
rect 10634 2144 10698 2148
rect 10714 2204 10778 2208
rect 10714 2148 10718 2204
rect 10718 2148 10774 2204
rect 10774 2148 10778 2204
rect 10714 2144 10778 2148
rect 17190 2204 17254 2208
rect 17190 2148 17194 2204
rect 17194 2148 17250 2204
rect 17250 2148 17254 2204
rect 17190 2144 17254 2148
rect 17270 2204 17334 2208
rect 17270 2148 17274 2204
rect 17274 2148 17330 2204
rect 17330 2148 17334 2204
rect 17270 2144 17334 2148
rect 17350 2204 17414 2208
rect 17350 2148 17354 2204
rect 17354 2148 17410 2204
rect 17410 2148 17414 2204
rect 17350 2144 17414 2148
rect 17430 2204 17494 2208
rect 17430 2148 17434 2204
rect 17434 2148 17490 2204
rect 17490 2148 17494 2204
rect 17430 2144 17494 2148
rect 23906 2204 23970 2208
rect 23906 2148 23910 2204
rect 23910 2148 23966 2204
rect 23966 2148 23970 2204
rect 23906 2144 23970 2148
rect 23986 2204 24050 2208
rect 23986 2148 23990 2204
rect 23990 2148 24046 2204
rect 24046 2148 24050 2204
rect 23986 2144 24050 2148
rect 24066 2204 24130 2208
rect 24066 2148 24070 2204
rect 24070 2148 24126 2204
rect 24126 2148 24130 2204
rect 24066 2144 24130 2148
rect 24146 2204 24210 2208
rect 24146 2148 24150 2204
rect 24150 2148 24206 2204
rect 24206 2148 24210 2204
rect 24146 2144 24210 2148
rect 7116 1660 7180 1664
rect 7116 1604 7120 1660
rect 7120 1604 7176 1660
rect 7176 1604 7180 1660
rect 7116 1600 7180 1604
rect 7196 1660 7260 1664
rect 7196 1604 7200 1660
rect 7200 1604 7256 1660
rect 7256 1604 7260 1660
rect 7196 1600 7260 1604
rect 7276 1660 7340 1664
rect 7276 1604 7280 1660
rect 7280 1604 7336 1660
rect 7336 1604 7340 1660
rect 7276 1600 7340 1604
rect 7356 1660 7420 1664
rect 7356 1604 7360 1660
rect 7360 1604 7416 1660
rect 7416 1604 7420 1660
rect 7356 1600 7420 1604
rect 13832 1660 13896 1664
rect 13832 1604 13836 1660
rect 13836 1604 13892 1660
rect 13892 1604 13896 1660
rect 13832 1600 13896 1604
rect 13912 1660 13976 1664
rect 13912 1604 13916 1660
rect 13916 1604 13972 1660
rect 13972 1604 13976 1660
rect 13912 1600 13976 1604
rect 13992 1660 14056 1664
rect 13992 1604 13996 1660
rect 13996 1604 14052 1660
rect 14052 1604 14056 1660
rect 13992 1600 14056 1604
rect 14072 1660 14136 1664
rect 14072 1604 14076 1660
rect 14076 1604 14132 1660
rect 14132 1604 14136 1660
rect 14072 1600 14136 1604
rect 20548 1660 20612 1664
rect 20548 1604 20552 1660
rect 20552 1604 20608 1660
rect 20608 1604 20612 1660
rect 20548 1600 20612 1604
rect 20628 1660 20692 1664
rect 20628 1604 20632 1660
rect 20632 1604 20688 1660
rect 20688 1604 20692 1660
rect 20628 1600 20692 1604
rect 20708 1660 20772 1664
rect 20708 1604 20712 1660
rect 20712 1604 20768 1660
rect 20768 1604 20772 1660
rect 20708 1600 20772 1604
rect 20788 1660 20852 1664
rect 20788 1604 20792 1660
rect 20792 1604 20848 1660
rect 20848 1604 20852 1660
rect 20788 1600 20852 1604
rect 27264 1660 27328 1664
rect 27264 1604 27268 1660
rect 27268 1604 27324 1660
rect 27324 1604 27328 1660
rect 27264 1600 27328 1604
rect 27344 1660 27408 1664
rect 27344 1604 27348 1660
rect 27348 1604 27404 1660
rect 27404 1604 27408 1660
rect 27344 1600 27408 1604
rect 27424 1660 27488 1664
rect 27424 1604 27428 1660
rect 27428 1604 27484 1660
rect 27484 1604 27488 1660
rect 27424 1600 27488 1604
rect 27504 1660 27568 1664
rect 27504 1604 27508 1660
rect 27508 1604 27564 1660
rect 27564 1604 27568 1660
rect 27504 1600 27568 1604
rect 3758 1116 3822 1120
rect 3758 1060 3762 1116
rect 3762 1060 3818 1116
rect 3818 1060 3822 1116
rect 3758 1056 3822 1060
rect 3838 1116 3902 1120
rect 3838 1060 3842 1116
rect 3842 1060 3898 1116
rect 3898 1060 3902 1116
rect 3838 1056 3902 1060
rect 3918 1116 3982 1120
rect 3918 1060 3922 1116
rect 3922 1060 3978 1116
rect 3978 1060 3982 1116
rect 3918 1056 3982 1060
rect 3998 1116 4062 1120
rect 3998 1060 4002 1116
rect 4002 1060 4058 1116
rect 4058 1060 4062 1116
rect 3998 1056 4062 1060
rect 10474 1116 10538 1120
rect 10474 1060 10478 1116
rect 10478 1060 10534 1116
rect 10534 1060 10538 1116
rect 10474 1056 10538 1060
rect 10554 1116 10618 1120
rect 10554 1060 10558 1116
rect 10558 1060 10614 1116
rect 10614 1060 10618 1116
rect 10554 1056 10618 1060
rect 10634 1116 10698 1120
rect 10634 1060 10638 1116
rect 10638 1060 10694 1116
rect 10694 1060 10698 1116
rect 10634 1056 10698 1060
rect 10714 1116 10778 1120
rect 10714 1060 10718 1116
rect 10718 1060 10774 1116
rect 10774 1060 10778 1116
rect 10714 1056 10778 1060
rect 17190 1116 17254 1120
rect 17190 1060 17194 1116
rect 17194 1060 17250 1116
rect 17250 1060 17254 1116
rect 17190 1056 17254 1060
rect 17270 1116 17334 1120
rect 17270 1060 17274 1116
rect 17274 1060 17330 1116
rect 17330 1060 17334 1116
rect 17270 1056 17334 1060
rect 17350 1116 17414 1120
rect 17350 1060 17354 1116
rect 17354 1060 17410 1116
rect 17410 1060 17414 1116
rect 17350 1056 17414 1060
rect 17430 1116 17494 1120
rect 17430 1060 17434 1116
rect 17434 1060 17490 1116
rect 17490 1060 17494 1116
rect 17430 1056 17494 1060
rect 23906 1116 23970 1120
rect 23906 1060 23910 1116
rect 23910 1060 23966 1116
rect 23966 1060 23970 1116
rect 23906 1056 23970 1060
rect 23986 1116 24050 1120
rect 23986 1060 23990 1116
rect 23990 1060 24046 1116
rect 24046 1060 24050 1116
rect 23986 1056 24050 1060
rect 24066 1116 24130 1120
rect 24066 1060 24070 1116
rect 24070 1060 24126 1116
rect 24126 1060 24130 1116
rect 24066 1056 24130 1060
rect 24146 1116 24210 1120
rect 24146 1060 24150 1116
rect 24150 1060 24206 1116
rect 24206 1060 24210 1116
rect 24146 1056 24210 1060
rect 7116 572 7180 576
rect 7116 516 7120 572
rect 7120 516 7176 572
rect 7176 516 7180 572
rect 7116 512 7180 516
rect 7196 572 7260 576
rect 7196 516 7200 572
rect 7200 516 7256 572
rect 7256 516 7260 572
rect 7196 512 7260 516
rect 7276 572 7340 576
rect 7276 516 7280 572
rect 7280 516 7336 572
rect 7336 516 7340 572
rect 7276 512 7340 516
rect 7356 572 7420 576
rect 7356 516 7360 572
rect 7360 516 7416 572
rect 7416 516 7420 572
rect 7356 512 7420 516
rect 13832 572 13896 576
rect 13832 516 13836 572
rect 13836 516 13892 572
rect 13892 516 13896 572
rect 13832 512 13896 516
rect 13912 572 13976 576
rect 13912 516 13916 572
rect 13916 516 13972 572
rect 13972 516 13976 572
rect 13912 512 13976 516
rect 13992 572 14056 576
rect 13992 516 13996 572
rect 13996 516 14052 572
rect 14052 516 14056 572
rect 13992 512 14056 516
rect 14072 572 14136 576
rect 14072 516 14076 572
rect 14076 516 14132 572
rect 14132 516 14136 572
rect 14072 512 14136 516
rect 20548 572 20612 576
rect 20548 516 20552 572
rect 20552 516 20608 572
rect 20608 516 20612 572
rect 20548 512 20612 516
rect 20628 572 20692 576
rect 20628 516 20632 572
rect 20632 516 20688 572
rect 20688 516 20692 572
rect 20628 512 20692 516
rect 20708 572 20772 576
rect 20708 516 20712 572
rect 20712 516 20768 572
rect 20768 516 20772 572
rect 20708 512 20772 516
rect 20788 572 20852 576
rect 20788 516 20792 572
rect 20792 516 20848 572
rect 20848 516 20852 572
rect 20788 512 20852 516
rect 27264 572 27328 576
rect 27264 516 27268 572
rect 27268 516 27324 572
rect 27324 516 27328 572
rect 27264 512 27328 516
rect 27344 572 27408 576
rect 27344 516 27348 572
rect 27348 516 27404 572
rect 27404 516 27408 572
rect 27344 512 27408 516
rect 27424 572 27488 576
rect 27424 516 27428 572
rect 27428 516 27484 572
rect 27484 516 27488 572
rect 27424 512 27488 516
rect 27504 572 27568 576
rect 27504 516 27508 572
rect 27508 516 27564 572
rect 27564 516 27568 572
rect 27504 512 27568 516
<< metal4 >>
rect 3750 17440 4070 17456
rect 3750 17376 3758 17440
rect 3822 17376 3838 17440
rect 3902 17376 3918 17440
rect 3982 17376 3998 17440
rect 4062 17376 4070 17440
rect 3750 16352 4070 17376
rect 3750 16288 3758 16352
rect 3822 16288 3838 16352
rect 3902 16288 3918 16352
rect 3982 16288 3998 16352
rect 4062 16288 4070 16352
rect 3750 15264 4070 16288
rect 3750 15200 3758 15264
rect 3822 15200 3838 15264
rect 3902 15200 3918 15264
rect 3982 15200 3998 15264
rect 4062 15200 4070 15264
rect 3750 14176 4070 15200
rect 3750 14112 3758 14176
rect 3822 14112 3838 14176
rect 3902 14112 3918 14176
rect 3982 14112 3998 14176
rect 4062 14112 4070 14176
rect 3750 13088 4070 14112
rect 3750 13024 3758 13088
rect 3822 13024 3838 13088
rect 3902 13024 3918 13088
rect 3982 13024 3998 13088
rect 4062 13024 4070 13088
rect 3750 12000 4070 13024
rect 3750 11936 3758 12000
rect 3822 11936 3838 12000
rect 3902 11936 3918 12000
rect 3982 11936 3998 12000
rect 4062 11936 4070 12000
rect 3750 10912 4070 11936
rect 3750 10848 3758 10912
rect 3822 10848 3838 10912
rect 3902 10848 3918 10912
rect 3982 10848 3998 10912
rect 4062 10848 4070 10912
rect 3750 9824 4070 10848
rect 3750 9760 3758 9824
rect 3822 9760 3838 9824
rect 3902 9760 3918 9824
rect 3982 9760 3998 9824
rect 4062 9760 4070 9824
rect 3750 8736 4070 9760
rect 3750 8672 3758 8736
rect 3822 8672 3838 8736
rect 3902 8672 3918 8736
rect 3982 8672 3998 8736
rect 4062 8672 4070 8736
rect 3750 7648 4070 8672
rect 3750 7584 3758 7648
rect 3822 7584 3838 7648
rect 3902 7584 3918 7648
rect 3982 7584 3998 7648
rect 4062 7584 4070 7648
rect 3750 6560 4070 7584
rect 3750 6496 3758 6560
rect 3822 6496 3838 6560
rect 3902 6496 3918 6560
rect 3982 6496 3998 6560
rect 4062 6496 4070 6560
rect 3750 5472 4070 6496
rect 3750 5408 3758 5472
rect 3822 5408 3838 5472
rect 3902 5408 3918 5472
rect 3982 5408 3998 5472
rect 4062 5408 4070 5472
rect 3750 4384 4070 5408
rect 3750 4320 3758 4384
rect 3822 4320 3838 4384
rect 3902 4320 3918 4384
rect 3982 4320 3998 4384
rect 4062 4320 4070 4384
rect 3750 3296 4070 4320
rect 3750 3232 3758 3296
rect 3822 3232 3838 3296
rect 3902 3232 3918 3296
rect 3982 3232 3998 3296
rect 4062 3232 4070 3296
rect 3750 2208 4070 3232
rect 3750 2144 3758 2208
rect 3822 2144 3838 2208
rect 3902 2144 3918 2208
rect 3982 2144 3998 2208
rect 4062 2144 4070 2208
rect 3750 1120 4070 2144
rect 3750 1056 3758 1120
rect 3822 1056 3838 1120
rect 3902 1056 3918 1120
rect 3982 1056 3998 1120
rect 4062 1056 4070 1120
rect 3750 496 4070 1056
rect 7108 16896 7428 17456
rect 7108 16832 7116 16896
rect 7180 16832 7196 16896
rect 7260 16832 7276 16896
rect 7340 16832 7356 16896
rect 7420 16832 7428 16896
rect 7108 15808 7428 16832
rect 7108 15744 7116 15808
rect 7180 15744 7196 15808
rect 7260 15744 7276 15808
rect 7340 15744 7356 15808
rect 7420 15744 7428 15808
rect 7108 14720 7428 15744
rect 7108 14656 7116 14720
rect 7180 14656 7196 14720
rect 7260 14656 7276 14720
rect 7340 14656 7356 14720
rect 7420 14656 7428 14720
rect 7108 13632 7428 14656
rect 7108 13568 7116 13632
rect 7180 13568 7196 13632
rect 7260 13568 7276 13632
rect 7340 13568 7356 13632
rect 7420 13568 7428 13632
rect 7108 12544 7428 13568
rect 7108 12480 7116 12544
rect 7180 12480 7196 12544
rect 7260 12480 7276 12544
rect 7340 12480 7356 12544
rect 7420 12480 7428 12544
rect 7108 11456 7428 12480
rect 10466 17440 10786 17456
rect 10466 17376 10474 17440
rect 10538 17376 10554 17440
rect 10618 17376 10634 17440
rect 10698 17376 10714 17440
rect 10778 17376 10786 17440
rect 10466 16352 10786 17376
rect 10466 16288 10474 16352
rect 10538 16288 10554 16352
rect 10618 16288 10634 16352
rect 10698 16288 10714 16352
rect 10778 16288 10786 16352
rect 10466 15264 10786 16288
rect 10466 15200 10474 15264
rect 10538 15200 10554 15264
rect 10618 15200 10634 15264
rect 10698 15200 10714 15264
rect 10778 15200 10786 15264
rect 10466 14176 10786 15200
rect 10466 14112 10474 14176
rect 10538 14112 10554 14176
rect 10618 14112 10634 14176
rect 10698 14112 10714 14176
rect 10778 14112 10786 14176
rect 10466 13088 10786 14112
rect 10466 13024 10474 13088
rect 10538 13024 10554 13088
rect 10618 13024 10634 13088
rect 10698 13024 10714 13088
rect 10778 13024 10786 13088
rect 10179 12204 10245 12205
rect 10179 12140 10180 12204
rect 10244 12140 10245 12204
rect 10179 12139 10245 12140
rect 7108 11392 7116 11456
rect 7180 11392 7196 11456
rect 7260 11392 7276 11456
rect 7340 11392 7356 11456
rect 7420 11392 7428 11456
rect 7108 10368 7428 11392
rect 7108 10304 7116 10368
rect 7180 10304 7196 10368
rect 7260 10304 7276 10368
rect 7340 10304 7356 10368
rect 7420 10304 7428 10368
rect 7108 9280 7428 10304
rect 10182 9621 10242 12139
rect 10466 12000 10786 13024
rect 10466 11936 10474 12000
rect 10538 11936 10554 12000
rect 10618 11936 10634 12000
rect 10698 11936 10714 12000
rect 10778 11936 10786 12000
rect 10466 10912 10786 11936
rect 10466 10848 10474 10912
rect 10538 10848 10554 10912
rect 10618 10848 10634 10912
rect 10698 10848 10714 10912
rect 10778 10848 10786 10912
rect 10466 9824 10786 10848
rect 10466 9760 10474 9824
rect 10538 9760 10554 9824
rect 10618 9760 10634 9824
rect 10698 9760 10714 9824
rect 10778 9760 10786 9824
rect 10179 9620 10245 9621
rect 10179 9556 10180 9620
rect 10244 9556 10245 9620
rect 10179 9555 10245 9556
rect 7108 9216 7116 9280
rect 7180 9216 7196 9280
rect 7260 9216 7276 9280
rect 7340 9216 7356 9280
rect 7420 9216 7428 9280
rect 7108 8192 7428 9216
rect 7108 8128 7116 8192
rect 7180 8128 7196 8192
rect 7260 8128 7276 8192
rect 7340 8128 7356 8192
rect 7420 8128 7428 8192
rect 7108 7104 7428 8128
rect 7108 7040 7116 7104
rect 7180 7040 7196 7104
rect 7260 7040 7276 7104
rect 7340 7040 7356 7104
rect 7420 7040 7428 7104
rect 7108 6016 7428 7040
rect 10182 6357 10242 9555
rect 10466 8736 10786 9760
rect 10466 8672 10474 8736
rect 10538 8672 10554 8736
rect 10618 8672 10634 8736
rect 10698 8672 10714 8736
rect 10778 8672 10786 8736
rect 10466 7648 10786 8672
rect 10466 7584 10474 7648
rect 10538 7584 10554 7648
rect 10618 7584 10634 7648
rect 10698 7584 10714 7648
rect 10778 7584 10786 7648
rect 10466 6560 10786 7584
rect 10466 6496 10474 6560
rect 10538 6496 10554 6560
rect 10618 6496 10634 6560
rect 10698 6496 10714 6560
rect 10778 6496 10786 6560
rect 10179 6356 10245 6357
rect 10179 6292 10180 6356
rect 10244 6292 10245 6356
rect 10179 6291 10245 6292
rect 7108 5952 7116 6016
rect 7180 5952 7196 6016
rect 7260 5952 7276 6016
rect 7340 5952 7356 6016
rect 7420 5952 7428 6016
rect 7108 4928 7428 5952
rect 7108 4864 7116 4928
rect 7180 4864 7196 4928
rect 7260 4864 7276 4928
rect 7340 4864 7356 4928
rect 7420 4864 7428 4928
rect 7108 3840 7428 4864
rect 7108 3776 7116 3840
rect 7180 3776 7196 3840
rect 7260 3776 7276 3840
rect 7340 3776 7356 3840
rect 7420 3776 7428 3840
rect 7108 2752 7428 3776
rect 7108 2688 7116 2752
rect 7180 2688 7196 2752
rect 7260 2688 7276 2752
rect 7340 2688 7356 2752
rect 7420 2688 7428 2752
rect 7108 1664 7428 2688
rect 7108 1600 7116 1664
rect 7180 1600 7196 1664
rect 7260 1600 7276 1664
rect 7340 1600 7356 1664
rect 7420 1600 7428 1664
rect 7108 576 7428 1600
rect 7108 512 7116 576
rect 7180 512 7196 576
rect 7260 512 7276 576
rect 7340 512 7356 576
rect 7420 512 7428 576
rect 7108 496 7428 512
rect 10466 5472 10786 6496
rect 10466 5408 10474 5472
rect 10538 5408 10554 5472
rect 10618 5408 10634 5472
rect 10698 5408 10714 5472
rect 10778 5408 10786 5472
rect 10466 4384 10786 5408
rect 10466 4320 10474 4384
rect 10538 4320 10554 4384
rect 10618 4320 10634 4384
rect 10698 4320 10714 4384
rect 10778 4320 10786 4384
rect 10466 3296 10786 4320
rect 10466 3232 10474 3296
rect 10538 3232 10554 3296
rect 10618 3232 10634 3296
rect 10698 3232 10714 3296
rect 10778 3232 10786 3296
rect 10466 2208 10786 3232
rect 10466 2144 10474 2208
rect 10538 2144 10554 2208
rect 10618 2144 10634 2208
rect 10698 2144 10714 2208
rect 10778 2144 10786 2208
rect 10466 1120 10786 2144
rect 10466 1056 10474 1120
rect 10538 1056 10554 1120
rect 10618 1056 10634 1120
rect 10698 1056 10714 1120
rect 10778 1056 10786 1120
rect 10466 496 10786 1056
rect 13824 16896 14144 17456
rect 13824 16832 13832 16896
rect 13896 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14144 16896
rect 13824 15808 14144 16832
rect 13824 15744 13832 15808
rect 13896 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14144 15808
rect 13824 14720 14144 15744
rect 13824 14656 13832 14720
rect 13896 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14144 14720
rect 13824 13632 14144 14656
rect 13824 13568 13832 13632
rect 13896 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14144 13632
rect 13824 12544 14144 13568
rect 13824 12480 13832 12544
rect 13896 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14144 12544
rect 13824 11456 14144 12480
rect 13824 11392 13832 11456
rect 13896 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14144 11456
rect 13824 10368 14144 11392
rect 13824 10304 13832 10368
rect 13896 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14144 10368
rect 13824 9280 14144 10304
rect 13824 9216 13832 9280
rect 13896 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14144 9280
rect 13824 8192 14144 9216
rect 13824 8128 13832 8192
rect 13896 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14144 8192
rect 13824 7104 14144 8128
rect 13824 7040 13832 7104
rect 13896 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14144 7104
rect 13824 6016 14144 7040
rect 13824 5952 13832 6016
rect 13896 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14144 6016
rect 13824 4928 14144 5952
rect 13824 4864 13832 4928
rect 13896 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14144 4928
rect 13824 3840 14144 4864
rect 13824 3776 13832 3840
rect 13896 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14144 3840
rect 13824 2752 14144 3776
rect 13824 2688 13832 2752
rect 13896 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14144 2752
rect 13824 1664 14144 2688
rect 13824 1600 13832 1664
rect 13896 1600 13912 1664
rect 13976 1600 13992 1664
rect 14056 1600 14072 1664
rect 14136 1600 14144 1664
rect 13824 576 14144 1600
rect 13824 512 13832 576
rect 13896 512 13912 576
rect 13976 512 13992 576
rect 14056 512 14072 576
rect 14136 512 14144 576
rect 13824 496 14144 512
rect 17182 17440 17502 17456
rect 17182 17376 17190 17440
rect 17254 17376 17270 17440
rect 17334 17376 17350 17440
rect 17414 17376 17430 17440
rect 17494 17376 17502 17440
rect 17182 16352 17502 17376
rect 17182 16288 17190 16352
rect 17254 16288 17270 16352
rect 17334 16288 17350 16352
rect 17414 16288 17430 16352
rect 17494 16288 17502 16352
rect 17182 15264 17502 16288
rect 20540 16896 20860 17456
rect 20540 16832 20548 16896
rect 20612 16832 20628 16896
rect 20692 16832 20708 16896
rect 20772 16832 20788 16896
rect 20852 16832 20860 16896
rect 20540 15808 20860 16832
rect 20540 15744 20548 15808
rect 20612 15744 20628 15808
rect 20692 15744 20708 15808
rect 20772 15744 20788 15808
rect 20852 15744 20860 15808
rect 17723 15468 17789 15469
rect 17723 15404 17724 15468
rect 17788 15404 17789 15468
rect 17723 15403 17789 15404
rect 17182 15200 17190 15264
rect 17254 15200 17270 15264
rect 17334 15200 17350 15264
rect 17414 15200 17430 15264
rect 17494 15200 17502 15264
rect 17182 14176 17502 15200
rect 17182 14112 17190 14176
rect 17254 14112 17270 14176
rect 17334 14112 17350 14176
rect 17414 14112 17430 14176
rect 17494 14112 17502 14176
rect 17182 13088 17502 14112
rect 17182 13024 17190 13088
rect 17254 13024 17270 13088
rect 17334 13024 17350 13088
rect 17414 13024 17430 13088
rect 17494 13024 17502 13088
rect 17182 12000 17502 13024
rect 17726 12613 17786 15403
rect 20540 14720 20860 15744
rect 20540 14656 20548 14720
rect 20612 14656 20628 14720
rect 20692 14656 20708 14720
rect 20772 14656 20788 14720
rect 20852 14656 20860 14720
rect 20540 13632 20860 14656
rect 23898 17440 24218 17456
rect 23898 17376 23906 17440
rect 23970 17376 23986 17440
rect 24050 17376 24066 17440
rect 24130 17376 24146 17440
rect 24210 17376 24218 17440
rect 23898 16352 24218 17376
rect 23898 16288 23906 16352
rect 23970 16288 23986 16352
rect 24050 16288 24066 16352
rect 24130 16288 24146 16352
rect 24210 16288 24218 16352
rect 23898 15264 24218 16288
rect 23898 15200 23906 15264
rect 23970 15200 23986 15264
rect 24050 15200 24066 15264
rect 24130 15200 24146 15264
rect 24210 15200 24218 15264
rect 23898 14176 24218 15200
rect 23898 14112 23906 14176
rect 23970 14112 23986 14176
rect 24050 14112 24066 14176
rect 24130 14112 24146 14176
rect 24210 14112 24218 14176
rect 22323 13836 22389 13837
rect 22323 13772 22324 13836
rect 22388 13772 22389 13836
rect 22323 13771 22389 13772
rect 20540 13568 20548 13632
rect 20612 13568 20628 13632
rect 20692 13568 20708 13632
rect 20772 13568 20788 13632
rect 20852 13568 20860 13632
rect 17723 12612 17789 12613
rect 17723 12548 17724 12612
rect 17788 12548 17789 12612
rect 17723 12547 17789 12548
rect 17182 11936 17190 12000
rect 17254 11936 17270 12000
rect 17334 11936 17350 12000
rect 17414 11936 17430 12000
rect 17494 11936 17502 12000
rect 17182 10912 17502 11936
rect 17182 10848 17190 10912
rect 17254 10848 17270 10912
rect 17334 10848 17350 10912
rect 17414 10848 17430 10912
rect 17494 10848 17502 10912
rect 17182 9824 17502 10848
rect 17182 9760 17190 9824
rect 17254 9760 17270 9824
rect 17334 9760 17350 9824
rect 17414 9760 17430 9824
rect 17494 9760 17502 9824
rect 17182 8736 17502 9760
rect 17182 8672 17190 8736
rect 17254 8672 17270 8736
rect 17334 8672 17350 8736
rect 17414 8672 17430 8736
rect 17494 8672 17502 8736
rect 17182 7648 17502 8672
rect 17726 8397 17786 12547
rect 20540 12544 20860 13568
rect 20540 12480 20548 12544
rect 20612 12480 20628 12544
rect 20692 12480 20708 12544
rect 20772 12480 20788 12544
rect 20852 12480 20860 12544
rect 18643 11524 18709 11525
rect 18643 11460 18644 11524
rect 18708 11460 18709 11524
rect 18643 11459 18709 11460
rect 18275 11116 18341 11117
rect 18275 11052 18276 11116
rect 18340 11052 18341 11116
rect 18275 11051 18341 11052
rect 17723 8396 17789 8397
rect 17723 8332 17724 8396
rect 17788 8332 17789 8396
rect 17723 8331 17789 8332
rect 17182 7584 17190 7648
rect 17254 7584 17270 7648
rect 17334 7584 17350 7648
rect 17414 7584 17430 7648
rect 17494 7584 17502 7648
rect 17182 6560 17502 7584
rect 17182 6496 17190 6560
rect 17254 6496 17270 6560
rect 17334 6496 17350 6560
rect 17414 6496 17430 6560
rect 17494 6496 17502 6560
rect 17182 5472 17502 6496
rect 17182 5408 17190 5472
rect 17254 5408 17270 5472
rect 17334 5408 17350 5472
rect 17414 5408 17430 5472
rect 17494 5408 17502 5472
rect 17182 4384 17502 5408
rect 17182 4320 17190 4384
rect 17254 4320 17270 4384
rect 17334 4320 17350 4384
rect 17414 4320 17430 4384
rect 17494 4320 17502 4384
rect 17182 3296 17502 4320
rect 18278 4045 18338 11051
rect 18646 9621 18706 11459
rect 20540 11456 20860 12480
rect 20540 11392 20548 11456
rect 20612 11392 20628 11456
rect 20692 11392 20708 11456
rect 20772 11392 20788 11456
rect 20852 11392 20860 11456
rect 20540 10368 20860 11392
rect 20540 10304 20548 10368
rect 20612 10304 20628 10368
rect 20692 10304 20708 10368
rect 20772 10304 20788 10368
rect 20852 10304 20860 10368
rect 18643 9620 18709 9621
rect 18643 9556 18644 9620
rect 18708 9556 18709 9620
rect 18643 9555 18709 9556
rect 20299 9620 20365 9621
rect 20299 9556 20300 9620
rect 20364 9556 20365 9620
rect 20299 9555 20365 9556
rect 20302 5269 20362 9555
rect 20540 9280 20860 10304
rect 20540 9216 20548 9280
rect 20612 9216 20628 9280
rect 20692 9216 20708 9280
rect 20772 9216 20788 9280
rect 20852 9216 20860 9280
rect 20540 8192 20860 9216
rect 20540 8128 20548 8192
rect 20612 8128 20628 8192
rect 20692 8128 20708 8192
rect 20772 8128 20788 8192
rect 20852 8128 20860 8192
rect 20540 7104 20860 8128
rect 20540 7040 20548 7104
rect 20612 7040 20628 7104
rect 20692 7040 20708 7104
rect 20772 7040 20788 7104
rect 20852 7040 20860 7104
rect 20540 6016 20860 7040
rect 20540 5952 20548 6016
rect 20612 5952 20628 6016
rect 20692 5952 20708 6016
rect 20772 5952 20788 6016
rect 20852 5952 20860 6016
rect 20299 5268 20365 5269
rect 20299 5204 20300 5268
rect 20364 5204 20365 5268
rect 20299 5203 20365 5204
rect 20540 4928 20860 5952
rect 20540 4864 20548 4928
rect 20612 4864 20628 4928
rect 20692 4864 20708 4928
rect 20772 4864 20788 4928
rect 20852 4864 20860 4928
rect 18275 4044 18341 4045
rect 18275 3980 18276 4044
rect 18340 3980 18341 4044
rect 18275 3979 18341 3980
rect 17182 3232 17190 3296
rect 17254 3232 17270 3296
rect 17334 3232 17350 3296
rect 17414 3232 17430 3296
rect 17494 3232 17502 3296
rect 17182 2208 17502 3232
rect 17182 2144 17190 2208
rect 17254 2144 17270 2208
rect 17334 2144 17350 2208
rect 17414 2144 17430 2208
rect 17494 2144 17502 2208
rect 17182 1120 17502 2144
rect 17182 1056 17190 1120
rect 17254 1056 17270 1120
rect 17334 1056 17350 1120
rect 17414 1056 17430 1120
rect 17494 1056 17502 1120
rect 17182 496 17502 1056
rect 20540 3840 20860 4864
rect 22326 4045 22386 13771
rect 23898 13088 24218 14112
rect 23898 13024 23906 13088
rect 23970 13024 23986 13088
rect 24050 13024 24066 13088
rect 24130 13024 24146 13088
rect 24210 13024 24218 13088
rect 23898 12000 24218 13024
rect 27256 16896 27576 17456
rect 27256 16832 27264 16896
rect 27328 16832 27344 16896
rect 27408 16832 27424 16896
rect 27488 16832 27504 16896
rect 27568 16832 27576 16896
rect 27256 15808 27576 16832
rect 27256 15744 27264 15808
rect 27328 15744 27344 15808
rect 27408 15744 27424 15808
rect 27488 15744 27504 15808
rect 27568 15744 27576 15808
rect 27256 14720 27576 15744
rect 27256 14656 27264 14720
rect 27328 14656 27344 14720
rect 27408 14656 27424 14720
rect 27488 14656 27504 14720
rect 27568 14656 27576 14720
rect 27256 13632 27576 14656
rect 27256 13568 27264 13632
rect 27328 13568 27344 13632
rect 27408 13568 27424 13632
rect 27488 13568 27504 13632
rect 27568 13568 27576 13632
rect 27256 12544 27576 13568
rect 27256 12480 27264 12544
rect 27328 12480 27344 12544
rect 27408 12480 27424 12544
rect 27488 12480 27504 12544
rect 27568 12480 27576 12544
rect 26187 12340 26253 12341
rect 26187 12276 26188 12340
rect 26252 12276 26253 12340
rect 26187 12275 26253 12276
rect 23898 11936 23906 12000
rect 23970 11936 23986 12000
rect 24050 11936 24066 12000
rect 24130 11936 24146 12000
rect 24210 11936 24218 12000
rect 23898 10912 24218 11936
rect 23898 10848 23906 10912
rect 23970 10848 23986 10912
rect 24050 10848 24066 10912
rect 24130 10848 24146 10912
rect 24210 10848 24218 10912
rect 23898 9824 24218 10848
rect 23898 9760 23906 9824
rect 23970 9760 23986 9824
rect 24050 9760 24066 9824
rect 24130 9760 24146 9824
rect 24210 9760 24218 9824
rect 23898 8736 24218 9760
rect 26190 9485 26250 12275
rect 27256 11456 27576 12480
rect 27256 11392 27264 11456
rect 27328 11392 27344 11456
rect 27408 11392 27424 11456
rect 27488 11392 27504 11456
rect 27568 11392 27576 11456
rect 27256 10368 27576 11392
rect 27256 10304 27264 10368
rect 27328 10304 27344 10368
rect 27408 10304 27424 10368
rect 27488 10304 27504 10368
rect 27568 10304 27576 10368
rect 26187 9484 26253 9485
rect 26187 9420 26188 9484
rect 26252 9420 26253 9484
rect 26187 9419 26253 9420
rect 23898 8672 23906 8736
rect 23970 8672 23986 8736
rect 24050 8672 24066 8736
rect 24130 8672 24146 8736
rect 24210 8672 24218 8736
rect 23898 7648 24218 8672
rect 23898 7584 23906 7648
rect 23970 7584 23986 7648
rect 24050 7584 24066 7648
rect 24130 7584 24146 7648
rect 24210 7584 24218 7648
rect 23898 6560 24218 7584
rect 23898 6496 23906 6560
rect 23970 6496 23986 6560
rect 24050 6496 24066 6560
rect 24130 6496 24146 6560
rect 24210 6496 24218 6560
rect 23898 5472 24218 6496
rect 23898 5408 23906 5472
rect 23970 5408 23986 5472
rect 24050 5408 24066 5472
rect 24130 5408 24146 5472
rect 24210 5408 24218 5472
rect 23898 4384 24218 5408
rect 23898 4320 23906 4384
rect 23970 4320 23986 4384
rect 24050 4320 24066 4384
rect 24130 4320 24146 4384
rect 24210 4320 24218 4384
rect 22323 4044 22389 4045
rect 22323 3980 22324 4044
rect 22388 3980 22389 4044
rect 22323 3979 22389 3980
rect 20540 3776 20548 3840
rect 20612 3776 20628 3840
rect 20692 3776 20708 3840
rect 20772 3776 20788 3840
rect 20852 3776 20860 3840
rect 20540 2752 20860 3776
rect 20540 2688 20548 2752
rect 20612 2688 20628 2752
rect 20692 2688 20708 2752
rect 20772 2688 20788 2752
rect 20852 2688 20860 2752
rect 20540 1664 20860 2688
rect 20540 1600 20548 1664
rect 20612 1600 20628 1664
rect 20692 1600 20708 1664
rect 20772 1600 20788 1664
rect 20852 1600 20860 1664
rect 20540 576 20860 1600
rect 20540 512 20548 576
rect 20612 512 20628 576
rect 20692 512 20708 576
rect 20772 512 20788 576
rect 20852 512 20860 576
rect 20540 496 20860 512
rect 23898 3296 24218 4320
rect 23898 3232 23906 3296
rect 23970 3232 23986 3296
rect 24050 3232 24066 3296
rect 24130 3232 24146 3296
rect 24210 3232 24218 3296
rect 23898 2208 24218 3232
rect 23898 2144 23906 2208
rect 23970 2144 23986 2208
rect 24050 2144 24066 2208
rect 24130 2144 24146 2208
rect 24210 2144 24218 2208
rect 23898 1120 24218 2144
rect 23898 1056 23906 1120
rect 23970 1056 23986 1120
rect 24050 1056 24066 1120
rect 24130 1056 24146 1120
rect 24210 1056 24218 1120
rect 23898 496 24218 1056
rect 27256 9280 27576 10304
rect 27256 9216 27264 9280
rect 27328 9216 27344 9280
rect 27408 9216 27424 9280
rect 27488 9216 27504 9280
rect 27568 9216 27576 9280
rect 27256 8192 27576 9216
rect 27256 8128 27264 8192
rect 27328 8128 27344 8192
rect 27408 8128 27424 8192
rect 27488 8128 27504 8192
rect 27568 8128 27576 8192
rect 27256 7104 27576 8128
rect 27256 7040 27264 7104
rect 27328 7040 27344 7104
rect 27408 7040 27424 7104
rect 27488 7040 27504 7104
rect 27568 7040 27576 7104
rect 27256 6016 27576 7040
rect 27256 5952 27264 6016
rect 27328 5952 27344 6016
rect 27408 5952 27424 6016
rect 27488 5952 27504 6016
rect 27568 5952 27576 6016
rect 27256 4928 27576 5952
rect 27256 4864 27264 4928
rect 27328 4864 27344 4928
rect 27408 4864 27424 4928
rect 27488 4864 27504 4928
rect 27568 4864 27576 4928
rect 27256 3840 27576 4864
rect 27256 3776 27264 3840
rect 27328 3776 27344 3840
rect 27408 3776 27424 3840
rect 27488 3776 27504 3840
rect 27568 3776 27576 3840
rect 27256 2752 27576 3776
rect 27256 2688 27264 2752
rect 27328 2688 27344 2752
rect 27408 2688 27424 2752
rect 27488 2688 27504 2752
rect 27568 2688 27576 2752
rect 27256 1664 27576 2688
rect 27256 1600 27264 1664
rect 27328 1600 27344 1664
rect 27408 1600 27424 1664
rect 27488 1600 27504 1664
rect 27568 1600 27576 1664
rect 27256 576 27576 1600
rect 27256 512 27264 576
rect 27328 512 27344 576
rect 27408 512 27424 576
rect 27488 512 27504 576
rect 27568 512 27576 576
rect 27256 496 27576 512
use sky130_fd_sc_hd__inv_2  _382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16376 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _383_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15824 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _384_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15548 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _385_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _386_
timestamp 1704896540
transform 1 0 9752 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1704896540
transform 1 0 25484 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1704896540
transform 1 0 25208 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _389_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 18124 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _390_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 25668 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 25668 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _392_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 24748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _393_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 26864 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _394_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 24748 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _395_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22908 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _396_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 23460 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 24748 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _398_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 25300 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _399_
timestamp 1704896540
transform 1 0 21988 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _400_
timestamp 1704896540
transform -1 0 23368 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _401_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17756 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _402_
timestamp 1704896540
transform 1 0 17572 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _403_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21804 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _404_
timestamp 1704896540
transform 1 0 17940 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _405_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 23276 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _406_
timestamp 1704896540
transform -1 0 22724 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _407_
timestamp 1704896540
transform -1 0 23460 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _408_
timestamp 1704896540
transform -1 0 23184 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _409_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22172 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _410_
timestamp 1704896540
transform 1 0 23184 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _411_
timestamp 1704896540
transform -1 0 24564 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _412_
timestamp 1704896540
transform 1 0 17020 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _413_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2116 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _414_
timestamp 1704896540
transform -1 0 1932 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _415_
timestamp 1704896540
transform -1 0 16008 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _416_
timestamp 1704896540
transform -1 0 10672 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17480 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _418_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 19964 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_4  _419_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15640 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1704896540
transform -1 0 14904 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _421_
timestamp 1704896540
transform 1 0 23460 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _422_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4324 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_2  _423_
timestamp 1704896540
transform -1 0 23276 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _424_
timestamp 1704896540
transform 1 0 4416 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_2  _425_
timestamp 1704896540
transform -1 0 23184 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _426_
timestamp 1704896540
transform 1 0 5612 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_2  _427_
timestamp 1704896540
transform -1 0 23460 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _428_
timestamp 1704896540
transform 1 0 7360 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_2  _429_
timestamp 1704896540
transform -1 0 22908 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _430_
timestamp 1704896540
transform 1 0 9108 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_2  _431_
timestamp 1704896540
transform -1 0 22356 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _432_
timestamp 1704896540
transform 1 0 10672 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_2  _433_
timestamp 1704896540
transform 1 0 21252 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _434_
timestamp 1704896540
transform 1 0 12788 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__a2bb2o_4  _435_
timestamp 1704896540
transform 1 0 14260 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  _436_
timestamp 1704896540
transform 1 0 16100 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _437_
timestamp 1704896540
transform 1 0 16100 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _438_
timestamp 1704896540
transform -1 0 18768 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _439_
timestamp 1704896540
transform -1 0 20700 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _440_
timestamp 1704896540
transform -1 0 22540 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _441_
timestamp 1704896540
transform -1 0 22264 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _442_
timestamp 1704896540
transform -1 0 22540 0 1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _443_
timestamp 1704896540
transform -1 0 22540 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _444_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14536 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _445_
timestamp 1704896540
transform -1 0 14720 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _446_
timestamp 1704896540
transform 1 0 16100 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _447_
timestamp 1704896540
transform 1 0 15088 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _448_
timestamp 1704896540
transform 1 0 14720 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _449_
timestamp 1704896540
transform -1 0 14536 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _450_
timestamp 1704896540
transform 1 0 14720 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _451_
timestamp 1704896540
transform 1 0 14536 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _452_
timestamp 1704896540
transform -1 0 14076 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _453_
timestamp 1704896540
transform 1 0 14444 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _454_
timestamp 1704896540
transform 1 0 13892 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _455_
timestamp 1704896540
transform -1 0 13708 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _456_
timestamp 1704896540
transform 1 0 13524 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _457_
timestamp 1704896540
transform 1 0 12604 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _458_
timestamp 1704896540
transform 1 0 12696 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _459_
timestamp 1704896540
transform 1 0 13156 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _460_
timestamp 1704896540
transform 1 0 12328 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _461_
timestamp 1704896540
transform 1 0 12236 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp 1704896540
transform 1 0 13156 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _463_
timestamp 1704896540
transform 1 0 12328 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _464_
timestamp 1704896540
transform -1 0 11776 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _465_
timestamp 1704896540
transform 1 0 13064 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _466_
timestamp 1704896540
transform -1 0 15180 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _467_
timestamp 1704896540
transform 1 0 11960 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _468_
timestamp 1704896540
transform -1 0 11408 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _469_
timestamp 1704896540
transform -1 0 6992 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _470_
timestamp 1704896540
transform -1 0 6532 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_2  _471_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17296 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _472_
timestamp 1704896540
transform -1 0 5520 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _473_
timestamp 1704896540
transform -1 0 4232 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _474_
timestamp 1704896540
transform -1 0 19044 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _475_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4600 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _476_
timestamp 1704896540
transform -1 0 3404 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _477_
timestamp 1704896540
transform -1 0 5152 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _478_
timestamp 1704896540
transform -1 0 24104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _479_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3128 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _480_
timestamp 1704896540
transform 1 0 2484 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _481_
timestamp 1704896540
transform -1 0 1932 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _482_
timestamp 1704896540
transform 1 0 3956 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _483_
timestamp 1704896540
transform -1 0 2300 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _484_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6164 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _485_
timestamp 1704896540
transform 1 0 4876 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4600 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _487_
timestamp 1704896540
transform 1 0 5244 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _488_
timestamp 1704896540
transform -1 0 4140 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _489_
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _490_
timestamp 1704896540
transform 1 0 3404 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _491_
timestamp 1704896540
transform -1 0 4692 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _492_
timestamp 1704896540
transform -1 0 5336 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _493_
timestamp 1704896540
transform -1 0 4600 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _494_
timestamp 1704896540
transform -1 0 6440 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _495_
timestamp 1704896540
transform -1 0 5704 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _496_
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _497_
timestamp 1704896540
transform -1 0 7544 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _498_
timestamp 1704896540
transform 1 0 5336 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _499_
timestamp 1704896540
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _500_
timestamp 1704896540
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _501_
timestamp 1704896540
transform 1 0 7820 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _502_
timestamp 1704896540
transform 1 0 7544 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _503_
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _504_
timestamp 1704896540
transform 1 0 8464 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _505_
timestamp 1704896540
transform 1 0 9476 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _506_
timestamp 1704896540
transform -1 0 9292 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_1  _507_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7360 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _508_
timestamp 1704896540
transform -1 0 6716 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _509_
timestamp 1704896540
transform -1 0 6440 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _510_
timestamp 1704896540
transform -1 0 7084 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _511_
timestamp 1704896540
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _512_
timestamp 1704896540
transform -1 0 6532 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _513_
timestamp 1704896540
transform -1 0 5704 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _514_
timestamp 1704896540
transform 1 0 5244 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _515_
timestamp 1704896540
transform 1 0 8096 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _516_
timestamp 1704896540
transform 1 0 8556 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _517_
timestamp 1704896540
transform 1 0 8372 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _518_
timestamp 1704896540
transform -1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _519_
timestamp 1704896540
transform -1 0 8648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _520_
timestamp 1704896540
transform -1 0 10212 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _521_
timestamp 1704896540
transform -1 0 9200 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _522_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6808 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _523_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7912 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _524_
timestamp 1704896540
transform -1 0 8280 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _525_
timestamp 1704896540
transform -1 0 7728 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _526_
timestamp 1704896540
transform -1 0 10028 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _527_
timestamp 1704896540
transform -1 0 10304 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _528_
timestamp 1704896540
transform -1 0 9936 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _529_
timestamp 1704896540
transform 1 0 9200 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _530_
timestamp 1704896540
transform 1 0 11224 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _531_
timestamp 1704896540
transform 1 0 13064 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _532_
timestamp 1704896540
transform 1 0 13800 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _533_
timestamp 1704896540
transform -1 0 11316 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _534_
timestamp 1704896540
transform 1 0 11316 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _535_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11224 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _536_
timestamp 1704896540
transform -1 0 12696 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _537_
timestamp 1704896540
transform 1 0 10120 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _538_
timestamp 1704896540
transform 1 0 10396 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _539_
timestamp 1704896540
transform -1 0 13800 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _540_
timestamp 1704896540
transform -1 0 12696 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _541_
timestamp 1704896540
transform -1 0 12788 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _542_
timestamp 1704896540
transform -1 0 12604 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _543_
timestamp 1704896540
transform -1 0 13616 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _544_
timestamp 1704896540
transform -1 0 12420 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _545_
timestamp 1704896540
transform 1 0 12420 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _546_
timestamp 1704896540
transform -1 0 11776 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1704896540
transform -1 0 11040 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _548_
timestamp 1704896540
transform 1 0 13800 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _549_
timestamp 1704896540
transform -1 0 12236 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _550_
timestamp 1704896540
transform 1 0 11224 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _551_
timestamp 1704896540
transform 1 0 11684 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _552_
timestamp 1704896540
transform -1 0 11224 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _553_
timestamp 1704896540
transform -1 0 24380 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _554_
timestamp 1704896540
transform -1 0 24380 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _555_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 23276 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _556_
timestamp 1704896540
transform -1 0 23368 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _557_
timestamp 1704896540
transform -1 0 22172 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _558_
timestamp 1704896540
transform 1 0 22540 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _559_
timestamp 1704896540
transform 1 0 21804 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _560_
timestamp 1704896540
transform 1 0 25668 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 23920 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _562_
timestamp 1704896540
transform 1 0 24748 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _563_
timestamp 1704896540
transform -1 0 17296 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _564_
timestamp 1704896540
transform 1 0 16284 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _565_
timestamp 1704896540
transform 1 0 23460 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _566_
timestamp 1704896540
transform -1 0 24380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _567_
timestamp 1704896540
transform 1 0 25300 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _568_
timestamp 1704896540
transform 1 0 24840 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _569_
timestamp 1704896540
transform -1 0 25392 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _570_
timestamp 1704896540
transform 1 0 25116 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _571_
timestamp 1704896540
transform 1 0 24564 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _572_
timestamp 1704896540
transform -1 0 26220 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _573_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 25944 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _574_
timestamp 1704896540
transform 1 0 25760 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _575_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 25760 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _576_
timestamp 1704896540
transform -1 0 25852 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _577_
timestamp 1704896540
transform -1 0 26312 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _578_
timestamp 1704896540
transform 1 0 24380 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _579_
timestamp 1704896540
transform 1 0 25852 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _580_
timestamp 1704896540
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _581_
timestamp 1704896540
transform -1 0 24380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _582_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _583_
timestamp 1704896540
transform 1 0 24564 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _584_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 24748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _585_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 23644 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _586_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 23828 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _587_
timestamp 1704896540
transform 1 0 17388 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _588_
timestamp 1704896540
transform -1 0 23736 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _589_
timestamp 1704896540
transform 1 0 24564 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _590_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 24564 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _591_
timestamp 1704896540
transform 1 0 19596 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _592_
timestamp 1704896540
transform -1 0 20700 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _593_
timestamp 1704896540
transform -1 0 23736 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _594_
timestamp 1704896540
transform -1 0 20424 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 20056 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _596_
timestamp 1704896540
transform -1 0 24932 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _597_
timestamp 1704896540
transform -1 0 24472 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _598_
timestamp 1704896540
transform -1 0 20608 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _599_
timestamp 1704896540
transform 1 0 19228 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21344 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _601_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17940 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _602_
timestamp 1704896540
transform -1 0 24104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _603_
timestamp 1704896540
transform 1 0 17112 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _604_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18308 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _605_
timestamp 1704896540
transform 1 0 19872 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _606_
timestamp 1704896540
transform -1 0 21160 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _607_
timestamp 1704896540
transform 1 0 11132 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _608_
timestamp 1704896540
transform -1 0 12696 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _609_
timestamp 1704896540
transform 1 0 11224 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _610_
timestamp 1704896540
transform -1 0 13432 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _611_
timestamp 1704896540
transform 1 0 11040 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _612_
timestamp 1704896540
transform -1 0 12512 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _613_
timestamp 1704896540
transform 1 0 11500 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _614_
timestamp 1704896540
transform -1 0 14260 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _615_
timestamp 1704896540
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _616_
timestamp 1704896540
transform 1 0 16836 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _617_
timestamp 1704896540
transform 1 0 11960 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _618_
timestamp 1704896540
transform -1 0 13432 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _619_
timestamp 1704896540
transform 1 0 11316 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _620_
timestamp 1704896540
transform 1 0 12236 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _621_
timestamp 1704896540
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _622_
timestamp 1704896540
transform -1 0 14996 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _623_
timestamp 1704896540
transform 1 0 16008 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _624_
timestamp 1704896540
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _625_
timestamp 1704896540
transform 1 0 18676 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _626_
timestamp 1704896540
transform 1 0 23092 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _627_
timestamp 1704896540
transform -1 0 22908 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _628_
timestamp 1704896540
transform 1 0 18860 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _629_
timestamp 1704896540
transform -1 0 20884 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _630_
timestamp 1704896540
transform -1 0 23644 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _631_
timestamp 1704896540
transform 1 0 21988 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _632_
timestamp 1704896540
transform 1 0 20240 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _633_
timestamp 1704896540
transform 1 0 21988 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _634_
timestamp 1704896540
transform -1 0 24564 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _635_
timestamp 1704896540
transform -1 0 22724 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _636_
timestamp 1704896540
transform -1 0 21988 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _637_
timestamp 1704896540
transform 1 0 21252 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _638_
timestamp 1704896540
transform -1 0 22724 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _639_
timestamp 1704896540
transform -1 0 22264 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _640_
timestamp 1704896540
transform 1 0 22264 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _641_
timestamp 1704896540
transform -1 0 23736 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _642_
timestamp 1704896540
transform 1 0 24564 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _643_
timestamp 1704896540
transform -1 0 26772 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _644_
timestamp 1704896540
transform 1 0 23828 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _645_
timestamp 1704896540
transform -1 0 26036 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _646_
timestamp 1704896540
transform 1 0 22724 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _647_
timestamp 1704896540
transform -1 0 24564 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _648_
timestamp 1704896540
transform 1 0 22356 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _649_
timestamp 1704896540
transform 1 0 16744 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _650_
timestamp 1704896540
transform -1 0 24196 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _651_
timestamp 1704896540
transform 1 0 22356 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _652_
timestamp 1704896540
transform -1 0 23644 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _653_
timestamp 1704896540
transform 1 0 21252 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _654_
timestamp 1704896540
transform -1 0 22540 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _655_
timestamp 1704896540
transform -1 0 21620 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _656_
timestamp 1704896540
transform -1 0 21160 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _657_
timestamp 1704896540
transform -1 0 18492 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _658_
timestamp 1704896540
transform -1 0 18584 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _659_
timestamp 1704896540
transform -1 0 18492 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _660_
timestamp 1704896540
transform 1 0 5428 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _661_
timestamp 1704896540
transform -1 0 17480 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _662_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16284 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _663_
timestamp 1704896540
transform 1 0 5796 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _664_
timestamp 1704896540
transform -1 0 8648 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _665_
timestamp 1704896540
transform 1 0 7176 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _666_
timestamp 1704896540
transform 1 0 5796 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _667_
timestamp 1704896540
transform -1 0 9108 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _668_
timestamp 1704896540
transform -1 0 8280 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _669_
timestamp 1704896540
transform 1 0 6164 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _670_
timestamp 1704896540
transform -1 0 10120 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _671_
timestamp 1704896540
transform -1 0 7544 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _672_
timestamp 1704896540
transform 1 0 6164 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _673_
timestamp 1704896540
transform -1 0 10120 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _674_
timestamp 1704896540
transform 1 0 8372 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _675_
timestamp 1704896540
transform 1 0 6624 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _676_
timestamp 1704896540
transform -1 0 9568 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _677_
timestamp 1704896540
transform -1 0 8188 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _678_
timestamp 1704896540
transform 1 0 7452 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _679_
timestamp 1704896540
transform -1 0 13984 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _680_
timestamp 1704896540
transform 1 0 11224 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _681_
timestamp 1704896540
transform -1 0 9384 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _682_
timestamp 1704896540
transform -1 0 10120 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _683_
timestamp 1704896540
transform 1 0 8648 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _684_
timestamp 1704896540
transform -1 0 9200 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _685_
timestamp 1704896540
transform 1 0 13064 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _686_
timestamp 1704896540
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _687_
timestamp 1704896540
transform -1 0 14904 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _688_
timestamp 1704896540
transform 1 0 14904 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _689_
timestamp 1704896540
transform -1 0 14904 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _690_
timestamp 1704896540
transform 1 0 16836 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _691_
timestamp 1704896540
transform -1 0 14536 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _692_
timestamp 1704896540
transform 1 0 14812 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _693_
timestamp 1704896540
transform -1 0 14812 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _694_
timestamp 1704896540
transform 1 0 15916 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _695_
timestamp 1704896540
transform -1 0 16652 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _696_
timestamp 1704896540
transform -1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _697_
timestamp 1704896540
transform -1 0 16008 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _698_
timestamp 1704896540
transform -1 0 15272 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _699_
timestamp 1704896540
transform -1 0 15640 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _700_
timestamp 1704896540
transform -1 0 14352 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _701_
timestamp 1704896540
transform 1 0 16836 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _702_
timestamp 1704896540
transform -1 0 14904 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _703_
timestamp 1704896540
transform -1 0 20148 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _704_
timestamp 1704896540
transform -1 0 15180 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _705_
timestamp 1704896540
transform 1 0 18676 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _706_
timestamp 1704896540
transform -1 0 15824 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _707_
timestamp 1704896540
transform -1 0 18584 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _708_
timestamp 1704896540
transform 1 0 12420 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _709_
timestamp 1704896540
transform -1 0 13064 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _710_
timestamp 1704896540
transform -1 0 19136 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _711_
timestamp 1704896540
transform -1 0 13616 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _712_
timestamp 1704896540
transform 1 0 16836 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _713_
timestamp 1704896540
transform -1 0 14812 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _714_
timestamp 1704896540
transform -1 0 18584 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _715_
timestamp 1704896540
transform -1 0 14260 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _716_
timestamp 1704896540
transform -1 0 18400 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _717_
timestamp 1704896540
transform 1 0 16560 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17112 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _719_
timestamp 1704896540
transform 1 0 17756 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _720_
timestamp 1704896540
transform 1 0 19964 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _721_
timestamp 1704896540
transform 1 0 20332 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _722_
timestamp 1704896540
transform 1 0 9476 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _723_
timestamp 1704896540
transform 1 0 10120 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _724_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9752 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _725_
timestamp 1704896540
transform 1 0 5796 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _726_
timestamp 1704896540
transform -1 0 10120 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _727_
timestamp 1704896540
transform 1 0 7268 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _728_
timestamp 1704896540
transform -1 0 10488 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _729_
timestamp 1704896540
transform 1 0 5336 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _730_
timestamp 1704896540
transform -1 0 10120 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _731_
timestamp 1704896540
transform 1 0 4968 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _732_
timestamp 1704896540
transform -1 0 10764 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _733_
timestamp 1704896540
transform 1 0 5060 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _734_
timestamp 1704896540
transform -1 0 9844 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _735_
timestamp 1704896540
transform 1 0 8372 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _736_
timestamp 1704896540
transform 1 0 11316 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _737_
timestamp 1704896540
transform 1 0 10672 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _738_
timestamp 1704896540
transform 1 0 11224 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _739_
timestamp 1704896540
transform 1 0 10948 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _740_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9292 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _741_
timestamp 1704896540
transform 1 0 8648 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _742_
timestamp 1704896540
transform -1 0 18124 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _743_
timestamp 1704896540
transform -1 0 4876 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _744_
timestamp 1704896540
transform -1 0 3680 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _745_
timestamp 1704896540
transform -1 0 3036 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _746_
timestamp 1704896540
transform -1 0 5520 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _747_
timestamp 1704896540
transform 1 0 4600 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _748_
timestamp 1704896540
transform 1 0 5796 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _749_
timestamp 1704896540
transform -1 0 4784 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _750_
timestamp 1704896540
transform -1 0 4140 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _751_
timestamp 1704896540
transform 1 0 2852 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _752_
timestamp 1704896540
transform -1 0 4876 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _753_
timestamp 1704896540
transform -1 0 3772 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _754_
timestamp 1704896540
transform -1 0 3128 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _755_
timestamp 1704896540
transform -1 0 4968 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _756_
timestamp 1704896540
transform -1 0 4232 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _757_
timestamp 1704896540
transform 1 0 2760 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _758_
timestamp 1704896540
transform 1 0 16744 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _759_
timestamp 1704896540
transform -1 0 9752 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _760_
timestamp 1704896540
transform 1 0 7820 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _761_
timestamp 1704896540
transform 1 0 8372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _762_
timestamp 1704896540
transform 1 0 11684 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _763_
timestamp 1704896540
transform -1 0 12512 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _764_
timestamp 1704896540
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _765_
timestamp 1704896540
transform 1 0 12420 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _766_
timestamp 1704896540
transform 1 0 12512 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _767_
timestamp 1704896540
transform -1 0 13248 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _768_
timestamp 1704896540
transform 1 0 9476 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _769_
timestamp 1704896540
transform -1 0 10580 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _770_
timestamp 1704896540
transform -1 0 8924 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _771_
timestamp 1704896540
transform 1 0 17204 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _772_
timestamp 1704896540
transform 1 0 17848 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _773_
timestamp 1704896540
transform -1 0 18584 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _774_
timestamp 1704896540
transform 1 0 16100 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _775_
timestamp 1704896540
transform -1 0 17204 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _776_
timestamp 1704896540
transform -1 0 16192 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _777_
timestamp 1704896540
transform 1 0 16008 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _778_
timestamp 1704896540
transform 1 0 16928 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _779_
timestamp 1704896540
transform -1 0 18584 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _780_
timestamp 1704896540
transform 1 0 17572 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _781_
timestamp 1704896540
transform 1 0 18124 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _782_
timestamp 1704896540
transform -1 0 19412 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _783_
timestamp 1704896540
transform 1 0 16928 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _784_
timestamp 1704896540
transform 1 0 18676 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _785_
timestamp 1704896540
transform -1 0 19596 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _786_
timestamp 1704896540
transform 1 0 17112 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _787_
timestamp 1704896540
transform 1 0 18400 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _788_
timestamp 1704896540
transform -1 0 19688 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _789_
timestamp 1704896540
transform 1 0 17664 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _790_
timestamp 1704896540
transform 1 0 18676 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _791_
timestamp 1704896540
transform -1 0 19228 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _792_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3220 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _793_
timestamp 1704896540
transform 1 0 1656 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _794_
timestamp 1704896540
transform 1 0 1472 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _795_
timestamp 1704896540
transform 1 0 4232 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _796_
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _797_
timestamp 1704896540
transform 1 0 3496 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _798_
timestamp 1704896540
transform 1 0 5796 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _799_
timestamp 1704896540
transform -1 0 5704 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _800_
timestamp 1704896540
transform 1 0 8280 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _801_
timestamp 1704896540
transform 1 0 6808 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _802_
timestamp 1704896540
transform 1 0 4600 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _803_
timestamp 1704896540
transform 1 0 4600 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _804_
timestamp 1704896540
transform 1 0 9016 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _805_
timestamp 1704896540
transform 1 0 6808 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _806_
timestamp 1704896540
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _807_
timestamp 1704896540
transform 1 0 8740 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _808_
timestamp 1704896540
transform -1 0 13432 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _809_
timestamp 1704896540
transform 1 0 10948 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _810_
timestamp 1704896540
transform 1 0 12696 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _811_
timestamp 1704896540
transform 1 0 11500 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _812_
timestamp 1704896540
transform 1 0 11040 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _813_
timestamp 1704896540
transform -1 0 12788 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _814_
timestamp 1704896540
transform 1 0 11592 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _815_
timestamp 1704896540
transform 1 0 25484 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _816_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 25208 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _817_
timestamp 1704896540
transform -1 0 22724 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _818_
timestamp 1704896540
transform 1 0 21252 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _819_
timestamp 1704896540
transform 1 0 24932 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _820_
timestamp 1704896540
transform -1 0 25300 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _821_
timestamp 1704896540
transform 1 0 21804 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _822_
timestamp 1704896540
transform 1 0 24012 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _823_
timestamp 1704896540
transform -1 0 26312 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _824_
timestamp 1704896540
transform 1 0 25484 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _825_
timestamp 1704896540
transform 1 0 24564 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _826_
timestamp 1704896540
transform 1 0 24288 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _827_
timestamp 1704896540
transform 1 0 23828 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _828_
timestamp 1704896540
transform 1 0 20240 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _829_
timestamp 1704896540
transform 1 0 18952 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _830_
timestamp 1704896540
transform -1 0 20148 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _831_
timestamp 1704896540
transform 1 0 12328 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _832_
timestamp 1704896540
transform 1 0 14168 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _833_
timestamp 1704896540
transform 1 0 12512 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _834_
timestamp 1704896540
transform 1 0 14260 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _835_
timestamp 1704896540
transform -1 0 17296 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _836_
timestamp 1704896540
transform -1 0 15640 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _837_
timestamp 1704896540
transform 1 0 12052 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _838_
timestamp 1704896540
transform 1 0 14536 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _839_
timestamp 1704896540
transform 1 0 17848 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _840_
timestamp 1704896540
transform -1 0 21068 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _841_
timestamp 1704896540
transform 1 0 20792 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _842_
timestamp 1704896540
transform -1 0 24196 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _843_
timestamp 1704896540
transform 1 0 19872 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _844_
timestamp 1704896540
transform 1 0 20056 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _845_
timestamp 1704896540
transform 1 0 21896 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _846_
timestamp 1704896540
transform -1 0 24840 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _847_
timestamp 1704896540
transform 1 0 23920 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _848_
timestamp 1704896540
transform 1 0 24196 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _849_
timestamp 1704896540
transform -1 0 25300 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _850_
timestamp 1704896540
transform -1 0 24840 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _851_
timestamp 1704896540
transform -1 0 22724 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _852_
timestamp 1704896540
transform -1 0 22724 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _853_
timestamp 1704896540
transform 1 0 18676 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _854_
timestamp 1704896540
transform 1 0 16192 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _855_
timestamp 1704896540
transform 1 0 6716 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _856_
timestamp 1704896540
transform 1 0 8372 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _857_
timestamp 1704896540
transform 1 0 7360 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _858_
timestamp 1704896540
transform 1 0 8188 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _859_
timestamp 1704896540
transform 1 0 8372 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _860_
timestamp 1704896540
transform 1 0 10948 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _861_
timestamp 1704896540
transform 1 0 9384 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _862_
timestamp 1704896540
transform 1 0 9936 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _863_
timestamp 1704896540
transform 1 0 14536 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _864_
timestamp 1704896540
transform 1 0 15732 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _865_
timestamp 1704896540
transform 1 0 14536 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _866_
timestamp 1704896540
transform 1 0 16652 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _867_
timestamp 1704896540
transform 1 0 16100 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _868_
timestamp 1704896540
transform 1 0 15640 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _869_
timestamp 1704896540
transform 1 0 16100 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _870_
timestamp 1704896540
transform 1 0 19136 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _871_
timestamp 1704896540
transform -1 0 19136 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _872_
timestamp 1704896540
transform 1 0 18492 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _873_
timestamp 1704896540
transform 1 0 18952 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _874_
timestamp 1704896540
transform 1 0 17112 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _875_
timestamp 1704896540
transform 1 0 18676 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _876_
timestamp 1704896540
transform 1 0 18676 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _877_
timestamp 1704896540
transform -1 0 21160 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _878_
timestamp 1704896540
transform -1 0 6440 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _879_
timestamp 1704896540
transform -1 0 7912 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _880_
timestamp 1704896540
transform -1 0 5336 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _881_
timestamp 1704896540
transform 1 0 5796 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _882_
timestamp 1704896540
transform 1 0 5796 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _883_
timestamp 1704896540
transform 1 0 7544 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _884_
timestamp 1704896540
transform 1 0 10212 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _885_
timestamp 1704896540
transform 1 0 10948 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _886_
timestamp 1704896540
transform 1 0 8004 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _887_
timestamp 1704896540
transform 1 0 3956 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _888_
timestamp 1704896540
transform 1 0 4232 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _889_
timestamp 1704896540
transform 1 0 2484 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _890_
timestamp 1704896540
transform 1 0 3220 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _891_
timestamp 1704896540
transform 1 0 2300 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _892_
timestamp 1704896540
transform 1 0 7544 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _893_
timestamp 1704896540
transform 1 0 11776 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _894_
timestamp 1704896540
transform -1 0 13432 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _895_
timestamp 1704896540
transform 1 0 8924 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _896_
timestamp 1704896540
transform -1 0 19596 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _897_
timestamp 1704896540
transform 1 0 16192 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _898_
timestamp 1704896540
transform 1 0 18676 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _899_
timestamp 1704896540
transform 1 0 19504 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _900_
timestamp 1704896540
transform 1 0 19780 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _901_
timestamp 1704896540
transform 1 0 19688 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _902_
timestamp 1704896540
transform 1 0 19136 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  _912_
timestamp 1704896540
transform -1 0 24564 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _913_
timestamp 1704896540
transform -1 0 10396 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _914_
timestamp 1704896540
transform -1 0 25116 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15824 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1704896540
transform -1 0 8188 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1704896540
transform 1 0 9844 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1704896540
transform -1 0 8280 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1704896540
transform 1 0 10948 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1704896540
transform -1 0 19504 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1704896540
transform 1 0 21068 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1704896540
transform 1 0 18676 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1704896540
transform 1 0 21528 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  digital_top_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4324 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_15
timestamp 1704896540
transform -1 0 3036 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_16
timestamp 1704896540
transform -1 0 2392 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_17
timestamp 1704896540
transform -1 0 9568 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_18
timestamp 1704896540
transform -1 0 8188 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_19
timestamp 1704896540
transform -1 0 7544 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_20
timestamp 1704896540
transform 1 0 5336 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_21
timestamp 1704896540
transform 1 0 4692 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_22
timestamp 1704896540
transform 1 0 3404 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1704896540
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1704896540
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1704896540
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_125 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12052 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_132 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12696 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1704896540
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1704896540
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_181 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17204 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_187
timestamp 1704896540
transform 1 0 17756 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_213
timestamp 1704896540
transform 1 0 20148 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1704896540
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_225
timestamp 1704896540
transform 1 0 21252 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_269
timestamp 1704896540
transform 1 0 25300 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1704896540
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_281
timestamp 1704896540
transform 1 0 26404 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8004 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1704896540
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_148
timestamp 1704896540
transform 1 0 14168 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_152
timestamp 1704896540
transform 1 0 14536 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_159
timestamp 1704896540
transform 1 0 15180 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_185
timestamp 1704896540
transform 1 0 17572 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_218
timestamp 1704896540
transform 1 0 20608 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_225
timestamp 1704896540
transform 1 0 21252 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_231
timestamp 1704896540
transform 1 0 21804 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_281
timestamp 1704896540
transform 1 0 26404 0 -1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1704896540
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8372 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_93
timestamp 1704896540
transform 1 0 9108 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_102 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9936 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_141
timestamp 1704896540
transform 1 0 13524 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_205
timestamp 1704896540
transform 1 0 19412 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_211
timestamp 1704896540
transform 1 0 19964 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_285
timestamp 1704896540
transform 1 0 26772 0 1 1632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_69
timestamp 1704896540
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_78
timestamp 1704896540
transform 1 0 7728 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_90
timestamp 1704896540
transform 1 0 8832 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_106
timestamp 1704896540
transform 1 0 10304 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 1704896540
transform 1 0 10948 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_148
timestamp 1704896540
transform 1 0 14168 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 1704896540
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_193
timestamp 1704896540
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_219
timestamp 1704896540
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1704896540
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_249
timestamp 1704896540
transform 1 0 23460 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_253
timestamp 1704896540
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_278
timestamp 1704896540
transform 1 0 26128 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5428 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_61
timestamp 1704896540
transform 1 0 6164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_88
timestamp 1704896540
transform 1 0 8648 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_94
timestamp 1704896540
transform 1 0 9200 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_106
timestamp 1704896540
transform 1 0 10304 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_114
timestamp 1704896540
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_121
timestamp 1704896540
transform 1 0 11684 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1704896540
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_165
timestamp 1704896540
transform 1 0 15732 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_173
timestamp 1704896540
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1704896540
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_205
timestamp 1704896540
transform 1 0 19412 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_209
timestamp 1704896540
transform 1 0 19780 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_234
timestamp 1704896540
transform 1 0 22080 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_248
timestamp 1704896540
transform 1 0 23368 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1704896540
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5244 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_65
timestamp 1704896540
transform 1 0 6532 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1704896540
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_113
timestamp 1704896540
transform 1 0 10948 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_142
timestamp 1704896540
transform 1 0 13616 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_193
timestamp 1704896540
transform 1 0 18308 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_202
timestamp 1704896540
transform 1 0 19136 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_206
timestamp 1704896540
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1704896540
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1704896540
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1704896540
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_281
timestamp 1704896540
transform 1 0 26404 0 -1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4324 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_60
timestamp 1704896540
transform 1 0 6072 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_90
timestamp 1704896540
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_108
timestamp 1704896540
transform 1 0 10488 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1704896540
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_163
timestamp 1704896540
transform 1 0 15548 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_191
timestamp 1704896540
transform 1 0 18124 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1704896540
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_197
timestamp 1704896540
transform 1 0 18676 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_216
timestamp 1704896540
transform 1 0 20424 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_236
timestamp 1704896540
transform 1 0 22264 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_249
timestamp 1704896540
transform 1 0 23460 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_269
timestamp 1704896540
transform 1 0 25300 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_281
timestamp 1704896540
transform 1 0 26404 0 1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1704896540
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_57
timestamp 1704896540
transform 1 0 5796 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_65
timestamp 1704896540
transform 1 0 6532 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_73
timestamp 1704896540
transform 1 0 7268 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8004 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_90
timestamp 1704896540
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_95
timestamp 1704896540
transform 1 0 9292 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_103
timestamp 1704896540
transform 1 0 10028 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1704896540
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_122
timestamp 1704896540
transform 1 0 11776 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_142
timestamp 1704896540
transform 1 0 13616 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_185
timestamp 1704896540
transform 1 0 17572 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 1704896540
transform 1 0 20976 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_265
timestamp 1704896540
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_277
timestamp 1704896540
transform 1 0 26036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_281
timestamp 1704896540
transform 1 0 26404 0 -1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_60
timestamp 1704896540
transform 1 0 6072 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_72
timestamp 1704896540
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1704896540
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_95
timestamp 1704896540
transform 1 0 9292 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_107
timestamp 1704896540
transform 1 0 10396 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_115
timestamp 1704896540
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1704896540
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1704896540
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_159
timestamp 1704896540
transform 1 0 15180 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_171
timestamp 1704896540
transform 1 0 16284 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_221
timestamp 1704896540
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1704896540
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1704896540
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4140 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_67
timestamp 1704896540
transform 1 0 6716 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_106
timestamp 1704896540
transform 1 0 10304 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_148
timestamp 1704896540
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_164
timestamp 1704896540
transform 1 0 15640 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_185
timestamp 1704896540
transform 1 0 17572 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_196
timestamp 1704896540
transform 1 0 18584 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1704896540
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_245
timestamp 1704896540
transform 1 0 23092 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_272
timestamp 1704896540
transform 1 0 25576 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_281
timestamp 1704896540
transform 1 0 26404 0 -1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4324 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_56
timestamp 1704896540
transform 1 0 5704 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_100
timestamp 1704896540
transform 1 0 9752 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_136
timestamp 1704896540
transform 1 0 13064 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_141
timestamp 1704896540
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_149
timestamp 1704896540
transform 1 0 14260 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_164
timestamp 1704896540
transform 1 0 15640 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_189
timestamp 1704896540
transform 1 0 17940 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_205
timestamp 1704896540
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_243
timestamp 1704896540
transform 1 0 22908 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1704896540
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1704896540
transform 1 0 26036 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1704896540
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_51
timestamp 1704896540
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_60
timestamp 1704896540
transform 1 0 6072 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_83
timestamp 1704896540
transform 1 0 8188 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_87
timestamp 1704896540
transform 1 0 8556 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_94
timestamp 1704896540
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1704896540
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_149
timestamp 1704896540
transform 1 0 14260 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_177
timestamp 1704896540
transform 1 0 16836 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_249
timestamp 1704896540
transform 1 0 23460 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_257
timestamp 1704896540
transform 1 0 24196 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1704896540
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3220 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_56
timestamp 1704896540
transform 1 0 5704 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_73
timestamp 1704896540
transform 1 0 7268 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1704896540
transform 1 0 8004 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8372 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_126
timestamp 1704896540
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_149
timestamp 1704896540
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_180
timestamp 1704896540
transform 1 0 17112 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_194
timestamp 1704896540
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_241
timestamp 1704896540
transform 1 0 22724 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_249
timestamp 1704896540
transform 1 0 23460 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_285
timestamp 1704896540
transform 1 0 26772 0 1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_39
timestamp 1704896540
transform 1 0 4140 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1704896540
transform 1 0 5428 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_72
timestamp 1704896540
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_84
timestamp 1704896540
transform 1 0 8280 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp 1704896540
transform 1 0 10948 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 1704896540
transform 1 0 15732 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_177
timestamp 1704896540
transform 1 0 16836 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_187
timestamp 1704896540
transform 1 0 17756 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_199
timestamp 1704896540
transform 1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_214
timestamp 1704896540
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_241
timestamp 1704896540
transform 1 0 22724 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_252
timestamp 1704896540
transform 1 0 23736 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1704896540
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_286
timestamp 1704896540
transform 1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_54
timestamp 1704896540
transform 1 0 5520 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_65
timestamp 1704896540
transform 1 0 6532 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_71
timestamp 1704896540
transform 1 0 7084 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_80
timestamp 1704896540
transform 1 0 7912 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_101
timestamp 1704896540
transform 1 0 9844 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_113
timestamp 1704896540
transform 1 0 10948 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_146
timestamp 1704896540
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_164
timestamp 1704896540
transform 1 0 15640 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_176
timestamp 1704896540
transform 1 0 16744 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_184
timestamp 1704896540
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1704896540
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_213
timestamp 1704896540
transform 1 0 20148 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_246
timestamp 1704896540
transform 1 0 23184 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_269
timestamp 1704896540
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_287
timestamp 1704896540
transform 1 0 26956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_3
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_9
timestamp 1704896540
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_26
timestamp 1704896540
transform 1 0 2944 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_38
timestamp 1704896540
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_57
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_66
timestamp 1704896540
transform 1 0 6624 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_74
timestamp 1704896540
transform 1 0 7360 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_104
timestamp 1704896540
transform 1 0 10120 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1704896540
transform 1 0 15732 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_196
timestamp 1704896540
transform 1 0 18584 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_204
timestamp 1704896540
transform 1 0 19320 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_219
timestamp 1704896540
transform 1 0 20700 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1704896540
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1704896540
transform 1 0 21252 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1704896540
transform 1 0 22356 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_249
timestamp 1704896540
transform 1 0 23460 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_257
timestamp 1704896540
transform 1 0 24196 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1704896540
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_3
timestamp 1704896540
transform 1 0 828 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_23
timestamp 1704896540
transform 1 0 2668 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_44
timestamp 1704896540
transform 1 0 4600 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_66
timestamp 1704896540
transform 1 0 6624 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_98
timestamp 1704896540
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_108
timestamp 1704896540
transform 1 0 10488 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_116
timestamp 1704896540
transform 1 0 11224 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_135
timestamp 1704896540
transform 1 0 12972 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1704896540
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_141
timestamp 1704896540
transform 1 0 13524 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_145
timestamp 1704896540
transform 1 0 13892 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_182
timestamp 1704896540
transform 1 0 17296 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_190
timestamp 1704896540
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_201
timestamp 1704896540
transform 1 0 19044 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_212
timestamp 1704896540
transform 1 0 20056 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_231
timestamp 1704896540
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_239
timestamp 1704896540
transform 1 0 22540 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_246
timestamp 1704896540
transform 1 0 23184 0 1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1704896540
transform 1 0 26036 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1704896540
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_15
timestamp 1704896540
transform 1 0 1932 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_19
timestamp 1704896540
transform 1 0 2300 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_44
timestamp 1704896540
transform 1 0 4600 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1704896540
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_62
timestamp 1704896540
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_90
timestamp 1704896540
transform 1 0 8832 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_104
timestamp 1704896540
transform 1 0 10120 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_113
timestamp 1704896540
transform 1 0 10948 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_146
timestamp 1704896540
transform 1 0 13984 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_158
timestamp 1704896540
transform 1 0 15088 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1704896540
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_169
timestamp 1704896540
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_177
timestamp 1704896540
transform 1 0 16836 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_184
timestamp 1704896540
transform 1 0 17480 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_188
timestamp 1704896540
transform 1 0 17848 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_196
timestamp 1704896540
transform 1 0 18584 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_216
timestamp 1704896540
transform 1 0 20424 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_252
timestamp 1704896540
transform 1 0 23736 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_258
timestamp 1704896540
transform 1 0 24288 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_270
timestamp 1704896540
transform 1 0 25392 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_278
timestamp 1704896540
transform 1 0 26128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_281
timestamp 1704896540
transform 1 0 26404 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 1704896540
transform 1 0 828 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_11
timestamp 1704896540
transform 1 0 1564 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_58
timestamp 1704896540
transform 1 0 5888 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_70
timestamp 1704896540
transform 1 0 6992 0 1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_101
timestamp 1704896540
transform 1 0 9844 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_113
timestamp 1704896540
transform 1 0 10948 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_141
timestamp 1704896540
transform 1 0 13524 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_147
timestamp 1704896540
transform 1 0 14076 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_164
timestamp 1704896540
transform 1 0 15640 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_170
timestamp 1704896540
transform 1 0 16192 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_179
timestamp 1704896540
transform 1 0 17020 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_191
timestamp 1704896540
transform 1 0 18124 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1704896540
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_218
timestamp 1704896540
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_248
timestamp 1704896540
transform 1 0 23368 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_265
timestamp 1704896540
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_276
timestamp 1704896540
transform 1 0 25944 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_288
timestamp 1704896540
transform 1 0 27048 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1704896540
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_27
timestamp 1704896540
transform 1 0 3036 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_31
timestamp 1704896540
transform 1 0 3404 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_39
timestamp 1704896540
transform 1 0 4140 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_62
timestamp 1704896540
transform 1 0 6256 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_66
timestamp 1704896540
transform 1 0 6624 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_93
timestamp 1704896540
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_103
timestamp 1704896540
transform 1 0 10028 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1704896540
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 1704896540
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_123
timestamp 1704896540
transform 1 0 11868 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_127
timestamp 1704896540
transform 1 0 12236 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_144
timestamp 1704896540
transform 1 0 13800 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_156
timestamp 1704896540
transform 1 0 14904 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_169
timestamp 1704896540
transform 1 0 16100 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_186
timestamp 1704896540
transform 1 0 17664 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_192
timestamp 1704896540
transform 1 0 18216 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_202
timestamp 1704896540
transform 1 0 19136 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_211
timestamp 1704896540
transform 1 0 19964 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1704896540
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_225
timestamp 1704896540
transform 1 0 21252 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_248
timestamp 1704896540
transform 1 0 23368 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_261
timestamp 1704896540
transform 1 0 24564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1704896540
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_281
timestamp 1704896540
transform 1 0 26404 0 -1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_15
timestamp 1704896540
transform 1 0 1932 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_23
timestamp 1704896540
transform 1 0 2668 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_69
timestamp 1704896540
transform 1 0 6900 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_80
timestamp 1704896540
transform 1 0 7912 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_107
timestamp 1704896540
transform 1 0 10396 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 1704896540
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_165
timestamp 1704896540
transform 1 0 15732 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_187
timestamp 1704896540
transform 1 0 17756 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 1704896540
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_217
timestamp 1704896540
transform 1 0 20516 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_249
timestamp 1704896540
transform 1 0 23460 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_253
timestamp 1704896540
transform 1 0 23828 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_281
timestamp 1704896540
transform 1 0 26404 0 1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1704896540
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_15
timestamp 1704896540
transform 1 0 1932 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1704896540
transform 1 0 5428 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_65
timestamp 1704896540
transform 1 0 6532 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_73
timestamp 1704896540
transform 1 0 7268 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 1704896540
transform 1 0 10396 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1704896540
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_147
timestamp 1704896540
transform 1 0 14076 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_164
timestamp 1704896540
transform 1 0 15640 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_183
timestamp 1704896540
transform 1 0 17388 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_198
timestamp 1704896540
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_203
timestamp 1704896540
transform 1 0 19228 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_219
timestamp 1704896540
transform 1 0 20700 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1704896540
transform 1 0 21068 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_239
timestamp 1704896540
transform 1 0 22540 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_245
timestamp 1704896540
transform 1 0 23092 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_274
timestamp 1704896540
transform 1 0 25760 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_281
timestamp 1704896540
transform 1 0 26404 0 -1 12512
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1704896540
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_15
timestamp 1704896540
transform 1 0 1932 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_23
timestamp 1704896540
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_39
timestamp 1704896540
transform 1 0 4140 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_47
timestamp 1704896540
transform 1 0 4876 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_88
timestamp 1704896540
transform 1 0 8648 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_96
timestamp 1704896540
transform 1 0 9384 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_109
timestamp 1704896540
transform 1 0 10580 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_121
timestamp 1704896540
transform 1 0 11684 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_138
timestamp 1704896540
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1704896540
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_156
timestamp 1704896540
transform 1 0 14904 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_164
timestamp 1704896540
transform 1 0 15640 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_193
timestamp 1704896540
transform 1 0 18308 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_218
timestamp 1704896540
transform 1 0 20608 0 1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_236
timestamp 1704896540
transform 1 0 22264 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_248
timestamp 1704896540
transform 1 0 23368 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_253
timestamp 1704896540
transform 1 0 23828 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_287
timestamp 1704896540
transform 1 0 26956 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1704896540
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1704896540
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1704896540
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1704896540
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_65
timestamp 1704896540
transform 1 0 6532 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_73
timestamp 1704896540
transform 1 0 7268 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_100
timestamp 1704896540
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_145
timestamp 1704896540
transform 1 0 13892 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_151
timestamp 1704896540
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1704896540
transform 1 0 15364 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1704896540
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_181
timestamp 1704896540
transform 1 0 17204 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_190
timestamp 1704896540
transform 1 0 18032 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_202
timestamp 1704896540
transform 1 0 19136 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_214
timestamp 1704896540
transform 1 0 20240 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1704896540
transform 1 0 20976 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_239
timestamp 1704896540
transform 1 0 22540 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_251
timestamp 1704896540
transform 1 0 23644 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_259
timestamp 1704896540
transform 1 0 24380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_276
timestamp 1704896540
transform 1 0 25944 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_281
timestamp 1704896540
transform 1 0 26404 0 -1 13600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1704896540
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_15
timestamp 1704896540
transform 1 0 1932 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_23
timestamp 1704896540
transform 1 0 2668 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1704896540
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_29
timestamp 1704896540
transform 1 0 3220 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_35
timestamp 1704896540
transform 1 0 3772 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_60
timestamp 1704896540
transform 1 0 6072 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_72
timestamp 1704896540
transform 1 0 7176 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_78
timestamp 1704896540
transform 1 0 7728 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_108
timestamp 1704896540
transform 1 0 10488 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1704896540
transform 1 0 12788 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1704896540
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_141
timestamp 1704896540
transform 1 0 13524 0 1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_163
timestamp 1704896540
transform 1 0 15548 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_175
timestamp 1704896540
transform 1 0 16652 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_192
timestamp 1704896540
transform 1 0 18216 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_202
timestamp 1704896540
transform 1 0 19136 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_207
timestamp 1704896540
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_239
timestamp 1704896540
transform 1 0 22540 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1704896540
transform 1 0 23644 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_276
timestamp 1704896540
transform 1 0 25944 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_288
timestamp 1704896540
transform 1 0 27048 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1704896540
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_15
timestamp 1704896540
transform 1 0 1932 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_40
timestamp 1704896540
transform 1 0 4232 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_48
timestamp 1704896540
transform 1 0 4968 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_73
timestamp 1704896540
transform 1 0 7268 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_92
timestamp 1704896540
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_101
timestamp 1704896540
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1704896540
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1704896540
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_125
timestamp 1704896540
transform 1 0 12052 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_146
timestamp 1704896540
transform 1 0 13984 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1704896540
transform 1 0 15364 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1704896540
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16100 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_177
timestamp 1704896540
transform 1 0 16836 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_183
timestamp 1704896540
transform 1 0 17388 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_196
timestamp 1704896540
transform 1 0 18584 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_205
timestamp 1704896540
transform 1 0 19412 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_222
timestamp 1704896540
transform 1 0 20976 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_225
timestamp 1704896540
transform 1 0 21252 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_248
timestamp 1704896540
transform 1 0 23368 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_262
timestamp 1704896540
transform 1 0 24656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_281
timestamp 1704896540
transform 1 0 26404 0 -1 14688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1704896540
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1704896540
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1704896540
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_41
timestamp 1704896540
transform 1 0 4324 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1704896540
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1704896540
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1704896540
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_108
timestamp 1704896540
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_118
timestamp 1704896540
transform 1 0 11408 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_124
timestamp 1704896540
transform 1 0 11960 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_130
timestamp 1704896540
transform 1 0 12512 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_150
timestamp 1704896540
transform 1 0 14352 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_154
timestamp 1704896540
transform 1 0 14720 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_159
timestamp 1704896540
transform 1 0 15180 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_167
timestamp 1704896540
transform 1 0 15916 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_175
timestamp 1704896540
transform 1 0 16652 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_179
timestamp 1704896540
transform 1 0 17020 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_213
timestamp 1704896540
transform 1 0 20148 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_225
timestamp 1704896540
transform 1 0 21252 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_237
timestamp 1704896540
transform 1 0 22356 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_249
timestamp 1704896540
transform 1 0 23460 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_253
timestamp 1704896540
transform 1 0 23828 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_274
timestamp 1704896540
transform 1 0 25760 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_286
timestamp 1704896540
transform 1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1704896540
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1704896540
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_27
timestamp 1704896540
transform 1 0 3036 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_35
timestamp 1704896540
transform 1 0 3772 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_39
timestamp 1704896540
transform 1 0 4140 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_54
timestamp 1704896540
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1704896540
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_93
timestamp 1704896540
transform 1 0 9108 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_104
timestamp 1704896540
transform 1 0 10120 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_113
timestamp 1704896540
transform 1 0 10948 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_133
timestamp 1704896540
transform 1 0 12788 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_146
timestamp 1704896540
transform 1 0 13984 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_150
timestamp 1704896540
transform 1 0 14352 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1704896540
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_175
timestamp 1704896540
transform 1 0 16652 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_180
timestamp 1704896540
transform 1 0 17112 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_186
timestamp 1704896540
transform 1 0 17664 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_191
timestamp 1704896540
transform 1 0 18124 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_199
timestamp 1704896540
transform 1 0 18860 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_225
timestamp 1704896540
transform 1 0 21252 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_271
timestamp 1704896540
transform 1 0 25484 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1704896540
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_281
timestamp 1704896540
transform 1 0 26404 0 -1 15776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1704896540
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_15
timestamp 1704896540
transform 1 0 1932 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_23
timestamp 1704896540
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_45
timestamp 1704896540
transform 1 0 4692 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_80
timestamp 1704896540
transform 1 0 7912 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_85
timestamp 1704896540
transform 1 0 8372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_94
timestamp 1704896540
transform 1 0 9200 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_102
timestamp 1704896540
transform 1 0 9936 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_137
timestamp 1704896540
transform 1 0 13156 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_141
timestamp 1704896540
transform 1 0 13524 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_163
timestamp 1704896540
transform 1 0 15548 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_172
timestamp 1704896540
transform 1 0 16376 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_180
timestamp 1704896540
transform 1 0 17112 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_197
timestamp 1704896540
transform 1 0 18676 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_205
timestamp 1704896540
transform 1 0 19412 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_218
timestamp 1704896540
transform 1 0 20608 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_230
timestamp 1704896540
transform 1 0 21712 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_238
timestamp 1704896540
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_246
timestamp 1704896540
transform 1 0 23184 0 1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_256
timestamp 1704896540
transform 1 0 24104 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_268
timestamp 1704896540
transform 1 0 25208 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_280
timestamp 1704896540
transform 1 0 26312 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_288
timestamp 1704896540
transform 1 0 27048 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1704896540
transform 1 0 828 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_15
timestamp 1704896540
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_20
timestamp 1704896540
transform 1 0 2392 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_32
timestamp 1704896540
transform 1 0 3496 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_60
timestamp 1704896540
transform 1 0 6072 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_78
timestamp 1704896540
transform 1 0 7728 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_110
timestamp 1704896540
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_113
timestamp 1704896540
transform 1 0 10948 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_138
timestamp 1704896540
transform 1 0 13248 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_147
timestamp 1704896540
transform 1 0 14076 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_152
timestamp 1704896540
transform 1 0 14536 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_207
timestamp 1704896540
transform 1 0 19596 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_267
timestamp 1704896540
transform 1 0 25116 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1704896540
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_281
timestamp 1704896540
transform 1 0 26404 0 -1 16864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1704896540
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_15
timestamp 1704896540
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_20
timestamp 1704896540
transform 1 0 2392 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1704896540
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_29
timestamp 1704896540
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_34
timestamp 1704896540
transform 1 0 3680 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_41
timestamp 1704896540
transform 1 0 4324 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_48
timestamp 1704896540
transform 1 0 4968 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_55
timestamp 1704896540
transform 1 0 5612 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_57
timestamp 1704896540
transform 1 0 5796 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_69
timestamp 1704896540
transform 1 0 6900 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_76
timestamp 1704896540
transform 1 0 7544 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1704896540
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_85
timestamp 1704896540
transform 1 0 8372 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_98
timestamp 1704896540
transform 1 0 9568 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_102
timestamp 1704896540
transform 1 0 9936 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_107
timestamp 1704896540
transform 1 0 10396 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_111
timestamp 1704896540
transform 1 0 10764 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_113
timestamp 1704896540
transform 1 0 10948 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_121
timestamp 1704896540
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_126
timestamp 1704896540
transform 1 0 12144 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_131
timestamp 1704896540
transform 1 0 12604 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_136
timestamp 1704896540
transform 1 0 13064 0 1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1704896540
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_153
timestamp 1704896540
transform 1 0 14628 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_157
timestamp 1704896540
transform 1 0 14996 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_167
timestamp 1704896540
transform 1 0 15916 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_169
timestamp 1704896540
transform 1 0 16100 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_173
timestamp 1704896540
transform 1 0 16468 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_177
timestamp 1704896540
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_189
timestamp 1704896540
transform 1 0 17940 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_197
timestamp 1704896540
transform 1 0 18676 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_205
timestamp 1704896540
transform 1 0 19412 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1704896540
transform 1 0 19780 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_221
timestamp 1704896540
transform 1 0 20884 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_225
timestamp 1704896540
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_230
timestamp 1704896540
transform 1 0 21712 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_237
timestamp 1704896540
transform 1 0 22356 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 1704896540
transform 1 0 23552 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_259
timestamp 1704896540
transform 1 0 24380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_265
timestamp 1704896540
transform 1 0 24932 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_272
timestamp 1704896540
transform 1 0 25576 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_279
timestamp 1704896540
transform 1 0 26220 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_281
timestamp 1704896540
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_287
timestamp 1704896540
transform 1 0 26956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3772 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 12512 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform -1 0 13064 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform 1 0 22724 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 21988 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform -1 0 9384 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform -1 0 23736 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704896540
transform -1 0 23000 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1704896540
transform 1 0 4784 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1704896540
transform -1 0 12788 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1704896540
transform 1 0 21620 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1704896540
transform -1 0 23460 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1704896540
transform -1 0 20792 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1704896540
transform 1 0 17112 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1704896540
transform -1 0 6532 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1704896540
transform -1 0 22080 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1704896540
transform -1 0 21068 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1704896540
transform 1 0 20332 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1704896540
transform -1 0 21804 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1704896540
transform -1 0 16836 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1704896540
transform -1 0 15732 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1704896540
transform -1 0 25576 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1704896540
transform -1 0 24564 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1704896540
transform -1 0 16836 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1704896540
transform -1 0 15640 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1704896540
transform -1 0 19872 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1704896540
transform -1 0 22448 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1704896540
transform -1 0 23184 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1704896540
transform -1 0 10856 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1704896540
transform -1 0 20884 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1704896540
transform -1 0 20056 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1704896540
transform -1 0 6440 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1704896540
transform -1 0 6532 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1704896540
transform 1 0 25392 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1704896540
transform -1 0 27140 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1704896540
transform -1 0 24564 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1704896540
transform -1 0 25576 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1704896540
transform 1 0 6992 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1704896540
transform -1 0 17940 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1704896540
transform -1 0 16836 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1704896540
transform -1 0 24932 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1704896540
transform -1 0 26036 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1704896540
transform -1 0 24932 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1704896540
transform -1 0 14260 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1704896540
transform 1 0 24564 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1704896540
transform -1 0 26312 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1704896540
transform 1 0 9016 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1704896540
transform 1 0 6440 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1704896540
transform -1 0 7176 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1704896540
transform -1 0 23368 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1704896540
transform -1 0 25300 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1704896540
transform -1 0 12144 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1704896540
transform 1 0 9200 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1704896540
transform -1 0 22264 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1704896540
transform -1 0 26036 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1704896540
transform -1 0 25300 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1704896540
transform -1 0 20332 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1704896540
transform -1 0 20700 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1704896540
transform 1 0 18676 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1704896540
transform -1 0 20332 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1704896540
transform -1 0 13708 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1704896540
transform -1 0 11868 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1704896540
transform -1 0 25116 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1704896540
transform -1 0 17388 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1704896540
transform -1 0 18124 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1704896540
transform -1 0 18308 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1704896540
transform 1 0 17848 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1704896540
transform 1 0 18676 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1704896540
transform -1 0 16836 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1704896540
transform -1 0 20240 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1704896540
transform 1 0 16376 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1704896540
transform -1 0 13064 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1704896540
transform -1 0 17848 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1704896540
transform -1 0 16836 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1704896540
transform 1 0 8740 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1704896540
transform -1 0 8096 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1704896540
transform -1 0 18308 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1704896540
transform -1 0 13340 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1704896540
transform -1 0 25760 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1704896540
transform 1 0 4692 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1704896540
transform -1 0 3956 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1704896540
transform -1 0 2668 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1704896540
transform -1 0 5428 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1704896540
transform -1 0 27140 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1704896540
transform -1 0 9016 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1704896540
transform -1 0 4324 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1704896540
transform -1 0 27140 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1704896540
transform -1 0 26772 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1704896540
transform 1 0 12236 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1704896540
transform -1 0 18124 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1704896540
transform 1 0 9752 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1704896540
transform -1 0 10028 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1704896540
transform 1 0 8924 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1704896540
transform 1 0 7544 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1704896540
transform 1 0 8372 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1704896540
transform -1 0 26036 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1704896540
transform 1 0 4600 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1704896540
transform -1 0 6532 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1704896540
transform -1 0 24012 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1704896540
transform 1 0 12788 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1704896540
transform 1 0 24380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1704896540
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1704896540
transform -1 0 11960 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1704896540
transform -1 0 13800 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1704896540
transform 1 0 10120 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1704896540
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1704896540
transform -1 0 26956 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 26220 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1704896540
transform 1 0 25300 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform 1 0 24656 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1704896540
transform 1 0 24104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1704896540
transform 1 0 23828 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1704896540
transform 1 0 23276 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1704896540
transform 1 0 22080 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1704896540
transform 1 0 21436 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1704896540
transform 1 0 19504 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1704896540
transform 1 0 18216 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1704896540
transform -1 0 17940 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1704896540
transform -1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_31
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 27416 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_32
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 27416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_33
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 27416 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_34
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 27416 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_35
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 27416 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_36
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 27416 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_37
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 27416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_38
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 27416 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_39
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 27416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_40
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 27416 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_41
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 27416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_42
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 27416 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_43
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 27416 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_44
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 27416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_45
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 27416 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_46
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 27416 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_47
timestamp 1704896540
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 27416 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_48
timestamp 1704896540
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 27416 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_49
timestamp 1704896540
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 27416 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_50
timestamp 1704896540
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 27416 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_51
timestamp 1704896540
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 27416 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_52
timestamp 1704896540
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 27416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_53
timestamp 1704896540
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 27416 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_54
timestamp 1704896540
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 27416 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_55
timestamp 1704896540
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 27416 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_56
timestamp 1704896540
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 27416 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_57
timestamp 1704896540
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 27416 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_58
timestamp 1704896540
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 27416 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_59
timestamp 1704896540
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 27416 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_60
timestamp 1704896540
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 27416 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_61
timestamp 1704896540
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 27416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp 1704896540
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp 1704896540
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp 1704896540
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68
timestamp 1704896540
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1704896540
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1704896540
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1704896540
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_72
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_73
timestamp 1704896540
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_74
timestamp 1704896540
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_75
timestamp 1704896540
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_76
timestamp 1704896540
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_77
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_78
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_79
timestamp 1704896540
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_80
timestamp 1704896540
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_81
timestamp 1704896540
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_82
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_83
timestamp 1704896540
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_84
timestamp 1704896540
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_85
timestamp 1704896540
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_86
timestamp 1704896540
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_87
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_88
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_89
timestamp 1704896540
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_90
timestamp 1704896540
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_91
timestamp 1704896540
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_92
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_93
timestamp 1704896540
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_94
timestamp 1704896540
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_95
timestamp 1704896540
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_96
timestamp 1704896540
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_97
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_98
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_99
timestamp 1704896540
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_100
timestamp 1704896540
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_101
timestamp 1704896540
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_102
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_103
timestamp 1704896540
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_104
timestamp 1704896540
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_105
timestamp 1704896540
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_106
timestamp 1704896540
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_107
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_108
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_109
timestamp 1704896540
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_110
timestamp 1704896540
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_111
timestamp 1704896540
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_112
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_113
timestamp 1704896540
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_114
timestamp 1704896540
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_115
timestamp 1704896540
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_116
timestamp 1704896540
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_117
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_118
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_119
timestamp 1704896540
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_120
timestamp 1704896540
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_121
timestamp 1704896540
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_122
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_123
timestamp 1704896540
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_124
timestamp 1704896540
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_125
timestamp 1704896540
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_126
timestamp 1704896540
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_127
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_128
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_129
timestamp 1704896540
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_130
timestamp 1704896540
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_131
timestamp 1704896540
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_132
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_133
timestamp 1704896540
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_134
timestamp 1704896540
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_135
timestamp 1704896540
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_136
timestamp 1704896540
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_137
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_138
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_139
timestamp 1704896540
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_140
timestamp 1704896540
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_141
timestamp 1704896540
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_142
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_143
timestamp 1704896540
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_144
timestamp 1704896540
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_145
timestamp 1704896540
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_146
timestamp 1704896540
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_147
timestamp 1704896540
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_148
timestamp 1704896540
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_149
timestamp 1704896540
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_150
timestamp 1704896540
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_151
timestamp 1704896540
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_152
timestamp 1704896540
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_153
timestamp 1704896540
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_154
timestamp 1704896540
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_155
timestamp 1704896540
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_156
timestamp 1704896540
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_157
timestamp 1704896540
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_158
timestamp 1704896540
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_159
timestamp 1704896540
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_160
timestamp 1704896540
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp 1704896540
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_162
timestamp 1704896540
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_163
timestamp 1704896540
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp 1704896540
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp 1704896540
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_166
timestamp 1704896540
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_167
timestamp 1704896540
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp 1704896540
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp 1704896540
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_170
timestamp 1704896540
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_171
timestamp 1704896540
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_172
timestamp 1704896540
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_173
timestamp 1704896540
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_174
timestamp 1704896540
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_175
timestamp 1704896540
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_176
timestamp 1704896540
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_177
timestamp 1704896540
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_178
timestamp 1704896540
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_179
timestamp 1704896540
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_180
timestamp 1704896540
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_181
timestamp 1704896540
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_182
timestamp 1704896540
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_183
timestamp 1704896540
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_184
timestamp 1704896540
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_185
timestamp 1704896540
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_186
timestamp 1704896540
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_187
timestamp 1704896540
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_188
timestamp 1704896540
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_189
timestamp 1704896540
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_190
timestamp 1704896540
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_191
timestamp 1704896540
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_192
timestamp 1704896540
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_193
timestamp 1704896540
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_194
timestamp 1704896540
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_195
timestamp 1704896540
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_196
timestamp 1704896540
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_197
timestamp 1704896540
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_198
timestamp 1704896540
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_199
timestamp 1704896540
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_200
timestamp 1704896540
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_201
timestamp 1704896540
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_202
timestamp 1704896540
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_203
timestamp 1704896540
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_204
timestamp 1704896540
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_205
timestamp 1704896540
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_206
timestamp 1704896540
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_207
timestamp 1704896540
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_208
timestamp 1704896540
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_209
timestamp 1704896540
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_210
timestamp 1704896540
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_211
timestamp 1704896540
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_212
timestamp 1704896540
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_213
timestamp 1704896540
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_214
timestamp 1704896540
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_215
timestamp 1704896540
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_216
timestamp 1704896540
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_217
timestamp 1704896540
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_218
timestamp 1704896540
transform 1 0 5704 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_219
timestamp 1704896540
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_220
timestamp 1704896540
transform 1 0 10856 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_221
timestamp 1704896540
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_222
timestamp 1704896540
transform 1 0 16008 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_223
timestamp 1704896540
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_224
timestamp 1704896540
transform 1 0 21160 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_225
timestamp 1704896540
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_226
timestamp 1704896540
transform 1 0 26312 0 1 16864
box -38 -48 130 592
<< labels >>
rlabel metal2 s 14064 16864 14064 16864 4 VGND
rlabel metal1 s 13984 17408 13984 17408 4 VPWR
rlabel metal2 s 25801 12750 25801 12750 4 _000_
rlabel metal2 s 24518 11798 24518 11798 4 _001_
rlabel metal2 s 22218 11186 22218 11186 4 _002_
rlabel metal1 s 21666 9690 21666 9690 4 _003_
rlabel metal2 s 25346 11458 25346 11458 4 _004_
rlabel metal1 s 3440 10574 3440 10574 4 _005_
rlabel metal1 s 2484 10234 2484 10234 4 _006_
rlabel metal1 s 2392 9554 2392 9554 4 _007_
rlabel metal2 s 5290 8636 5290 8636 4 _008_
rlabel metal1 s 2893 7990 2893 7990 4 _009_
rlabel metal1 s 4135 7242 4135 7242 4 _010_
rlabel metal2 s 5934 7106 5934 7106 4 _011_
rlabel metal2 s 5386 5746 5386 5746 4 _012_
rlabel metal2 s 8597 5746 8597 5746 4 _013_
rlabel metal2 s 7590 4964 7590 4964 4 _014_
rlabel metal1 s 5377 5134 5377 5134 4 _015_
rlabel metal2 s 4917 3978 4917 3978 4 _016_
rlabel metal2 s 9333 4046 9333 4046 4 _017_
rlabel metal2 s 6394 3604 6394 3604 4 _018_
rlabel metal1 s 7355 2890 7355 2890 4 _019_
rlabel metal1 s 9149 1462 9149 1462 4 _020_
rlabel metal1 s 13396 1870 13396 1870 4 _021_
rlabel metal1 s 11265 1394 11265 1394 4 _022_
rlabel metal1 s 12742 986 12742 986 4 _023_
rlabel metal1 s 13018 3536 13018 3536 4 _024_
rlabel metal1 s 11254 3978 11254 3978 4 _025_
rlabel metal2 s 12466 5882 12466 5882 4 _026_
rlabel metal1 s 11812 5746 11812 5746 4 _027_
rlabel metal1 s 24610 13498 24610 13498 4 _028_
rlabel metal2 s 22126 15062 22126 15062 4 _029_
rlabel metal2 s 24794 15334 24794 15334 4 _030_
rlabel metal2 s 25530 14246 25530 14246 4 _031_
rlabel metal2 s 25801 8398 25801 8398 4 _032_
rlabel metal1 s 25295 6222 25295 6222 4 _033_
rlabel metal2 s 24605 6902 24605 6902 4 _034_
rlabel metal2 s 23690 8194 23690 8194 4 _035_
rlabel metal1 s 20603 8330 20603 8330 4 _036_
rlabel metal2 s 19269 10166 19269 10166 4 _037_
rlabel metal1 s 19928 10574 19928 10574 4 _038_
rlabel metal2 s 12650 10982 12650 10982 4 _039_
rlabel metal1 s 13922 10506 13922 10506 4 _040_
rlabel metal1 s 12732 10098 12732 10098 4 _041_
rlabel metal1 s 14382 9078 14382 9078 4 _042_
rlabel metal2 s 16882 9282 16882 9282 4 _043_
rlabel metal1 s 14862 8398 14862 8398 4 _044_
rlabel metal2 s 12834 7038 12834 7038 4 _045_
rlabel metal1 s 15272 7854 15272 7854 4 _046_
rlabel metal1 s 18216 6426 18216 6426 4 _047_
rlabel metal1 s 21252 5338 21252 5338 4 _048_
rlabel metal1 s 21988 4590 21988 4590 4 _049_
rlabel metal1 s 23920 3706 23920 3706 4 _050_
rlabel metal1 s 21160 3502 21160 3502 4 _051_
rlabel metal1 s 22540 986 22540 986 4 _052_
rlabel metal1 s 24058 850 24058 850 4 _053_
rlabel metal1 s 26496 1394 26496 1394 4 _054_
rlabel metal2 s 25990 2244 25990 2244 4 _055_
rlabel metal1 s 24840 3026 24840 3026 4 _056_
rlabel metal1 s 25024 4794 25024 4794 4 _057_
rlabel metal1 s 24518 5338 24518 5338 4 _058_
rlabel metal1 s 22908 6426 22908 6426 4 _059_
rlabel metal2 s 23046 8228 23046 8228 4 _060_
rlabel metal1 s 18706 8330 18706 8330 4 _061_
rlabel metal1 s 16422 10778 16422 10778 4 _062_
rlabel metal2 s 7033 11254 7033 11254 4 _063_
rlabel metal1 s 8448 10506 8448 10506 4 _064_
rlabel metal1 s 7544 9486 7544 9486 4 _065_
rlabel metal2 s 8505 9010 8505 9010 4 _066_
rlabel metal1 s 8402 8330 8402 8330 4 _067_
rlabel metal2 s 11270 8806 11270 8806 4 _068_
rlabel metal1 s 9885 6834 9885 6834 4 _069_
rlabel metal1 s 9200 7378 9200 7378 4 _070_
rlabel metal2 s 14950 6052 14950 6052 4 _071_
rlabel metal1 s 16836 5678 16836 5678 4 _072_
rlabel metal2 s 14858 4454 14858 4454 4 _073_
rlabel metal1 s 18078 3570 18078 3570 4 _074_
rlabel metal1 s 16320 3570 16320 3570 4 _075_
rlabel metal2 s 16698 2244 16698 2244 4 _076_
rlabel metal2 s 16882 1870 16882 1870 4 _077_
rlabel metal1 s 19964 986 19964 986 4 _078_
rlabel metal2 s 18722 1292 18722 1292 4 _079_
rlabel metal1 s 18630 2074 18630 2074 4 _080_
rlabel metal2 s 19090 3842 19090 3842 4 _081_
rlabel metal2 s 16882 4862 16882 4862 4 _082_
rlabel metal2 s 18993 5066 18993 5066 4 _083_
rlabel metal2 s 19918 7004 19918 7004 4 _084_
rlabel metal1 s 20608 16218 20608 16218 4 _085_
rlabel metal1 s 5984 12682 5984 12682 4 _086_
rlabel metal1 s 7406 15674 7406 15674 4 _087_
rlabel metal1 s 5213 13770 5213 13770 4 _088_
rlabel metal1 s 6016 15538 6016 15538 4 _089_
rlabel metal1 s 6016 14450 6016 14450 4 _090_
rlabel metal2 s 8418 14212 8418 14212 4 _091_
rlabel metal1 s 10534 15130 10534 15130 4 _092_
rlabel metal1 s 11040 12954 11040 12954 4 _093_
rlabel metal2 s 8694 16422 8694 16422 4 _094_
rlabel metal1 s 3634 11866 3634 11866 4 _095_
rlabel metal1 s 5193 16626 5193 16626 4 _096_
rlabel metal1 s 2852 12614 2852 12614 4 _097_
rlabel metal1 s 3296 15946 3296 15946 4 _098_
rlabel metal2 s 2622 14246 2622 14246 4 _099_
rlabel metal2 s 8418 13158 8418 13158 4 _100_
rlabel metal1 s 11990 16694 11990 16694 4 _101_
rlabel metal1 s 13340 12614 13340 12614 4 _102_
rlabel metal1 s 9052 12274 9052 12274 4 _103_
rlabel metal2 s 18538 16422 18538 16422 4 _104_
rlabel metal1 s 16488 12682 16488 12682 4 _105_
rlabel metal1 s 18942 14858 18942 14858 4 _106_
rlabel metal1 s 19770 14518 19770 14518 4 _107_
rlabel metal1 s 20000 13838 20000 13838 4 _108_
rlabel metal1 s 19810 15606 19810 15606 4 _109_
rlabel metal2 s 19453 12682 19453 12682 4 _110_
rlabel metal2 s 15686 15232 15686 15232 4 _111_
rlabel metal2 s 11822 14688 11822 14688 4 _112_
rlabel metal1 s 15962 5100 15962 5100 4 _113_
rlabel metal2 s 10396 1972 10396 1972 4 _114_
rlabel metal1 s 25576 13498 25576 13498 4 _115_
rlabel metal1 s 25162 13328 25162 13328 4 _116_
rlabel metal1 s 17526 11628 17526 11628 4 _117_
rlabel metal1 s 25208 13430 25208 13430 4 _118_
rlabel metal2 s 23966 14654 23966 14654 4 _119_
rlabel metal1 s 25622 7752 25622 7752 4 _120_
rlabel metal1 s 22954 9452 22954 9452 4 _121_
rlabel metal1 s 23828 12886 23828 12886 4 _122_
rlabel metal1 s 25438 11118 25438 11118 4 _123_
rlabel metal1 s 25484 10982 25484 10982 4 _124_
rlabel metal1 s 21528 9486 21528 9486 4 _125_
rlabel metal2 s 22862 10030 22862 10030 4 _126_
rlabel metal1 s 17572 10166 17572 10166 4 _127_
rlabel metal1 s 19734 816 19734 816 4 _128_
rlabel metal1 s 16238 8806 16238 8806 4 _129_
rlabel metal2 s 21850 5763 21850 5763 4 _130_
rlabel metal1 s 11594 10098 11594 10098 4 _131_
rlabel metal1 s 23084 11526 23084 11526 4 _132_
rlabel metal1 s 22678 10575 22678 10575 4 _133_
rlabel metal2 s 23644 12580 23644 12580 4 _134_
rlabel metal1 s 2346 16660 2346 16660 4 _135_
rlabel metal1 s 2162 16694 2162 16694 4 _136_
rlabel metal1 s 14214 16728 14214 16728 4 _137_
rlabel metal1 s 21712 13362 21712 13362 4 _138_
rlabel metal1 s 19458 15946 19458 15946 4 _139_
rlabel metal1 s 14490 12614 14490 12614 4 _140_
rlabel metal1 s 16882 12172 16882 12172 4 _141_
rlabel metal1 s 18400 12274 18400 12274 4 _142_
rlabel metal1 s 20286 12274 20286 12274 4 _143_
rlabel metal1 s 21758 13260 21758 13260 4 _144_
rlabel metal2 s 21482 12070 21482 12070 4 _145_
rlabel metal2 s 21942 15266 21942 15266 4 _146_
rlabel metal1 s 12926 12206 12926 12206 4 _147_
rlabel metal1 s 19044 15878 19044 15878 4 _148_
rlabel metal1 s 14398 13498 14398 13498 4 _149_
rlabel metal1 s 14950 13974 14950 13974 4 _150_
rlabel metal1 s 15180 16762 15180 16762 4 _151_
rlabel metal1 s 14628 16626 14628 16626 4 _152_
rlabel metal2 s 14766 14212 14766 14212 4 _153_
rlabel metal1 s 14398 14586 14398 14586 4 _154_
rlabel metal2 s 14490 15776 14490 15776 4 _155_
rlabel metal2 s 13938 16422 13938 16422 4 _156_
rlabel metal1 s 13340 14790 13340 14790 4 _157_
rlabel metal1 s 12696 15130 12696 15130 4 _158_
rlabel metal1 s 13018 14586 13018 14586 4 _159_
rlabel metal2 s 12374 15844 12374 15844 4 _160_
rlabel metal2 s 13202 15776 13202 15776 4 _161_
rlabel metal1 s 12052 16218 12052 16218 4 _162_
rlabel metal1 s 12788 13498 12788 13498 4 _163_
rlabel metal1 s 12834 13906 12834 13906 4 _164_
rlabel metal1 s 11684 14042 11684 14042 4 _165_
rlabel metal1 s 6532 16626 6532 16626 4 _166_
rlabel metal2 s 18078 12665 18078 12665 4 _167_
rlabel metal1 s 4416 13362 4416 13362 4 _168_
rlabel metal1 s 3036 9962 3036 9962 4 _169_
rlabel metal1 s 19044 9350 19044 9350 4 _170_
rlabel metal2 s 4278 10710 4278 10710 4 _171_
rlabel metal1 s 5106 9452 5106 9452 4 _172_
rlabel metal1 s 20516 16014 20516 16014 4 _173_
rlabel metal2 s 2898 9894 2898 9894 4 _174_
rlabel metal2 s 2070 9894 2070 9894 4 _175_
rlabel metal1 s 2254 10132 2254 10132 4 _176_
rlabel metal1 s 4876 8534 4876 8534 4 _177_
rlabel metal2 s 5014 8840 5014 8840 4 _178_
rlabel metal1 s 5336 8398 5336 8398 4 _179_
rlabel metal1 s 4462 7786 4462 7786 4 _180_
rlabel metal2 s 3450 8092 3450 8092 4 _181_
rlabel metal1 s 4830 8058 4830 8058 4 _182_
rlabel metal1 s 4830 7514 4830 7514 4 _183_
rlabel metal2 s 6026 7276 6026 7276 4 _184_
rlabel metal2 s 5842 7004 5842 7004 4 _185_
rlabel metal2 s 7130 6596 7130 6596 4 _186_
rlabel metal2 s 5566 6630 5566 6630 4 _187_
rlabel metal2 s 18262 14960 18262 14960 4 _188_
rlabel metal1 s 8510 5338 8510 5338 4 _189_
rlabel metal2 s 7820 4658 7820 4658 4 _190_
rlabel metal1 s 8740 5338 8740 5338 4 _191_
rlabel metal1 s 7774 4624 7774 4624 4 _192_
rlabel metal1 s 7682 4590 7682 4590 4 _193_
rlabel metal2 s 7590 3774 7590 3774 4 _194_
rlabel metal1 s 6670 6120 6670 6120 4 _195_
rlabel metal1 s 6072 5746 6072 5746 4 _196_
rlabel metal1 s 5796 4658 5796 4658 4 _197_
rlabel metal1 s 5336 3706 5336 3706 4 _198_
rlabel metal2 s 8602 4352 8602 4352 4 _199_
rlabel metal2 s 8610 3910 8610 3910 4 _200_
rlabel metal1 s 8924 4250 8924 4250 4 _201_
rlabel metal1 s 7590 2958 7590 2958 4 _202_
rlabel metal1 s 8356 2890 8356 2890 4 _203_
rlabel metal1 s 7636 2822 7636 2822 4 _204_
rlabel metal1 s 8740 2550 8740 2550 4 _205_
rlabel metal1 s 7820 2482 7820 2482 4 _206_
rlabel metal2 s 9706 2176 9706 2176 4 _207_
rlabel metal2 s 10166 1848 10166 1848 4 _208_
rlabel metal1 s 9476 1870 9476 1870 4 _209_
rlabel metal1 s 12420 3094 12420 3094 4 _210_
rlabel metal1 s 13892 2550 13892 2550 4 _211_
rlabel metal1 s 10534 2482 10534 2482 4 _212_
rlabel metal1 s 10718 1904 10718 1904 4 _213_
rlabel metal1 s 10534 1938 10534 1938 4 _214_
rlabel metal1 s 11178 2006 11178 2006 4 _215_
rlabel metal1 s 13416 2550 13416 2550 4 _216_
rlabel metal1 s 12926 782 12926 782 4 _217_
rlabel metal2 s 13202 3774 13202 3774 4 _218_
rlabel metal1 s 12144 2618 12144 2618 4 _219_
rlabel metal1 s 12926 5576 12926 5576 4 _220_
rlabel metal2 s 12466 3944 12466 3944 4 _221_
rlabel metal1 s 10856 4046 10856 4046 4 _222_
rlabel metal2 s 12190 6324 12190 6324 4 _223_
rlabel metal2 s 11270 6188 11270 6188 4 _224_
rlabel metal1 s 11178 5780 11178 5780 4 _225_
rlabel metal1 s 23874 12954 23874 12954 4 _226_
rlabel metal1 s 25392 12682 25392 12682 4 _227_
rlabel metal1 s 22126 14484 22126 14484 4 _228_
rlabel metal2 s 22218 13435 22218 13435 4 _229_
rlabel metal1 s 22310 14484 22310 14484 4 _230_
rlabel metal1 s 24334 14314 24334 14314 4 _231_
rlabel metal1 s 24794 14586 24794 14586 4 _232_
rlabel metal1 s 16652 11594 16652 11594 4 _233_
rlabel metal1 s 17618 12614 17618 12614 4 _234_
rlabel metal1 s 24380 12818 24380 12818 4 _235_
rlabel metal2 s 25438 14552 25438 14552 4 _236_
rlabel metal2 s 25346 9537 25346 9537 4 _237_
rlabel metal1 s 25668 10234 25668 10234 4 _238_
rlabel metal2 s 24978 13056 24978 13056 4 _239_
rlabel metal2 s 24794 11866 24794 11866 4 _240_
rlabel metal2 s 25898 10778 25898 10778 4 _241_
rlabel metal2 s 25622 7378 25622 7378 4 _242_
rlabel metal1 s 25116 9418 25116 9418 4 _243_
rlabel metal2 s 25346 9180 25346 9180 4 _244_
rlabel metal1 s 26450 6970 26450 6970 4 _245_
rlabel metal1 s 24978 9486 24978 9486 4 _246_
rlabel metal1 s 25990 7718 25990 7718 4 _247_
rlabel metal1 s 25346 7956 25346 7956 4 _248_
rlabel metal2 s 25070 7514 25070 7514 4 _249_
rlabel metal1 s 24056 7310 24056 7310 4 _250_
rlabel metal1 s 24196 7174 24196 7174 4 _251_
rlabel metal1 s 23552 7514 23552 7514 4 _252_
rlabel metal2 s 21114 7650 21114 7650 4 _253_
rlabel metal2 s 24045 9486 24045 9486 4 _254_
rlabel metal1 s 19826 9078 19826 9078 4 _255_
rlabel metal1 s 20470 8976 20470 8976 4 _256_
rlabel metal1 s 21114 9078 21114 9078 4 _257_
rlabel metal1 s 19872 8874 19872 8874 4 _258_
rlabel metal1 s 19504 9622 19504 9622 4 _259_
rlabel metal1 s 24426 10506 24426 10506 4 _260_
rlabel metal2 s 22127 6222 22127 6222 4 _261_
rlabel metal1 s 19964 10778 19964 10778 4 _262_
rlabel metal2 s 20930 10302 20930 10302 4 _263_
rlabel metal2 s 18538 10710 18538 10710 4 _264_
rlabel metal2 s 18630 10965 18630 10965 4 _265_
rlabel metal1 s 17480 8602 17480 8602 4 _266_
rlabel metal1 s 19642 5304 19642 5304 4 _267_
rlabel metal2 s 19182 6256 19182 6256 4 _268_
rlabel metal2 s 12190 10778 12190 10778 4 _269_
rlabel metal1 s 12880 10574 12880 10574 4 _270_
rlabel metal1 s 12006 10064 12006 10064 4 _271_
rlabel metal1 s 13754 9044 13754 9044 4 _272_
rlabel metal1 s 17342 8976 17342 8976 4 _273_
rlabel metal1 s 12926 8330 12926 8330 4 _274_
rlabel metal2 s 12742 7276 12742 7276 4 _275_
rlabel metal1 s 14490 7888 14490 7888 4 _276_
rlabel metal1 s 19182 6256 19182 6256 4 _277_
rlabel metal1 s 21620 782 21620 782 4 _278_
rlabel metal2 s 21479 2482 21479 2482 4 _279_
rlabel metal1 s 21988 2482 21988 2482 4 _280_
rlabel metal1 s 20332 5134 20332 5134 4 _281_
rlabel metal1 s 21850 714 21850 714 4 _282_
rlabel metal1 s 21666 2448 21666 2448 4 _283_
rlabel metal1 s 22494 4590 22494 4590 4 _284_
rlabel metal1 s 22218 3604 22218 3604 4 _285_
rlabel metal1 s 21528 2618 21528 2618 4 _286_
rlabel metal2 s 21758 1530 21758 1530 4 _287_
rlabel metal1 s 23230 748 23230 748 4 _288_
rlabel metal1 s 26266 1904 26266 1904 4 _289_
rlabel metal1 s 25530 1802 25530 1802 4 _290_
rlabel metal1 s 23736 2618 23736 2618 4 _291_
rlabel metal1 s 23138 3910 23138 3910 4 _292_
rlabel metal1 s 15732 7174 15732 7174 4 _293_
rlabel metal2 s 23138 5338 23138 5338 4 _294_
rlabel metal2 s 21942 6120 21942 6120 4 _295_
rlabel metal1 s 20792 7514 20792 7514 4 _296_
rlabel metal1 s 16698 2618 16698 2618 4 _297_
rlabel metal2 s 17986 8636 17986 8636 4 _298_
rlabel metal2 s 16698 10404 16698 10404 4 _299_
rlabel metal1 s 16928 10234 16928 10234 4 _300_
rlabel metal1 s 6900 11322 6900 11322 4 _301_
rlabel metal2 s 8234 11458 8234 11458 4 _302_
rlabel metal1 s 7038 10234 7038 10234 4 _303_
rlabel metal1 s 7774 10608 7774 10608 4 _304_
rlabel metal1 s 6854 9554 6854 9554 4 _305_
rlabel metal1 s 7038 9452 7038 9452 4 _306_
rlabel metal1 s 7682 9146 7682 9146 4 _307_
rlabel metal2 s 9706 9248 9706 9248 4 _308_
rlabel metal2 s 7038 8738 7038 8738 4 _309_
rlabel metal1 s 7682 9044 7682 9044 4 _310_
rlabel metal1 s 10718 8534 10718 8534 4 _311_
rlabel metal1 s 11730 8500 11730 8500 4 _312_
rlabel metal1 s 9614 7956 9614 7956 4 _313_
rlabel metal2 s 8694 7140 8694 7140 4 _314_
rlabel metal1 s 15318 2448 15318 2448 4 _315_
rlabel metal1 s 15594 2448 15594 2448 4 _316_
rlabel metal2 s 15410 5916 15410 5916 4 _317_
rlabel metal1 s 17342 5678 17342 5678 4 _318_
rlabel metal2 s 15318 4250 15318 4250 4 _319_
rlabel metal1 s 16146 4012 16146 4012 4 _320_
rlabel metal1 s 19412 1870 19412 1870 4 _321_
rlabel metal1 s 15502 3604 15502 3604 4 _322_
rlabel metal2 s 15134 2074 15134 2074 4 _323_
rlabel metal1 s 17342 2516 17342 2516 4 _324_
rlabel metal2 s 19642 1156 19642 1156 4 _325_
rlabel metal1 s 17434 1224 17434 1224 4 _326_
rlabel metal2 s 18078 2108 18078 2108 4 _327_
rlabel metal1 s 12834 9146 12834 9146 4 _328_
rlabel metal2 s 18630 4182 18630 4182 4 _329_
rlabel metal1 s 17342 4692 17342 4692 4 _330_
rlabel metal1 s 16422 5338 16422 5338 4 _331_
rlabel metal1 s 14490 6834 14490 6834 4 _332_
rlabel metal1 s 16652 16150 16652 16150 4 _333_
rlabel metal2 s 17802 13260 17802 13260 4 _334_
rlabel metal1 s 19734 16014 19734 16014 4 _335_
rlabel metal1 s 20378 16048 20378 16048 4 _336_
rlabel metal2 s 10074 16048 10074 16048 4 _337_
rlabel metal2 s 5474 14416 5474 14416 4 _338_
rlabel metal1 s 8234 13158 8234 13158 4 _339_
rlabel metal1 s 7774 15504 7774 15504 4 _340_
rlabel metal3 s 9614 13923 9614 13923 4 _341_
rlabel metal1 s 8878 15130 8878 15130 4 _342_
rlabel metal1 s 9338 14518 9338 14518 4 _343_
rlabel metal2 s 8878 14042 8878 14042 4 _344_
rlabel metal2 s 11178 15130 11178 15130 4 _345_
rlabel metal2 s 11454 13226 11454 13226 4 _346_
rlabel metal1 s 9016 16218 9016 16218 4 _347_
rlabel metal2 s 7866 14042 7866 14042 4 _348_
rlabel metal1 s 3450 12716 3450 12716 4 _349_
rlabel metal1 s 3036 11662 3036 11662 4 _350_
rlabel metal2 s 4830 15130 4830 15130 4 _351_
rlabel metal1 s 5520 15130 5520 15130 4 _352_
rlabel metal1 s 3910 12784 3910 12784 4 _353_
rlabel metal1 s 3082 12784 3082 12784 4 _354_
rlabel metal1 s 3910 15538 3910 15538 4 _355_
rlabel metal2 s 3358 15844 3358 15844 4 _356_
rlabel metal1 s 4186 14450 4186 14450 4 _357_
rlabel metal1 s 3174 13838 3174 13838 4 _358_
rlabel metal1 s 9338 13906 9338 13906 4 _359_
rlabel metal3 s 8050 13821 8050 13821 4 _360_
rlabel metal1 s 8418 12750 8418 12750 4 _361_
rlabel metal2 s 12282 15402 12282 15402 4 _362_
rlabel metal2 s 12098 16014 12098 16014 4 _363_
rlabel metal2 s 12742 12954 12742 12954 4 _364_
rlabel metal1 s 12972 12750 12972 12750 4 _365_
rlabel metal1 s 10212 12750 10212 12750 4 _366_
rlabel metal1 s 9430 12070 9430 12070 4 _367_
rlabel metal1 s 18078 16048 18078 16048 4 _368_
rlabel metal1 s 18308 16014 18308 16014 4 _369_
rlabel metal1 s 16974 13294 16974 13294 4 _370_
rlabel metal2 s 15962 12954 15962 12954 4 _371_
rlabel metal2 s 17158 14620 17158 14620 4 _372_
rlabel metal1 s 17848 14586 17848 14586 4 _373_
rlabel metal1 s 18262 14042 18262 14042 4 _374_
rlabel metal1 s 18860 14450 18860 14450 4 _375_
rlabel metal1 s 18906 13872 18906 13872 4 _376_
rlabel metal1 s 19228 13838 19228 13838 4 _377_
rlabel metal1 s 18170 15130 18170 15130 4 _378_
rlabel metal1 s 19136 15538 19136 15538 4 _379_
rlabel metal1 s 18860 12750 18860 12750 4 _380_
rlabel metal1 s 19044 12614 19044 12614 4 _381_
rlabel metal3 s 15778 9435 15778 9435 4 clk
rlabel metal3 s 14030 9571 14030 9571 4 clknet_0_clk
rlabel metal1 s 1748 7922 1748 7922 4 clknet_3_0__leaf_clk
rlabel metal1 s 10994 1258 10994 1258 4 clknet_3_1__leaf_clk
rlabel metal2 s 2530 11390 2530 11390 4 clknet_3_2__leaf_clk
rlabel metal1 s 14260 10574 14260 10574 4 clknet_3_3__leaf_clk
rlabel metal1 s 19136 1394 19136 1394 4 clknet_3_4__leaf_clk
rlabel metal1 s 20010 1938 20010 1938 4 clknet_3_5__leaf_clk
rlabel metal1 s 16284 12818 16284 12818 4 clknet_3_6__leaf_clk
rlabel metal1 s 21482 15538 21482 15538 4 clknet_3_7__leaf_clk
rlabel metal1 s 20102 15606 20102 15606 4 net1
rlabel metal1 s 19872 16966 19872 16966 4 net10
rlabel metal1 s 17158 2448 17158 2448 4 net100
rlabel metal1 s 11960 2346 11960 2346 4 net101
rlabel metal1 s 24334 14960 24334 14960 4 net102
rlabel metal2 s 5290 7514 5290 7514 4 net103
rlabel metal1 s 2024 9418 2024 9418 4 net104
rlabel metal1 s 1881 9078 1881 9078 4 net105
rlabel metal1 s 4646 10098 4646 10098 4 net106
rlabel metal1 s 25530 9044 25530 9044 4 net107
rlabel metal2 s 8326 3876 8326 3876 4 net108
rlabel metal1 s 3266 8364 3266 8364 4 net109
rlabel metal1 s 15916 17170 15916 17170 4 net11
rlabel metal1 s 26266 6834 26266 6834 4 net110
rlabel metal2 s 26082 7684 26082 7684 4 net111
rlabel metal2 s 12374 8483 12374 8483 4 net112
rlabel metal2 s 17250 10302 17250 10302 4 net113
rlabel metal1 s 11178 9350 11178 9350 4 net114
rlabel metal2 s 9706 10744 9706 10744 4 net115
rlabel metal1 s 10672 10166 10672 10166 4 net116
rlabel metal2 s 8234 9894 8234 9894 4 net117
rlabel metal1 s 8740 11526 8740 11526 4 net118
rlabel metal1 s 24886 7276 24886 7276 4 net119
rlabel metal1 s 17572 16694 17572 16694 4 net12
rlabel metal1 s 5336 6222 5336 6222 4 net120
rlabel metal1 s 5750 3570 5750 3570 4 net121
rlabel metal1 s 22816 14450 22816 14450 4 net122
rlabel metal1 s 14996 9146 14996 9146 4 net123
rlabel metal1 s 25300 12342 25300 12342 4 net124
rlabel metal1 s 6578 8398 6578 8398 4 net125
rlabel metal1 s 11086 2516 11086 2516 4 net126
rlabel metal2 s 12006 6052 12006 6052 4 net127
rlabel metal1 s 14122 4624 14122 4624 4 net128
rlabel metal1 s 14306 4998 14306 4998 4 net129
rlabel metal2 s 17526 16864 17526 16864 4 net13
rlabel metal1 s 3864 17306 3864 17306 4 net14
rlabel metal2 s 2714 17520 2714 17520 4 net15
rlabel metal2 s 2162 17527 2162 17527 4 net16
rlabel metal1 s 9246 17306 9246 17306 4 net17
rlabel metal1 s 7912 17306 7912 17306 4 net18
rlabel metal2 s 7314 17527 7314 17527 4 net19
rlabel metal1 s 20286 15980 20286 15980 4 net2
rlabel metal1 s 5336 17170 5336 17170 4 net20
rlabel metal1 s 4692 17170 4692 17170 4 net21
rlabel metal2 s 3450 17459 3450 17459 4 net22
rlabel metal1 s 3036 10030 3036 10030 4 net23
rlabel metal1 s 11270 12716 11270 12716 4 net24
rlabel metal1 s 13938 7242 13938 7242 4 net25
rlabel metal2 s 12374 7718 12374 7718 4 net26
rlabel metal1 s 23874 4454 23874 4454 4 net27
rlabel metal2 s 21109 4046 21109 4046 4 net28
rlabel metal2 s 8694 14314 8694 14314 4 net29
rlabel metal1 s 23690 16660 23690 16660 4 net3
rlabel metal2 s 22476 782 22476 782 4 net30
rlabel metal1 s 21339 1802 21339 1802 4 net31
rlabel metal2 s 5658 13668 5658 13668 4 net32
rlabel metal2 s 10994 15164 10994 15164 4 net33
rlabel metal1 s 21895 7242 21895 7242 4 net34
rlabel metal1 s 22596 6834 22596 6834 4 net35
rlabel metal2 s 18998 6426 18998 6426 4 net36
rlabel metal1 s 18114 6834 18114 6834 4 net37
rlabel metal1 s 5980 13158 5980 13158 4 net38
rlabel metal2 s 21574 3366 21574 3366 4 net39
rlabel metal1 s 23046 17170 23046 17170 4 net4
rlabel metal1 s 20281 2890 20281 2890 4 net40
rlabel metal1 s 20792 5134 20792 5134 4 net41
rlabel metal1 s 20945 6154 20945 6154 4 net42
rlabel metal1 s 15410 7922 15410 7922 4 net43
rlabel metal2 s 14853 7310 14853 7310 4 net44
rlabel metal1 s 24840 1530 24840 1530 4 net45
rlabel metal1 s 23552 986 23552 986 4 net46
rlabel metal2 s 15226 6188 15226 6188 4 net47
rlabel metal1 s 14904 6426 14904 6426 4 net48
rlabel metal2 s 18170 8228 18170 8228 4 net49
rlabel metal1 s 22954 16048 22954 16048 4 net5
rlabel metal1 s 20884 7922 20884 7922 4 net50
rlabel metal2 s 22406 7922 22406 7922 4 net51
rlabel metal1 s 9982 7922 9982 7922 4 net52
rlabel metal1 s 18078 7344 18078 7344 4 net53
rlabel metal2 s 19366 7038 19366 7038 4 net54
rlabel metal1 s 5290 15980 5290 15980 4 net55
rlabel metal1 s 5382 14960 5382 14960 4 net56
rlabel metal1 s 24886 2550 24886 2550 4 net57
rlabel metal1 s 25341 2482 25341 2482 4 net58
rlabel metal1 s 23414 5134 23414 5134 4 net59
rlabel metal1 s 23414 16626 23414 16626 4 net6
rlabel metal1 s 24620 5746 24620 5746 4 net60
rlabel metal2 s 7590 15980 7590 15980 4 net61
rlabel metal1 s 17158 5780 17158 5780 4 net62
rlabel metal2 s 16146 6018 16146 6018 4 net63
rlabel metal1 s 24058 4658 24058 4658 4 net64
rlabel metal1 s 25177 5066 25177 5066 4 net65
rlabel metal2 s 24334 11322 24334 11322 4 net66
rlabel metal2 s 12742 4352 12742 4352 4 net67
rlabel metal1 s 25530 986 25530 986 4 net68
rlabel metal1 s 25085 1462 25085 1462 4 net69
rlabel metal1 s 22816 16626 22816 16626 4 net7
rlabel metal1 s 12834 3400 12834 3400 4 net70
rlabel metal2 s 7125 3638 7125 3638 4 net71
rlabel metal1 s 6992 8058 6992 8058 4 net72
rlabel metal2 s 22402 3366 22402 3366 4 net73
rlabel metal1 s 24303 3638 24303 3638 4 net74
rlabel metal1 s 8878 7242 8878 7242 4 net75
rlabel metal1 s 10058 7242 10058 7242 4 net76
rlabel metal1 s 20378 782 20378 782 4 net77
rlabel metal1 s 24794 2958 24794 2958 4 net78
rlabel metal1 s 24564 3162 24564 3162 4 net79
rlabel metal2 s 22126 16796 22126 16796 4 net8
rlabel metal1 s 18262 5780 18262 5780 4 net80
rlabel metal1 s 18584 1870 18584 1870 4 net81
rlabel metal1 s 19085 2550 19085 2550 4 net82
rlabel metal1 s 19228 3570 19228 3570 4 net83
rlabel metal1 s 12098 6188 12098 6188 4 net84
rlabel metal2 s 10994 6188 10994 6188 4 net85
rlabel metal1 s 23414 7888 23414 7888 4 net86
rlabel metal2 s 15686 3366 15686 3366 4 net87
rlabel metal1 s 16330 4012 16330 4012 4 net88
rlabel metal2 s 17618 3842 17618 3842 4 net89
rlabel metal2 s 21482 16796 21482 16796 4 net9
rlabel metal2 s 18998 1428 18998 1428 4 net90
rlabel metal2 s 19366 1088 19366 1088 4 net91
rlabel metal2 s 15180 4046 15180 4046 4 net92
rlabel metal1 s 17158 4624 17158 4624 4 net93
rlabel metal1 s 17234 5066 17234 5066 4 net94
rlabel metal1 s 12190 6358 12190 6358 4 net95
rlabel metal1 s 15318 1836 15318 1836 4 net96
rlabel metal2 s 15957 1870 15957 1870 4 net97
rlabel metal1 s 9476 6222 9476 6222 4 net98
rlabel metal2 s 7406 5542 7406 5542 4 net99
rlabel metal2 s 874 1911 874 1911 4 o_digital[0]
rlabel metal4 s 18331 4012 18331 4012 4 o_digital[10]
rlabel metal2 s 20102 1557 20102 1557 4 o_digital[11]
rlabel metal2 s 21850 1367 21850 1367 4 o_digital[12]
rlabel metal1 s 22770 12682 22770 12682 4 o_digital[13]
rlabel metal4 s 22379 13804 22379 13804 4 o_digital[14]
rlabel metal1 s 25438 11866 25438 11866 4 o_digital[15]
rlabel metal2 s 2622 1690 2622 1690 4 o_digital[1]
rlabel metal1 s 4416 11118 4416 11118 4 o_digital[2]
rlabel metal2 s 6118 415 6118 415 4 o_digital[3]
rlabel metal2 s 7866 1557 7866 1557 4 o_digital[4]
rlabel metal2 s 9614 1557 9614 1557 4 o_digital[5]
rlabel metal2 s 11362 415 11362 415 4 o_digital[6]
rlabel metal2 s 13110 6212 13110 6212 4 o_digital[7]
rlabel metal2 s 14858 891 14858 891 4 o_digital[8]
rlabel metal2 s 16560 4148 16560 4148 4 o_digital[9]
rlabel metal2 s 26818 17425 26818 17425 4 rst_n
rlabel metal1 s 26036 17102 26036 17102 4 ui_in[0]
rlabel metal1 s 25392 17102 25392 17102 4 ui_in[1]
rlabel metal1 s 24748 17102 24748 17102 4 ui_in[2]
rlabel metal2 s 24334 17306 24334 17306 4 ui_in[3]
rlabel metal1 s 24058 17136 24058 17136 4 ui_in[4]
rlabel metal1 s 23506 17068 23506 17068 4 ui_in[5]
rlabel metal2 s 22034 17418 22034 17418 4 ui_in[6]
rlabel metal2 s 21666 17425 21666 17425 4 ui_in[7]
rlabel metal1 s 19596 17102 19596 17102 4 uio_in[2]
rlabel metal2 s 18262 17425 18262 17425 4 uio_in[4]
rlabel metal1 s 17756 17102 17756 17102 4 uio_in[5]
rlabel metal1 s 17434 17136 17434 17136 4 uio_in[6]
rlabel metal2 s 1426 14528 1426 14528 4 uio_oe[6]
rlabel metal1 s 1242 16762 1242 16762 4 uio_oe[7]
rlabel metal2 s 23782 15878 23782 15878 4 uio_out[0]
rlabel metal1 s 9982 17306 9982 17306 4 uio_out[1]
rlabel metal2 s 8510 16381 8510 16381 4 uio_out[3]
rlabel metal1 s 7682 17102 7682 17102 4 uio_out[6]
rlabel metal1 s 6118 16762 6118 16762 4 uio_out[7]
rlabel metal1 s 15962 16762 15962 16762 4 uo_out[0]
rlabel metal1 s 14306 16592 14306 16592 4 uo_out[1]
rlabel metal1 s 13984 16762 13984 16762 4 uo_out[2]
rlabel metal1 s 13570 16762 13570 16762 4 uo_out[3]
rlabel metal1 s 12972 17306 12972 17306 4 uo_out[4]
rlabel metal2 s 12374 17520 12374 17520 4 uo_out[5]
rlabel metal1 s 11638 16762 11638 16762 4 uo_out[6]
rlabel metal1 s 11132 16762 11132 16762 4 uo_out[7]
rlabel metal1 s 17710 16558 17710 16558 4 wrapped.o_busy
rlabel metal2 s 10350 17306 10350 17306 4 wrapped.o_copi
rlabel metal1 s 24794 14314 24794 14314 4 wrapped.o_cs_n
rlabel metal1 s 14352 13702 14352 13702 4 wrapped.o_data\[0\]
rlabel metal2 s 11270 11186 11270 11186 4 wrapped.o_data\[1\]
rlabel metal1 s 11418 10608 11418 10608 4 wrapped.o_data\[2\]
rlabel metal1 s 14030 15878 14030 15878 4 wrapped.o_data\[3\]
rlabel metal2 s 11712 9486 11712 9486 4 wrapped.o_data\[4\]
rlabel metal1 s 13938 8976 13938 8976 4 wrapped.o_data\[5\]
rlabel metal2 s 17526 14858 17526 14858 4 wrapped.o_data\[6\]
rlabel metal1 s 18078 12682 18078 12682 4 wrapped.o_data\[7\]
rlabel metal1 s 16974 16558 16974 16558 4 wrapped.o_data_valid
rlabel metal1 s 15088 13362 15088 13362 4 wrapped.o_digital$17\[0\]
rlabel metal2 s 16146 13532 16146 13532 4 wrapped.o_digital$17\[10\]
rlabel metal1 s 19918 15062 19918 15062 4 wrapped.o_digital$17\[11\]
rlabel metal1 s 17526 13838 17526 13838 4 wrapped.o_digital$17\[12\]
rlabel metal1 s 16928 13838 16928 13838 4 wrapped.o_digital$17\[13\]
rlabel metal2 s 21114 15062 21114 15062 4 wrapped.o_digital$17\[14\]
rlabel metal1 s 20976 12274 20976 12274 4 wrapped.o_digital$17\[15\]
rlabel metal2 s 5658 17136 5658 17136 4 wrapped.o_digital$17\[1\]
rlabel metal2 s 4738 13532 4738 13532 4 wrapped.o_digital$17\[2\]
rlabel metal1 s 5796 16150 5796 16150 4 wrapped.o_digital$17\[3\]
rlabel metal3 s 13938 14875 13938 14875 4 wrapped.o_digital$17\[4\]
rlabel metal1 s 9706 13804 9706 13804 4 wrapped.o_digital$17\[5\]
rlabel metal1 s 13386 16422 13386 16422 4 wrapped.o_digital$17\[6\]
rlabel metal2 s 13478 13226 13478 13226 4 wrapped.o_digital$17\[7\]
rlabel metal1 s 14812 13294 14812 13294 4 wrapped.o_digital$17\[8\]
rlabel metal1 s 17066 16014 17066 16014 4 wrapped.o_digital$17\[9\]
rlabel metal1 s 24610 14824 24610 14824 4 wrapped.o_sclk
rlabel metal1 s 13455 6154 13455 6154 4 wrapped.o_spi_address\[10\]
rlabel metal2 s 14490 5695 14490 5695 4 wrapped.o_spi_address\[11\]
rlabel metal2 s 9154 3706 9154 3706 4 wrapped.o_spi_address\[12\]
rlabel metal1 s 13409 3978 13409 3978 4 wrapped.o_spi_address\[13\]
rlabel metal1 s 9062 3468 9062 3468 4 wrapped.o_spi_address\[14\]
rlabel metal1 s 14536 2618 14536 2618 4 wrapped.o_spi_address\[15\]
rlabel metal1 s 12834 2924 12834 2924 4 wrapped.o_spi_address\[16\]
rlabel metal1 s 13662 2414 13662 2414 4 wrapped.o_spi_address\[17\]
rlabel metal1 s 13570 1190 13570 1190 4 wrapped.o_spi_address\[18\]
rlabel metal1 s 14122 1496 14122 1496 4 wrapped.o_spi_address\[19\]
rlabel metal1 s 5290 10676 5290 10676 4 wrapped.o_spi_address\[1\]
rlabel metal2 s 12558 2655 12558 2655 4 wrapped.o_spi_address\[20\]
rlabel metal1 s 12834 4250 12834 4250 4 wrapped.o_spi_address\[21\]
rlabel metal1 s 13570 5270 13570 5270 4 wrapped.o_spi_address\[22\]
rlabel metal2 s 13570 6154 13570 6154 4 wrapped.o_spi_address\[23\]
rlabel metal2 s 5106 10574 5106 10574 4 wrapped.o_spi_address\[2\]
rlabel metal2 s 3818 9316 3818 9316 4 wrapped.o_spi_address\[3\]
rlabel metal1 s 5750 9486 5750 9486 4 wrapped.o_spi_address\[4\]
rlabel metal2 s 6118 8466 6118 8466 4 wrapped.o_spi_address\[5\]
rlabel metal1 s 6072 8058 6072 8058 4 wrapped.o_spi_address\[6\]
rlabel metal1 s 6716 7854 6716 7854 4 wrapped.o_spi_address\[7\]
rlabel metal1 s 7498 6256 7498 6256 4 wrapped.o_spi_address\[8\]
rlabel metal2 s 9062 5338 9062 5338 4 wrapped.o_spi_address\[9\]
rlabel metal2 s 5014 13124 5014 13124 4 wrapped.player.buffer\[0\]
rlabel metal1 s 6670 16218 6670 16218 4 wrapped.player.buffer\[1\]
rlabel metal1 s 4370 13430 4370 13430 4 wrapped.player.buffer\[2\]
rlabel metal2 s 6302 15844 6302 15844 4 wrapped.player.buffer\[3\]
rlabel metal2 s 6394 14756 6394 14756 4 wrapped.player.buffer\[4\]
rlabel metal2 s 8970 14756 8970 14756 4 wrapped.player.buffer\[5\]
rlabel metal2 s 12006 15742 12006 15742 4 wrapped.player.buffer\[6\]
rlabel metal1 s 12650 13226 12650 13226 4 wrapped.player.buffer\[7\]
rlabel metal1 s 9246 17068 9246 17068 4 wrapped.player.received_samples
rlabel metal1 s 20010 8602 20010 8602 4 wrapped.spi_flash.address\[0\]
rlabel metal2 s 16422 7106 16422 7106 4 wrapped.spi_flash.address\[10\]
rlabel metal1 s 17986 6222 17986 6222 4 wrapped.spi_flash.address\[11\]
rlabel metal1 s 16790 4556 16790 4556 4 wrapped.spi_flash.address\[12\]
rlabel metal1 s 18078 2958 18078 2958 4 wrapped.spi_flash.address\[13\]
rlabel metal1 s 18814 2482 18814 2482 4 wrapped.spi_flash.address\[14\]
rlabel metal1 s 18308 1938 18308 1938 4 wrapped.spi_flash.address\[15\]
rlabel metal1 s 18262 2346 18262 2346 4 wrapped.spi_flash.address\[16\]
rlabel metal1 s 22310 1938 22310 1938 4 wrapped.spi_flash.address\[17\]
rlabel metal2 s 17710 1513 17710 1513 4 wrapped.spi_flash.address\[18\]
rlabel metal1 s 20654 2516 20654 2516 4 wrapped.spi_flash.address\[19\]
rlabel metal2 s 17986 10846 17986 10846 4 wrapped.spi_flash.address\[1\]
rlabel metal1 s 21574 3910 21574 3910 4 wrapped.spi_flash.address\[20\]
rlabel metal1 s 20056 4658 20056 4658 4 wrapped.spi_flash.address\[21\]
rlabel metal1 s 20930 5678 20930 5678 4 wrapped.spi_flash.address\[22\]
rlabel metal1 s 20746 7412 20746 7412 4 wrapped.spi_flash.address\[23\]
rlabel metal2 s 8142 11492 8142 11492 4 wrapped.spi_flash.address\[2\]
rlabel metal1 s 9844 10778 9844 10778 4 wrapped.spi_flash.address\[3\]
rlabel metal1 s 8970 9996 8970 9996 4 wrapped.spi_flash.address\[4\]
rlabel metal2 s 9614 9316 9614 9316 4 wrapped.spi_flash.address\[5\]
rlabel metal1 s 9798 8296 9798 8296 4 wrapped.spi_flash.address\[6\]
rlabel metal2 s 12374 9316 12374 9316 4 wrapped.spi_flash.address\[7\]
rlabel metal1 s 10810 7956 10810 7956 4 wrapped.spi_flash.address\[8\]
rlabel metal1 s 13202 7412 13202 7412 4 wrapped.spi_flash.address\[9\]
rlabel metal2 s 17710 11934 17710 11934 4 wrapped.spi_flash.fsm_state\[0\]
rlabel metal2 s 21114 9962 21114 9962 4 wrapped.spi_flash.fsm_state\[1\]
rlabel metal2 s 21298 11322 21298 11322 4 wrapped.spi_flash.fsm_state\[2\]
rlabel metal1 s 22632 9894 22632 9894 4 wrapped.spi_flash.fsm_state\[3\]
rlabel metal2 s 26174 11356 26174 11356 4 wrapped.spi_flash.fsm_state\[4\]
rlabel metal1 s 20746 6732 20746 6732 4 wrapped.spi_flash.shift_reg\[10\]
rlabel metal2 s 20378 5916 20378 5916 4 wrapped.spi_flash.shift_reg\[11\]
rlabel metal1 s 22494 4250 22494 4250 4 wrapped.spi_flash.shift_reg\[12\]
rlabel metal2 s 21849 2482 21849 2482 4 wrapped.spi_flash.shift_reg\[13\]
rlabel metal1 s 21942 3060 21942 3060 4 wrapped.spi_flash.shift_reg\[14\]
rlabel metal1 s 23074 1938 23074 1938 4 wrapped.spi_flash.shift_reg\[15\]
rlabel metal1 s 25438 1360 25438 1360 4 wrapped.spi_flash.shift_reg\[16\]
rlabel metal1 s 23460 1190 23460 1190 4 wrapped.spi_flash.shift_reg\[17\]
rlabel metal1 s 25438 2380 25438 2380 4 wrapped.spi_flash.shift_reg\[18\]
rlabel metal3 s 25622 3723 25622 3723 4 wrapped.spi_flash.shift_reg\[19\]
rlabel metal1 s 23828 5270 23828 5270 4 wrapped.spi_flash.shift_reg\[20\]
rlabel metal1 s 23920 5882 23920 5882 4 wrapped.spi_flash.shift_reg\[21\]
rlabel metal1 s 21482 6970 21482 6970 4 wrapped.spi_flash.shift_reg\[22\]
rlabel metal2 s 21298 9112 21298 9112 4 wrapped.spi_flash.shift_reg\[23\]
rlabel metal2 s 13570 7548 13570 7548 4 wrapped.spi_flash.shift_reg\[8\]
rlabel metal2 s 15962 7684 15962 7684 4 wrapped.spi_flash.shift_reg\[9\]
rlabel metal2 s 26818 7344 26818 7344 4 wrapped.spi_flash.timer\[0\]
rlabel metal2 s 27002 6596 27002 6596 4 wrapped.spi_flash.timer\[1\]
rlabel metal2 s 25898 7140 25898 7140 4 wrapped.spi_flash.timer\[2\]
rlabel metal1 s 24610 8908 24610 8908 4 wrapped.spi_flash.timer\[3\]
rlabel metal2 s 22494 9044 22494 9044 4 wrapped.spi_flash.timer\[4\]
flabel metal4 s 27256 496 27576 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 20540 496 20860 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 13824 496 14144 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7108 496 7428 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 23898 496 24218 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 17182 496 17502 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 10466 496 10786 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3750 496 4070 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 27158 17600 27214 18000 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal2 s 846 0 902 400 0 FreeSans 280 90 0 0 o_digital[0]
port 4 nsew
flabel metal2 s 18326 0 18382 400 0 FreeSans 280 90 0 0 o_digital[10]
port 5 nsew
flabel metal2 s 20074 0 20130 400 0 FreeSans 280 90 0 0 o_digital[11]
port 6 nsew
flabel metal2 s 21822 0 21878 400 0 FreeSans 280 90 0 0 o_digital[12]
port 7 nsew
flabel metal2 s 23570 0 23626 400 0 FreeSans 280 90 0 0 o_digital[13]
port 8 nsew
flabel metal2 s 25318 0 25374 400 0 FreeSans 280 90 0 0 o_digital[14]
port 9 nsew
flabel metal2 s 27066 0 27122 400 0 FreeSans 280 90 0 0 o_digital[15]
port 10 nsew
flabel metal2 s 2594 0 2650 400 0 FreeSans 280 90 0 0 o_digital[1]
port 11 nsew
flabel metal2 s 4342 0 4398 400 0 FreeSans 280 90 0 0 o_digital[2]
port 12 nsew
flabel metal2 s 6090 0 6146 400 0 FreeSans 280 90 0 0 o_digital[3]
port 13 nsew
flabel metal2 s 7838 0 7894 400 0 FreeSans 280 90 0 0 o_digital[4]
port 14 nsew
flabel metal2 s 9586 0 9642 400 0 FreeSans 280 90 0 0 o_digital[5]
port 15 nsew
flabel metal2 s 11334 0 11390 400 0 FreeSans 280 90 0 0 o_digital[6]
port 16 nsew
flabel metal2 s 13082 0 13138 400 0 FreeSans 280 90 0 0 o_digital[7]
port 17 nsew
flabel metal2 s 14830 0 14886 400 0 FreeSans 280 90 0 0 o_digital[8]
port 18 nsew
flabel metal2 s 16578 0 16634 400 0 FreeSans 280 90 0 0 o_digital[9]
port 19 nsew
flabel metal2 s 26514 17600 26570 18000 0 FreeSans 280 90 0 0 rst_n
port 20 nsew
flabel metal2 s 25870 17600 25926 18000 0 FreeSans 280 90 0 0 ui_in[0]
port 21 nsew
flabel metal2 s 25226 17600 25282 18000 0 FreeSans 280 90 0 0 ui_in[1]
port 22 nsew
flabel metal2 s 24582 17600 24638 18000 0 FreeSans 280 90 0 0 ui_in[2]
port 23 nsew
flabel metal2 s 23938 17600 23994 18000 0 FreeSans 280 90 0 0 ui_in[3]
port 24 nsew
flabel metal2 s 23294 17600 23350 18000 0 FreeSans 280 90 0 0 ui_in[4]
port 25 nsew
flabel metal2 s 22650 17600 22706 18000 0 FreeSans 280 90 0 0 ui_in[5]
port 26 nsew
flabel metal2 s 22006 17600 22062 18000 0 FreeSans 280 90 0 0 ui_in[6]
port 27 nsew
flabel metal2 s 21362 17600 21418 18000 0 FreeSans 280 90 0 0 ui_in[7]
port 28 nsew
flabel metal2 s 20718 17600 20774 18000 0 FreeSans 280 90 0 0 uio_in[0]
port 29 nsew
flabel metal2 s 20074 17600 20130 18000 0 FreeSans 280 90 0 0 uio_in[1]
port 30 nsew
flabel metal2 s 19430 17600 19486 18000 0 FreeSans 280 90 0 0 uio_in[2]
port 31 nsew
flabel metal2 s 18786 17600 18842 18000 0 FreeSans 280 90 0 0 uio_in[3]
port 32 nsew
flabel metal2 s 18142 17600 18198 18000 0 FreeSans 280 90 0 0 uio_in[4]
port 33 nsew
flabel metal2 s 17498 17600 17554 18000 0 FreeSans 280 90 0 0 uio_in[5]
port 34 nsew
flabel metal2 s 16854 17600 16910 18000 0 FreeSans 280 90 0 0 uio_in[6]
port 35 nsew
flabel metal2 s 16210 17600 16266 18000 0 FreeSans 280 90 0 0 uio_in[7]
port 36 nsew
flabel metal2 s 5262 17600 5318 18000 0 FreeSans 280 90 0 0 uio_oe[0]
port 37 nsew
flabel metal2 s 4618 17600 4674 18000 0 FreeSans 280 90 0 0 uio_oe[1]
port 38 nsew
flabel metal2 s 3974 17600 4030 18000 0 FreeSans 280 90 0 0 uio_oe[2]
port 39 nsew
flabel metal2 s 3330 17600 3386 18000 0 FreeSans 280 90 0 0 uio_oe[3]
port 40 nsew
flabel metal2 s 2686 17600 2742 18000 0 FreeSans 280 90 0 0 uio_oe[4]
port 41 nsew
flabel metal2 s 2042 17600 2098 18000 0 FreeSans 280 90 0 0 uio_oe[5]
port 42 nsew
flabel metal2 s 1398 17600 1454 18000 0 FreeSans 280 90 0 0 uio_oe[6]
port 43 nsew
flabel metal2 s 754 17600 810 18000 0 FreeSans 280 90 0 0 uio_oe[7]
port 44 nsew
flabel metal2 s 10414 17600 10470 18000 0 FreeSans 280 90 0 0 uio_out[0]
port 45 nsew
flabel metal2 s 9770 17600 9826 18000 0 FreeSans 280 90 0 0 uio_out[1]
port 46 nsew
flabel metal2 s 9126 17600 9182 18000 0 FreeSans 280 90 0 0 uio_out[2]
port 47 nsew
flabel metal2 s 8482 17600 8538 18000 0 FreeSans 280 90 0 0 uio_out[3]
port 48 nsew
flabel metal2 s 7838 17600 7894 18000 0 FreeSans 280 90 0 0 uio_out[4]
port 49 nsew
flabel metal2 s 7194 17600 7250 18000 0 FreeSans 280 90 0 0 uio_out[5]
port 50 nsew
flabel metal2 s 6550 17600 6606 18000 0 FreeSans 280 90 0 0 uio_out[6]
port 51 nsew
flabel metal2 s 5906 17600 5962 18000 0 FreeSans 280 90 0 0 uio_out[7]
port 52 nsew
flabel metal2 s 15566 17600 15622 18000 0 FreeSans 280 90 0 0 uo_out[0]
port 53 nsew
flabel metal2 s 14922 17600 14978 18000 0 FreeSans 280 90 0 0 uo_out[1]
port 54 nsew
flabel metal2 s 14278 17600 14334 18000 0 FreeSans 280 90 0 0 uo_out[2]
port 55 nsew
flabel metal2 s 13634 17600 13690 18000 0 FreeSans 280 90 0 0 uo_out[3]
port 56 nsew
flabel metal2 s 12990 17600 13046 18000 0 FreeSans 280 90 0 0 uo_out[4]
port 57 nsew
flabel metal2 s 12346 17600 12402 18000 0 FreeSans 280 90 0 0 uo_out[5]
port 58 nsew
flabel metal2 s 11702 17600 11758 18000 0 FreeSans 280 90 0 0 uo_out[6]
port 59 nsew
flabel metal2 s 11058 17600 11114 18000 0 FreeSans 280 90 0 0 uo_out[7]
port 60 nsew
<< properties >>
string FIXED_BBOX 0 0 28000 18000
string GDS_END 1923552
string GDS_FILE ../gds/digital_top.gds
string GDS_START 376800
<< end >>
