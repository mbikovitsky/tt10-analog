magic
tech sky130A
magscale 1 2
timestamp 1757953533
<< checkpaint >>
rect -746 -1260 28836 19260
<< viali >>
rect 857 17289 891 17323
rect 1501 17289 1535 17323
rect 4077 17289 4111 17323
rect 5641 17289 5675 17323
rect 6837 17289 6871 17323
rect 9229 17289 9263 17323
rect 12449 17289 12483 17323
rect 13185 17289 13219 17323
rect 16313 17289 16347 17323
rect 23397 17289 23431 17323
rect 6653 17221 6687 17255
rect 12817 17221 12851 17255
rect 15669 17221 15703 17255
rect 17601 17221 17635 17255
rect 19993 17221 20027 17255
rect 2789 17153 2823 17187
rect 3433 17153 3467 17187
rect 4721 17153 4755 17187
rect 5365 17153 5399 17187
rect 6285 17153 6319 17187
rect 6469 17085 6503 17119
rect 10057 17085 10091 17119
rect 10149 17085 10183 17119
rect 10241 17085 10275 17119
rect 10425 17085 10459 17119
rect 11529 17085 11563 17119
rect 12633 17085 12667 17119
rect 13001 17085 13035 17119
rect 13369 17085 13403 17119
rect 14381 17085 14415 17119
rect 15301 17085 15335 17119
rect 15485 17085 15519 17119
rect 16129 17085 16163 17119
rect 16497 17085 16531 17119
rect 16957 17085 16991 17119
rect 17785 17085 17819 17119
rect 20453 17085 20487 17119
rect 21649 17085 21683 17119
rect 22293 17085 22327 17119
rect 22937 17085 22971 17119
rect 23581 17085 23615 17119
rect 24225 17085 24259 17119
rect 24869 17085 24903 17119
rect 25789 17085 25823 17119
rect 26157 17085 26191 17119
rect 26617 17085 26651 17119
rect 6009 17017 6043 17051
rect 10977 17017 11011 17051
rect 19625 17017 19659 17051
rect 9781 16949 9815 16983
rect 13737 16949 13771 16983
rect 14749 16949 14783 16983
rect 16681 16949 16715 16983
rect 17141 16949 17175 16983
rect 20085 16949 20119 16983
rect 20269 16949 20303 16983
rect 21465 16949 21499 16983
rect 22109 16949 22143 16983
rect 22753 16949 22787 16983
rect 24041 16949 24075 16983
rect 24685 16949 24719 16983
rect 25237 16949 25271 16983
rect 25973 16949 26007 16983
rect 26801 16949 26835 16983
rect 10977 16745 11011 16779
rect 12173 16745 12207 16779
rect 12633 16745 12667 16779
rect 14197 16745 14231 16779
rect 17141 16745 17175 16779
rect 17969 16745 18003 16779
rect 19073 16745 19107 16779
rect 20085 16745 20119 16779
rect 20361 16745 20395 16779
rect 21741 16745 21775 16779
rect 9588 16677 9622 16711
rect 11253 16677 11287 16711
rect 16221 16677 16255 16711
rect 20821 16677 20855 16711
rect 21281 16677 21315 16711
rect 25145 16677 25179 16711
rect 26801 16677 26835 16711
rect 4537 16609 4571 16643
rect 4905 16609 4939 16643
rect 6101 16609 6135 16643
rect 6368 16609 6402 16643
rect 7757 16609 7791 16643
rect 8024 16609 8058 16643
rect 9321 16609 9355 16643
rect 10977 16609 11011 16643
rect 11989 16609 12023 16643
rect 12357 16609 12391 16643
rect 12449 16609 12483 16643
rect 13073 16609 13107 16643
rect 14473 16609 14507 16643
rect 15678 16609 15712 16643
rect 15945 16609 15979 16643
rect 16405 16609 16439 16643
rect 17601 16609 17635 16643
rect 18429 16609 18463 16643
rect 19533 16609 19567 16643
rect 24501 16609 24535 16643
rect 24685 16609 24719 16643
rect 24777 16609 24811 16643
rect 24869 16609 24903 16643
rect 25789 16609 25823 16643
rect 26157 16609 26191 16643
rect 26433 16609 26467 16643
rect 26526 16609 26560 16643
rect 26709 16609 26743 16643
rect 26898 16609 26932 16643
rect 12817 16541 12851 16575
rect 19625 16541 19659 16575
rect 10701 16473 10735 16507
rect 11069 16473 11103 16507
rect 11805 16473 11839 16507
rect 14565 16473 14599 16507
rect 17325 16473 17359 16507
rect 18153 16473 18187 16507
rect 19257 16473 19291 16507
rect 19993 16473 20027 16507
rect 20545 16473 20579 16507
rect 21649 16473 21683 16507
rect 7481 16405 7515 16439
rect 9137 16405 9171 16439
rect 14381 16405 14415 16439
rect 25237 16405 25271 16439
rect 25973 16405 26007 16439
rect 27077 16405 27111 16439
rect 6009 16201 6043 16235
rect 6377 16201 6411 16235
rect 8953 16201 8987 16235
rect 9781 16201 9815 16235
rect 10057 16201 10091 16235
rect 11161 16201 11195 16235
rect 11805 16201 11839 16235
rect 12725 16201 12759 16235
rect 13185 16201 13219 16235
rect 15025 16201 15059 16235
rect 8769 16133 8803 16167
rect 11713 16133 11747 16167
rect 12173 16133 12207 16167
rect 13369 16133 13403 16167
rect 15485 16133 15519 16167
rect 8033 16065 8067 16099
rect 10701 16065 10735 16099
rect 12817 16065 12851 16099
rect 13001 16065 13035 16099
rect 6653 15997 6687 16031
rect 6745 15997 6779 16031
rect 6837 15997 6871 16031
rect 7021 15997 7055 16031
rect 8493 15997 8527 16031
rect 9137 15997 9171 16031
rect 9505 15997 9539 16031
rect 10182 15997 10216 16031
rect 10609 15997 10643 16031
rect 10977 15997 11011 16031
rect 11161 15997 11195 16031
rect 11437 15997 11471 16031
rect 11713 15997 11747 16031
rect 11989 15997 12023 16031
rect 12265 15997 12299 16031
rect 12357 15997 12391 16031
rect 12541 15997 12575 16031
rect 13225 15997 13259 16031
rect 14197 15997 14231 16031
rect 14381 15997 14415 16031
rect 14565 15997 14599 16031
rect 14657 15997 14691 16031
rect 14749 15997 14783 16031
rect 15301 15997 15335 16031
rect 18797 15997 18831 16031
rect 20085 15997 20119 16031
rect 20269 15997 20303 16031
rect 21741 15997 21775 16031
rect 24961 15997 24995 16031
rect 25329 15997 25363 16031
rect 25513 15997 25547 16031
rect 25605 15997 25639 16031
rect 25697 15997 25731 16031
rect 26341 15997 26375 16031
rect 26893 15997 26927 16031
rect 5917 15929 5951 15963
rect 12909 15929 12943 15963
rect 15117 15929 15151 15963
rect 7481 15861 7515 15895
rect 9965 15861 9999 15895
rect 10241 15861 10275 15895
rect 10793 15861 10827 15895
rect 11529 15861 11563 15895
rect 13645 15861 13679 15895
rect 19349 15861 19383 15895
rect 19441 15861 19475 15895
rect 20821 15861 20855 15895
rect 21097 15861 21131 15895
rect 24409 15861 24443 15895
rect 25973 15861 26007 15895
rect 4537 15657 4571 15691
rect 6653 15657 6687 15691
rect 7113 15657 7147 15691
rect 8861 15657 8895 15691
rect 10517 15657 10551 15691
rect 14473 15657 14507 15691
rect 18797 15657 18831 15691
rect 20269 15657 20303 15691
rect 21005 15657 21039 15691
rect 23673 15657 23707 15691
rect 25697 15657 25731 15691
rect 5089 15589 5123 15623
rect 7481 15589 7515 15623
rect 9413 15589 9447 15623
rect 13001 15589 13035 15623
rect 13338 15589 13372 15623
rect 19156 15589 19190 15623
rect 22394 15589 22428 15623
rect 23029 15589 23063 15623
rect 24584 15589 24618 15623
rect 3424 15521 3458 15555
rect 6469 15521 6503 15555
rect 6653 15521 6687 15555
rect 7297 15521 7331 15555
rect 7573 15521 7607 15555
rect 8493 15521 8527 15555
rect 8677 15521 8711 15555
rect 9137 15521 9171 15555
rect 9321 15521 9355 15555
rect 9597 15521 9631 15555
rect 9689 15521 9723 15555
rect 9781 15521 9815 15555
rect 9919 15521 9953 15555
rect 10149 15521 10183 15555
rect 10333 15521 10367 15555
rect 10609 15521 10643 15555
rect 12265 15521 12299 15555
rect 12357 15521 12391 15555
rect 12541 15521 12575 15555
rect 12633 15521 12667 15555
rect 12725 15521 12759 15555
rect 16267 15521 16301 15555
rect 16405 15521 16439 15555
rect 16497 15521 16531 15555
rect 16680 15521 16714 15555
rect 16773 15521 16807 15555
rect 17684 15521 17718 15555
rect 20361 15521 20395 15555
rect 20545 15521 20579 15555
rect 20637 15521 20671 15555
rect 20729 15521 20763 15555
rect 22932 15521 22966 15555
rect 23121 15521 23155 15555
rect 23304 15521 23338 15555
rect 23397 15521 23431 15555
rect 23949 15521 23983 15555
rect 26985 15521 27019 15555
rect 3157 15453 3191 15487
rect 10057 15453 10091 15487
rect 12173 15453 12207 15487
rect 13093 15453 13127 15487
rect 17417 15453 17451 15487
rect 18889 15453 18923 15487
rect 22661 15453 22695 15487
rect 24317 15453 24351 15487
rect 5181 15317 5215 15351
rect 9321 15317 9355 15351
rect 16129 15317 16163 15351
rect 21281 15317 21315 15351
rect 22753 15317 22787 15351
rect 26433 15317 26467 15351
rect 4905 15113 4939 15147
rect 5181 15113 5215 15147
rect 6009 15113 6043 15147
rect 9505 15113 9539 15147
rect 10241 15113 10275 15147
rect 10793 15113 10827 15147
rect 13553 15113 13587 15147
rect 13737 15113 13771 15147
rect 18705 15113 18739 15147
rect 24501 15113 24535 15147
rect 4721 15045 4755 15079
rect 5825 15045 5859 15079
rect 9137 15045 9171 15079
rect 16313 15045 16347 15079
rect 20177 15045 20211 15079
rect 17693 14977 17727 15011
rect 19533 14977 19567 15011
rect 1685 14909 1719 14943
rect 4445 14909 4479 14943
rect 5365 14909 5399 14943
rect 5549 14909 5583 14943
rect 6377 14909 6411 14943
rect 6653 14909 6687 14943
rect 6837 14909 6871 14943
rect 9413 14909 9447 14943
rect 9689 14909 9723 14943
rect 9965 14909 9999 14943
rect 10425 14909 10459 14943
rect 13829 14909 13863 14943
rect 14105 14909 14139 14943
rect 14933 14909 14967 14943
rect 16957 14909 16991 14943
rect 18015 14909 18049 14943
rect 18428 14909 18462 14943
rect 18521 14909 18555 14943
rect 18981 14909 19015 14943
rect 19073 14909 19107 14943
rect 19165 14909 19199 14943
rect 19349 14909 19383 14943
rect 20315 14909 20349 14943
rect 20545 14909 20579 14943
rect 20728 14909 20762 14943
rect 20821 14909 20855 14943
rect 21097 14909 21131 14943
rect 22569 14909 22603 14943
rect 25881 14909 25915 14943
rect 26525 14909 26559 14943
rect 1952 14841 1986 14875
rect 5089 14841 5123 14875
rect 6193 14841 6227 14875
rect 8769 14841 8803 14875
rect 10149 14841 10183 14875
rect 10609 14841 10643 14875
rect 15200 14841 15234 14875
rect 16405 14841 16439 14875
rect 18153 14841 18187 14875
rect 18245 14841 18279 14875
rect 20453 14841 20487 14875
rect 21364 14841 21398 14875
rect 25636 14841 25670 14875
rect 3065 14773 3099 14807
rect 5733 14773 5767 14807
rect 5983 14773 6017 14807
rect 6469 14773 6503 14807
rect 6745 14773 6779 14807
rect 9229 14773 9263 14807
rect 9873 14773 9907 14807
rect 17141 14773 17175 14807
rect 17877 14773 17911 14807
rect 20085 14773 20119 14807
rect 22477 14773 22511 14807
rect 23213 14773 23247 14807
rect 25973 14773 26007 14807
rect 3985 14569 4019 14603
rect 4445 14569 4479 14603
rect 5365 14569 5399 14603
rect 9965 14569 9999 14603
rect 11253 14569 11287 14603
rect 15945 14569 15979 14603
rect 16497 14569 16531 14603
rect 19257 14569 19291 14603
rect 20085 14569 20119 14603
rect 22753 14569 22787 14603
rect 24501 14569 24535 14603
rect 25329 14569 25363 14603
rect 27077 14569 27111 14603
rect 8033 14501 8067 14535
rect 8249 14501 8283 14535
rect 8852 14501 8886 14535
rect 11621 14501 11655 14535
rect 21649 14501 21683 14535
rect 23121 14501 23155 14535
rect 25605 14501 25639 14535
rect 1952 14433 1986 14467
rect 3801 14433 3835 14467
rect 4169 14433 4203 14467
rect 4629 14433 4663 14467
rect 4813 14433 4847 14467
rect 4905 14433 4939 14467
rect 5273 14433 5307 14467
rect 5457 14433 5491 14467
rect 8585 14433 8619 14467
rect 10241 14433 10275 14467
rect 10425 14433 10459 14467
rect 11713 14433 11747 14467
rect 14105 14433 14139 14467
rect 14197 14433 14231 14467
rect 14289 14433 14323 14467
rect 14473 14433 14507 14467
rect 15301 14433 15335 14467
rect 15485 14433 15519 14467
rect 15577 14433 15611 14467
rect 15669 14433 15703 14467
rect 16129 14433 16163 14467
rect 18144 14433 18178 14467
rect 19349 14433 19383 14467
rect 20361 14433 20395 14467
rect 20453 14433 20487 14467
rect 20545 14433 20579 14467
rect 20729 14433 20763 14467
rect 21460 14433 21494 14467
rect 21557 14433 21591 14467
rect 21832 14433 21866 14467
rect 21925 14433 21959 14467
rect 22932 14433 22966 14467
rect 23029 14433 23063 14467
rect 23249 14433 23283 14467
rect 23397 14433 23431 14467
rect 23857 14433 23891 14467
rect 24041 14433 24075 14467
rect 24133 14433 24167 14467
rect 24225 14433 24259 14467
rect 24869 14433 24903 14467
rect 24961 14433 24995 14467
rect 25053 14433 25087 14467
rect 25237 14433 25271 14467
rect 25508 14433 25542 14467
rect 25697 14433 25731 14467
rect 25852 14433 25886 14467
rect 25984 14433 26018 14467
rect 26433 14433 26467 14467
rect 26581 14433 26615 14467
rect 26709 14433 26743 14467
rect 26801 14433 26835 14467
rect 26898 14433 26932 14467
rect 1685 14365 1719 14399
rect 11805 14365 11839 14399
rect 12817 14365 12851 14399
rect 14565 14365 14599 14399
rect 15117 14365 15151 14399
rect 17049 14365 17083 14399
rect 17877 14365 17911 14399
rect 19901 14365 19935 14399
rect 22017 14365 22051 14399
rect 22569 14365 22603 14399
rect 21281 14297 21315 14331
rect 3065 14229 3099 14263
rect 3249 14229 3283 14263
rect 8217 14229 8251 14263
rect 8401 14229 8435 14263
rect 10609 14229 10643 14263
rect 12265 14229 12299 14263
rect 13829 14229 13863 14263
rect 16313 14229 16347 14263
rect 24593 14229 24627 14263
rect 3249 14025 3283 14059
rect 4077 14025 4111 14059
rect 4537 14025 4571 14059
rect 9781 14025 9815 14059
rect 9873 14025 9907 14059
rect 14933 14025 14967 14059
rect 16497 14025 16531 14059
rect 18705 14025 18739 14059
rect 20361 14025 20395 14059
rect 22293 14025 22327 14059
rect 26893 14025 26927 14059
rect 4261 13957 4295 13991
rect 4353 13957 4387 13991
rect 5457 13957 5491 13991
rect 5917 13957 5951 13991
rect 18521 13957 18555 13991
rect 3433 13889 3467 13923
rect 3617 13889 3651 13923
rect 3709 13889 3743 13923
rect 5089 13889 5123 13923
rect 6101 13889 6135 13923
rect 6469 13889 6503 13923
rect 7205 13889 7239 13923
rect 7481 13889 7515 13923
rect 8401 13889 8435 13923
rect 11437 13889 11471 13923
rect 13553 13889 13587 13923
rect 19441 13889 19475 13923
rect 21465 13889 21499 13923
rect 23121 13889 23155 13923
rect 23673 13889 23707 13923
rect 3525 13821 3559 13855
rect 5273 13821 5307 13855
rect 5549 13821 5583 13855
rect 5641 13821 5675 13855
rect 5917 13821 5951 13855
rect 6285 13821 6319 13855
rect 6561 13821 6595 13855
rect 6745 13821 6779 13855
rect 8668 13821 8702 13855
rect 9873 13821 9907 13855
rect 10057 13821 10091 13855
rect 11704 13821 11738 13855
rect 13820 13821 13854 13855
rect 15117 13821 15151 13855
rect 17141 13821 17175 13855
rect 19349 13821 19383 13855
rect 19993 13821 20027 13855
rect 20177 13821 20211 13855
rect 21557 13821 21591 13855
rect 22569 13821 22603 13855
rect 22661 13821 22695 13855
rect 22753 13821 22787 13855
rect 22937 13821 22971 13855
rect 24501 13821 24535 13855
rect 24593 13821 24627 13855
rect 25513 13821 25547 13855
rect 25780 13821 25814 13855
rect 3893 13753 3927 13787
rect 4505 13753 4539 13787
rect 4721 13753 4755 13787
rect 6929 13753 6963 13787
rect 15384 13753 15418 13787
rect 17408 13753 17442 13787
rect 4093 13685 4127 13719
rect 5733 13685 5767 13719
rect 10241 13685 10275 13719
rect 12817 13685 12851 13719
rect 20821 13685 20855 13719
rect 22201 13685 22235 13719
rect 23857 13685 23891 13719
rect 25237 13685 25271 13719
rect 4077 13481 4111 13515
rect 4261 13481 4295 13515
rect 4629 13481 4663 13515
rect 6285 13481 6319 13515
rect 8585 13481 8619 13515
rect 8953 13481 8987 13515
rect 11621 13481 11655 13515
rect 11897 13481 11931 13515
rect 16129 13481 16163 13515
rect 17049 13481 17083 13515
rect 18153 13481 18187 13515
rect 19625 13481 19659 13515
rect 20545 13481 20579 13515
rect 21281 13481 21315 13515
rect 24409 13481 24443 13515
rect 25973 13481 26007 13515
rect 3433 13413 3467 13447
rect 4813 13413 4847 13447
rect 8769 13413 8803 13447
rect 12633 13413 12667 13447
rect 14381 13413 14415 13447
rect 22394 13413 22428 13447
rect 24860 13413 24894 13447
rect 3801 13345 3835 13379
rect 3893 13345 3927 13379
rect 4169 13345 4203 13379
rect 4445 13345 4479 13379
rect 4727 13345 4761 13379
rect 4905 13345 4939 13379
rect 6193 13345 6227 13379
rect 6285 13345 6319 13379
rect 6469 13345 6503 13379
rect 6837 13345 6871 13379
rect 8125 13345 8159 13379
rect 8677 13345 8711 13379
rect 8861 13345 8895 13379
rect 9137 13345 9171 13379
rect 9229 13345 9263 13379
rect 9413 13345 9447 13379
rect 10057 13345 10091 13379
rect 11805 13345 11839 13379
rect 12173 13345 12207 13379
rect 12265 13345 12299 13379
rect 12357 13345 12391 13379
rect 12541 13345 12575 13379
rect 13185 13345 13219 13379
rect 14192 13345 14226 13379
rect 14289 13345 14323 13379
rect 14564 13345 14598 13379
rect 14657 13345 14691 13379
rect 16405 13345 16439 13379
rect 16497 13345 16531 13379
rect 16589 13345 16623 13379
rect 16773 13345 16807 13379
rect 16865 13345 16899 13379
rect 17509 13345 17543 13379
rect 17693 13345 17727 13379
rect 17785 13345 17819 13379
rect 17877 13345 17911 13379
rect 18234 13345 18268 13379
rect 18393 13345 18427 13379
rect 18521 13345 18555 13379
rect 18613 13345 18647 13379
rect 18710 13345 18744 13379
rect 18981 13345 19015 13379
rect 19144 13345 19178 13379
rect 19257 13345 19291 13379
rect 19349 13345 19383 13379
rect 19901 13345 19935 13379
rect 20085 13345 20119 13379
rect 20177 13345 20211 13379
rect 20269 13345 20303 13379
rect 20637 13345 20671 13379
rect 22661 13345 22695 13379
rect 22937 13345 22971 13379
rect 23029 13345 23063 13379
rect 23296 13345 23330 13379
rect 24593 13345 24627 13379
rect 27077 13345 27111 13379
rect 3249 13277 3283 13311
rect 8217 13277 8251 13311
rect 8309 13277 8343 13311
rect 8401 13277 8435 13311
rect 14749 13277 14783 13311
rect 9321 13209 9355 13243
rect 14013 13209 14047 13243
rect 20821 13209 20855 13243
rect 2697 13141 2731 13175
rect 3893 13141 3927 13175
rect 6101 13141 6135 13175
rect 7021 13141 7055 13175
rect 9873 13141 9907 13175
rect 15393 13141 15427 13175
rect 18889 13141 18923 13175
rect 22845 13141 22879 13175
rect 26433 13141 26467 13175
rect 4077 12937 4111 12971
rect 17509 12937 17543 12971
rect 23489 12937 23523 12971
rect 26065 12937 26099 12971
rect 2789 12869 2823 12903
rect 6193 12869 6227 12903
rect 19165 12869 19199 12903
rect 22017 12869 22051 12903
rect 24501 12869 24535 12903
rect 25973 12869 26007 12903
rect 2973 12801 3007 12835
rect 4629 12801 4663 12835
rect 6377 12801 6411 12835
rect 15209 12801 15243 12835
rect 16589 12801 16623 12835
rect 20637 12801 20671 12835
rect 22845 12801 22879 12835
rect 1409 12733 1443 12767
rect 3065 12733 3099 12767
rect 3893 12733 3927 12767
rect 4813 12733 4847 12767
rect 6561 12733 6595 12767
rect 7113 12733 7147 12767
rect 7481 12733 7515 12767
rect 7573 12733 7607 12767
rect 7941 12733 7975 12767
rect 8401 12733 8435 12767
rect 8493 12733 8527 12767
rect 8677 12733 8711 12767
rect 8769 12733 8803 12767
rect 9505 12733 9539 12767
rect 9689 12733 9723 12767
rect 9965 12733 9999 12767
rect 10113 12733 10147 12767
rect 10241 12733 10275 12767
rect 10333 12733 10367 12767
rect 10471 12733 10505 12767
rect 10701 12733 10735 12767
rect 11437 12733 11471 12767
rect 11621 12733 11655 12767
rect 11713 12733 11747 12767
rect 11805 12733 11839 12767
rect 12904 12733 12938 12767
rect 13276 12733 13310 12767
rect 13369 12733 13403 12767
rect 14953 12733 14987 12767
rect 15301 12733 15335 12767
rect 15485 12733 15519 12767
rect 15577 12733 15611 12767
rect 15669 12733 15703 12767
rect 16957 12733 16991 12767
rect 17325 12733 17359 12767
rect 18337 12733 18371 12767
rect 22109 12733 22143 12767
rect 22293 12733 22327 12767
rect 22385 12733 22419 12767
rect 22477 12733 22511 12767
rect 23857 12733 23891 12767
rect 23950 12733 23984 12767
rect 24133 12733 24167 12767
rect 24322 12733 24356 12767
rect 24593 12733 24627 12767
rect 24777 12733 24811 12767
rect 24869 12733 24903 12767
rect 24961 12733 24995 12767
rect 25329 12733 25363 12767
rect 25513 12733 25547 12767
rect 25605 12733 25639 12767
rect 25697 12733 25731 12767
rect 26203 12733 26237 12767
rect 26561 12733 26595 12767
rect 26709 12733 26743 12767
rect 1676 12665 1710 12699
rect 5058 12665 5092 12699
rect 6745 12665 6779 12699
rect 6929 12665 6963 12699
rect 13001 12665 13035 12699
rect 13093 12665 13127 12699
rect 15945 12665 15979 12699
rect 20453 12665 20487 12699
rect 20904 12665 20938 12699
rect 22753 12665 22787 12699
rect 24225 12665 24259 12699
rect 26341 12665 26375 12699
rect 26433 12665 26467 12699
rect 3341 12597 3375 12631
rect 7297 12597 7331 12631
rect 7757 12597 7791 12631
rect 8125 12597 8159 12631
rect 8953 12597 8987 12631
rect 9321 12597 9355 12631
rect 10609 12597 10643 12631
rect 11345 12597 11379 12631
rect 12081 12597 12115 12631
rect 12725 12597 12759 12631
rect 13829 12597 13863 12631
rect 16037 12597 16071 12631
rect 17141 12597 17175 12631
rect 17693 12597 17727 12631
rect 25237 12597 25271 12631
rect 7941 12393 7975 12427
rect 14657 12393 14691 12427
rect 16865 12393 16899 12427
rect 18981 12393 19015 12427
rect 26249 12393 26283 12427
rect 4261 12325 4295 12359
rect 4445 12325 4479 12359
rect 6009 12325 6043 12359
rect 10057 12325 10091 12359
rect 12725 12325 12759 12359
rect 21281 12325 21315 12359
rect 25136 12325 25170 12359
rect 1777 12257 1811 12291
rect 2044 12257 2078 12291
rect 3525 12257 3559 12291
rect 3709 12257 3743 12291
rect 3893 12257 3927 12291
rect 4537 12257 4571 12291
rect 5089 12257 5123 12291
rect 5365 12257 5399 12291
rect 6653 12257 6687 12291
rect 8677 12257 8711 12291
rect 8953 12257 8987 12291
rect 9045 12257 9079 12291
rect 9229 12257 9263 12291
rect 9597 12257 9631 12291
rect 9689 12257 9723 12291
rect 9873 12257 9907 12291
rect 10977 12257 11011 12291
rect 14887 12257 14921 12291
rect 15025 12257 15059 12291
rect 15117 12260 15151 12294
rect 15301 12257 15335 12291
rect 16681 12257 16715 12291
rect 17601 12257 17635 12291
rect 17694 12257 17728 12291
rect 17877 12257 17911 12291
rect 17969 12257 18003 12291
rect 18107 12257 18141 12291
rect 18337 12257 18371 12291
rect 18521 12257 18555 12291
rect 18613 12257 18647 12291
rect 18705 12257 18739 12291
rect 19524 12257 19558 12291
rect 22017 12257 22051 12291
rect 27077 12257 27111 12291
rect 3249 12189 3283 12223
rect 3433 12189 3467 12223
rect 3617 12189 3651 12223
rect 4169 12189 4203 12223
rect 5917 12189 5951 12223
rect 6101 12189 6135 12223
rect 8861 12189 8895 12223
rect 10149 12189 10183 12223
rect 10701 12189 10735 12223
rect 13185 12189 13219 12223
rect 14565 12189 14599 12223
rect 17417 12189 17451 12223
rect 19257 12189 19291 12223
rect 21833 12189 21867 12223
rect 23765 12189 23799 12223
rect 24409 12189 24443 12223
rect 24869 12189 24903 12223
rect 26433 12189 26467 12223
rect 4077 12121 4111 12155
rect 13921 12121 13955 12155
rect 18245 12121 18279 12155
rect 20637 12121 20671 12155
rect 3157 12053 3191 12087
rect 3985 12053 4019 12087
rect 4261 12053 4295 12087
rect 5549 12053 5583 12087
rect 6469 12053 6503 12087
rect 8493 12053 8527 12087
rect 9413 12053 9447 12087
rect 13829 12053 13863 12087
rect 16129 12053 16163 12087
rect 23857 12053 23891 12087
rect 3985 11849 4019 11883
rect 4813 11849 4847 11883
rect 5641 11849 5675 11883
rect 10057 11849 10091 11883
rect 14933 11849 14967 11883
rect 16589 11849 16623 11883
rect 18705 11849 18739 11883
rect 21373 11849 21407 11883
rect 23581 11849 23615 11883
rect 26433 11849 26467 11883
rect 12909 11781 12943 11815
rect 18337 11781 18371 11815
rect 19901 11781 19935 11815
rect 19257 11713 19291 11747
rect 21281 11713 21315 11747
rect 25053 11713 25087 11747
rect 3801 11645 3835 11679
rect 3985 11645 4019 11679
rect 4721 11645 4755 11679
rect 4905 11645 4939 11679
rect 5457 11645 5491 11679
rect 6653 11645 6687 11679
rect 6929 11645 6963 11679
rect 8585 11645 8619 11679
rect 11437 11645 11471 11679
rect 11529 11645 11563 11679
rect 13553 11645 13587 11679
rect 13820 11645 13854 11679
rect 15209 11645 15243 11679
rect 16957 11645 16991 11679
rect 17224 11645 17258 11679
rect 21925 11645 21959 11679
rect 22201 11645 22235 11679
rect 24409 11645 24443 11679
rect 7021 11577 7055 11611
rect 7665 11577 7699 11611
rect 8830 11577 8864 11611
rect 11192 11577 11226 11611
rect 11796 11577 11830 11611
rect 15476 11577 15510 11611
rect 21036 11577 21070 11611
rect 22468 11577 22502 11611
rect 23857 11577 23891 11611
rect 25320 11577 25354 11611
rect 7573 11509 7607 11543
rect 9965 11509 9999 11543
rect 11621 11305 11655 11339
rect 13093 11305 13127 11339
rect 14565 11305 14599 11339
rect 15301 11305 15335 11339
rect 17325 11305 17359 11339
rect 19533 11305 19567 11339
rect 22661 11305 22695 11339
rect 25513 11305 25547 11339
rect 3240 11237 3274 11271
rect 4537 11237 4571 11271
rect 10333 11237 10367 11271
rect 14933 11237 14967 11271
rect 20913 11237 20947 11271
rect 2973 11169 3007 11203
rect 4445 11169 4479 11203
rect 4629 11169 4663 11203
rect 4997 11169 5031 11203
rect 5181 11169 5215 11203
rect 5273 11169 5307 11203
rect 5457 11169 5491 11203
rect 5641 11169 5675 11203
rect 5825 11169 5859 11203
rect 6009 11169 6043 11203
rect 6101 11169 6135 11203
rect 6929 11169 6963 11203
rect 7196 11169 7230 11203
rect 9045 11169 9079 11203
rect 10149 11169 10183 11203
rect 10977 11169 11011 11203
rect 11161 11169 11195 11203
rect 11253 11169 11287 11203
rect 11345 11169 11379 11203
rect 12449 11169 12483 11203
rect 12633 11169 12667 11203
rect 12725 11169 12759 11203
rect 12817 11169 12851 11203
rect 13185 11169 13219 11203
rect 13452 11169 13486 11203
rect 14657 11169 14691 11203
rect 14750 11169 14784 11203
rect 15025 11169 15059 11203
rect 15122 11169 15156 11203
rect 18449 11169 18483 11203
rect 18705 11169 18739 11203
rect 19349 11169 19383 11203
rect 19809 11169 19843 11203
rect 19901 11169 19935 11203
rect 19993 11169 20027 11203
rect 20177 11169 20211 11203
rect 20269 11169 20303 11203
rect 20453 11169 20487 11203
rect 20545 11169 20579 11203
rect 20637 11169 20671 11203
rect 21281 11169 21315 11203
rect 21548 11169 21582 11203
rect 23305 11169 23339 11203
rect 24400 11169 24434 11203
rect 26249 11169 26283 11203
rect 26433 11169 26467 11203
rect 26617 11169 26651 11203
rect 26709 11169 26743 11203
rect 26801 11169 26835 11203
rect 8401 11101 8435 11135
rect 10517 11101 10551 11135
rect 24133 11101 24167 11135
rect 5825 11033 5859 11067
rect 8309 11033 8343 11067
rect 25605 11033 25639 11067
rect 4353 10965 4387 10999
rect 5549 10965 5583 10999
rect 18797 10965 18831 10999
rect 22753 10965 22787 10999
rect 27077 10965 27111 10999
rect 16589 10761 16623 10795
rect 18705 10761 18739 10795
rect 20821 10761 20855 10795
rect 21557 10761 21591 10795
rect 21649 10761 21683 10795
rect 23397 10761 23431 10795
rect 25053 10761 25087 10795
rect 6377 10693 6411 10727
rect 10057 10693 10091 10727
rect 12541 10693 12575 10727
rect 20085 10693 20119 10727
rect 4813 10625 4847 10659
rect 10333 10625 10367 10659
rect 11161 10625 11195 10659
rect 13185 10625 13219 10659
rect 14749 10625 14783 10659
rect 18337 10625 18371 10659
rect 19257 10625 19291 10659
rect 22201 10625 22235 10659
rect 24961 10625 24995 10659
rect 25605 10625 25639 10659
rect 26801 10625 26835 10659
rect 3801 10557 3835 10591
rect 4629 10557 4663 10591
rect 5457 10557 5491 10591
rect 6009 10557 6043 10591
rect 6285 10557 6319 10591
rect 6929 10557 6963 10591
rect 7113 10557 7147 10591
rect 7205 10557 7239 10591
rect 7297 10557 7331 10591
rect 8493 10557 8527 10591
rect 9275 10557 9309 10591
rect 9505 10557 9539 10591
rect 9688 10557 9722 10591
rect 9781 10557 9815 10591
rect 16129 10557 16163 10591
rect 16405 10557 16439 10591
rect 17693 10557 17727 10591
rect 17877 10557 17911 10591
rect 17969 10557 18003 10591
rect 18061 10557 18095 10591
rect 19901 10557 19935 10591
rect 20361 10557 20395 10591
rect 20637 10557 20671 10591
rect 20913 10557 20947 10591
rect 21097 10557 21131 10591
rect 21189 10557 21223 10591
rect 21281 10557 21315 10591
rect 22753 10557 22787 10591
rect 22937 10557 22971 10591
rect 23029 10557 23063 10591
rect 23121 10557 23155 10591
rect 24317 10557 24351 10591
rect 24501 10557 24535 10591
rect 24593 10557 24627 10591
rect 24685 10557 24719 10591
rect 3893 10489 3927 10523
rect 5089 10489 5123 10523
rect 5181 10489 5215 10523
rect 9413 10489 9447 10523
rect 11428 10489 11462 10523
rect 12633 10489 12667 10523
rect 4077 10421 4111 10455
rect 4997 10421 5031 10455
rect 5365 10421 5399 10455
rect 7573 10421 7607 10455
rect 9045 10421 9079 10455
rect 9137 10421 9171 10455
rect 9873 10421 9907 10455
rect 14197 10421 14231 10455
rect 16221 10421 16255 10455
rect 20453 10421 20487 10455
rect 26157 10421 26191 10455
rect 3985 10217 4019 10251
rect 8677 10217 8711 10251
rect 11989 10217 12023 10251
rect 13553 10217 13587 10251
rect 15209 10217 15243 10251
rect 17693 10217 17727 10251
rect 18981 10217 19015 10251
rect 19901 10217 19935 10251
rect 21281 10217 21315 10251
rect 23121 10217 23155 10251
rect 23489 10217 23523 10251
rect 24777 10217 24811 10251
rect 25605 10217 25639 10251
rect 15577 10149 15611 10183
rect 19533 10149 19567 10183
rect 20729 10149 20763 10183
rect 23857 10149 23891 10183
rect 24225 10149 24259 10183
rect 2605 10081 2639 10115
rect 2872 10081 2906 10115
rect 4077 10081 4111 10115
rect 4169 10081 4203 10115
rect 4721 10081 4755 10115
rect 5273 10081 5307 10115
rect 6009 10081 6043 10115
rect 6193 10081 6227 10115
rect 7205 10081 7239 10115
rect 7564 10081 7598 10115
rect 9137 10081 9171 10115
rect 9404 10081 9438 10115
rect 12265 10081 12299 10115
rect 12357 10081 12391 10115
rect 12449 10081 12483 10115
rect 12633 10081 12667 10115
rect 13001 10081 13035 10115
rect 13093 10081 13127 10115
rect 13185 10081 13219 10115
rect 13369 10081 13403 10115
rect 13809 10081 13843 10115
rect 13921 10081 13955 10115
rect 14034 10081 14068 10115
rect 14197 10081 14231 10115
rect 15393 10081 15427 10115
rect 15669 10081 15703 10115
rect 15761 10081 15795 10115
rect 15945 10081 15979 10115
rect 18613 10081 18647 10115
rect 18797 10081 18831 10115
rect 18889 10081 18923 10115
rect 19165 10081 19199 10115
rect 19349 10081 19383 10115
rect 19441 10081 19475 10115
rect 19717 10081 19751 10115
rect 19993 10081 20027 10115
rect 20177 10081 20211 10115
rect 20637 10081 20671 10115
rect 20913 10081 20947 10115
rect 21465 10081 21499 10115
rect 21649 10081 21683 10115
rect 21741 10081 21775 10115
rect 23305 10081 23339 10115
rect 23581 10081 23615 10115
rect 23765 10081 23799 10115
rect 24041 10081 24075 10115
rect 24317 10081 24351 10115
rect 24409 10081 24443 10115
rect 24593 10081 24627 10115
rect 24869 10081 24903 10115
rect 25053 10081 25087 10115
rect 25145 10081 25179 10115
rect 25237 10081 25271 10115
rect 26249 10081 26283 10115
rect 4353 10013 4387 10047
rect 4629 10013 4663 10047
rect 7297 10013 7331 10047
rect 11253 10013 11287 10047
rect 15853 10013 15887 10047
rect 16221 10013 16255 10047
rect 16957 10013 16991 10047
rect 18245 10013 18279 10047
rect 21097 10013 21131 10047
rect 26985 10013 27019 10047
rect 18429 9945 18463 9979
rect 25513 9945 25547 9979
rect 4261 9877 4295 9911
rect 4445 9877 4479 9911
rect 5825 9877 5859 9911
rect 6009 9877 6043 9911
rect 7021 9877 7055 9911
rect 10517 9877 10551 9911
rect 11897 9877 11931 9911
rect 12725 9877 12759 9911
rect 16865 9877 16899 9911
rect 17601 9877 17635 9911
rect 20453 9877 20487 9911
rect 26433 9877 26467 9911
rect 3893 9673 3927 9707
rect 6193 9673 6227 9707
rect 7573 9673 7607 9707
rect 9597 9673 9631 9707
rect 16129 9673 16163 9707
rect 26893 9673 26927 9707
rect 3617 9605 3651 9639
rect 4905 9605 4939 9639
rect 5641 9605 5675 9639
rect 10517 9605 10551 9639
rect 13369 9605 13403 9639
rect 18705 9605 18739 9639
rect 19441 9605 19475 9639
rect 20361 9605 20395 9639
rect 24685 9605 24719 9639
rect 7481 9537 7515 9571
rect 8125 9537 8159 9571
rect 14289 9537 14323 9571
rect 18245 9537 18279 9571
rect 23673 9537 23707 9571
rect 25513 9537 25547 9571
rect 3341 9469 3375 9503
rect 4169 9469 4203 9503
rect 4721 9469 4755 9503
rect 4813 9469 4847 9503
rect 5089 9469 5123 9503
rect 5273 9469 5307 9503
rect 5457 9469 5491 9503
rect 6377 9469 6411 9503
rect 6469 9469 6503 9503
rect 6653 9469 6687 9503
rect 6745 9469 6779 9503
rect 6837 9469 6871 9503
rect 7021 9469 7055 9503
rect 7113 9469 7147 9503
rect 7205 9469 7239 9503
rect 8401 9469 8435 9503
rect 8953 9469 8987 9503
rect 9137 9469 9171 9503
rect 9229 9469 9263 9503
rect 9321 9469 9355 9503
rect 11897 9469 11931 9503
rect 11989 9469 12023 9503
rect 13921 9469 13955 9503
rect 17242 9469 17276 9503
rect 17509 9469 17543 9503
rect 18889 9469 18923 9503
rect 19165 9469 19199 9503
rect 19625 9469 19659 9503
rect 19901 9469 19935 9503
rect 20545 9469 20579 9503
rect 20821 9469 20855 9503
rect 21557 9469 21591 9503
rect 23857 9469 23891 9503
rect 24869 9469 24903 9503
rect 25145 9469 25179 9503
rect 25780 9469 25814 9503
rect 3617 9401 3651 9435
rect 3893 9401 3927 9435
rect 11630 9401 11664 9435
rect 12234 9401 12268 9435
rect 16037 9401 16071 9435
rect 20729 9401 20763 9435
rect 21649 9401 21683 9435
rect 21833 9401 21867 9435
rect 23406 9401 23440 9435
rect 3433 9333 3467 9367
rect 4077 9333 4111 9367
rect 4537 9333 4571 9367
rect 8585 9333 8619 9367
rect 14105 9333 14139 9367
rect 17601 9333 17635 9367
rect 19073 9333 19107 9367
rect 19809 9333 19843 9367
rect 21281 9333 21315 9367
rect 21465 9333 21499 9367
rect 22293 9333 22327 9367
rect 23949 9333 23983 9367
rect 25053 9333 25087 9367
rect 6285 9129 6319 9163
rect 11069 9129 11103 9163
rect 12081 9129 12115 9163
rect 15025 9129 15059 9163
rect 15761 9129 15795 9163
rect 17509 9129 17543 9163
rect 19533 9129 19567 9163
rect 21833 9129 21867 9163
rect 23213 9129 23247 9163
rect 26249 9129 26283 9163
rect 26893 9129 26927 9163
rect 8953 9061 8987 9095
rect 19349 9061 19383 9095
rect 19901 9061 19935 9095
rect 26525 9061 26559 9095
rect 2136 8993 2170 9027
rect 6469 8993 6503 9027
rect 6561 8993 6595 9027
rect 6745 8993 6779 9027
rect 6837 8993 6871 9027
rect 7205 8993 7239 9027
rect 7297 8993 7331 9027
rect 7389 8993 7423 9027
rect 7573 8993 7607 9027
rect 8217 8993 8251 9027
rect 8310 8993 8344 9027
rect 8493 8993 8527 9027
rect 8585 8993 8619 9027
rect 8682 8993 8716 9027
rect 9137 8993 9171 9027
rect 9229 8993 9263 9027
rect 9413 8993 9447 9027
rect 9505 8993 9539 9027
rect 11713 8993 11747 9027
rect 12357 8993 12391 9027
rect 12449 8993 12483 9027
rect 12562 8993 12596 9027
rect 12725 8993 12759 9027
rect 14933 8993 14967 9027
rect 15209 8993 15243 9027
rect 15669 8993 15703 9027
rect 15945 8993 15979 9027
rect 16129 8993 16163 9027
rect 16385 8993 16419 9027
rect 17785 8993 17819 9027
rect 17877 8993 17911 9027
rect 19625 8993 19659 9027
rect 19717 8993 19751 9027
rect 23581 8993 23615 9027
rect 23673 8993 23707 9027
rect 23765 8993 23799 9027
rect 23949 8993 23983 9027
rect 24501 8993 24535 9027
rect 24869 8993 24903 9027
rect 25125 8993 25159 9027
rect 26433 8993 26467 9027
rect 26709 8993 26743 9027
rect 1869 8925 1903 8959
rect 3525 8925 3559 8959
rect 17601 8925 17635 8959
rect 17969 8925 18003 8959
rect 18061 8925 18095 8959
rect 22477 8925 22511 8959
rect 22661 8925 22695 8959
rect 23305 8925 23339 8959
rect 24041 8925 24075 8959
rect 24225 8925 24259 8959
rect 24317 8925 24351 8959
rect 24409 8925 24443 8959
rect 3249 8857 3283 8891
rect 8861 8857 8895 8891
rect 15209 8857 15243 8891
rect 15945 8857 15979 8891
rect 4169 8789 4203 8823
rect 6929 8789 6963 8823
rect 3985 8585 4019 8619
rect 7665 8585 7699 8619
rect 11989 8585 12023 8619
rect 16589 8585 16623 8619
rect 18337 8585 18371 8619
rect 20085 8585 20119 8619
rect 20177 8585 20211 8619
rect 22293 8585 22327 8619
rect 23581 8585 23615 8619
rect 23949 8585 23983 8619
rect 24501 8585 24535 8619
rect 25145 8585 25179 8619
rect 25421 8585 25455 8619
rect 4537 8517 4571 8551
rect 6837 8517 6871 8551
rect 10701 8517 10735 8551
rect 16681 8517 16715 8551
rect 17969 8517 18003 8551
rect 24685 8517 24719 8551
rect 25605 8517 25639 8551
rect 4353 8449 4387 8483
rect 4445 8449 4479 8483
rect 4905 8449 4939 8483
rect 7021 8449 7055 8483
rect 16497 8449 16531 8483
rect 18705 8449 18739 8483
rect 21741 8449 21775 8483
rect 22385 8457 22419 8491
rect 23949 8449 23983 8483
rect 1593 8381 1627 8415
rect 3893 8381 3927 8415
rect 4169 8381 4203 8415
rect 4721 8381 4755 8415
rect 5457 8381 5491 8415
rect 5724 8381 5758 8415
rect 8769 8381 8803 8415
rect 8953 8381 8987 8415
rect 9045 8381 9079 8415
rect 9137 8381 9171 8415
rect 10885 8381 10919 8415
rect 10977 8381 11011 8415
rect 11161 8381 11195 8415
rect 11253 8381 11287 8415
rect 11345 8381 11379 8415
rect 11493 8381 11527 8415
rect 11810 8381 11844 8415
rect 12909 8381 12943 8415
rect 13553 8381 13587 8415
rect 13737 8381 13771 8415
rect 13829 8381 13863 8415
rect 13921 8381 13955 8415
rect 16405 8381 16439 8415
rect 16773 8381 16807 8415
rect 21557 8381 21591 8415
rect 22569 8381 22603 8415
rect 22661 8381 22695 8415
rect 23029 8381 23063 8415
rect 23857 8381 23891 8415
rect 24961 8381 24995 8415
rect 25697 8381 25731 8415
rect 1860 8313 1894 8347
rect 11621 8313 11655 8347
rect 11713 8313 11747 8347
rect 18950 8313 18984 8347
rect 21290 8313 21324 8347
rect 24317 8313 24351 8347
rect 24517 8313 24551 8347
rect 24777 8313 24811 8347
rect 25237 8313 25271 8347
rect 25437 8313 25471 8347
rect 2973 8245 3007 8279
rect 3249 8245 3283 8279
rect 9413 8245 9447 8279
rect 12357 8245 12391 8279
rect 14197 8245 14231 8279
rect 15761 8245 15795 8279
rect 18337 8245 18371 8279
rect 18521 8245 18555 8279
rect 22385 8245 22419 8279
rect 24225 8245 24259 8279
rect 25881 8245 25915 8279
rect 2605 8041 2639 8075
rect 2789 8041 2823 8075
rect 12909 8041 12943 8075
rect 13645 8041 13679 8075
rect 18797 8041 18831 8075
rect 22201 8041 22235 8075
rect 24133 8041 24167 8075
rect 24869 8041 24903 8075
rect 3249 7973 3283 8007
rect 13277 7973 13311 8007
rect 13369 7973 13403 8007
rect 14381 7973 14415 8007
rect 20821 7973 20855 8007
rect 20913 7973 20947 8007
rect 22017 7973 22051 8007
rect 24317 7973 24351 8007
rect 2513 7905 2547 7939
rect 2697 7905 2731 7939
rect 2973 7905 3007 7939
rect 3157 7905 3191 7939
rect 3525 7905 3559 7939
rect 3985 7905 4019 7939
rect 4077 7905 4111 7939
rect 4261 7905 4295 7939
rect 6460 7905 6494 7939
rect 8401 7905 8435 7939
rect 8493 7905 8527 7939
rect 8585 7905 8619 7939
rect 8769 7905 8803 7939
rect 8861 7905 8895 7939
rect 9128 7905 9162 7939
rect 11529 7905 11563 7939
rect 11796 7905 11830 7939
rect 12990 7905 13024 7939
rect 13094 7905 13128 7939
rect 13466 7905 13500 7939
rect 14479 7905 14513 7939
rect 14657 7905 14691 7939
rect 14749 7905 14783 7939
rect 14841 7905 14875 7939
rect 15215 7905 15249 7939
rect 15393 7905 15427 7939
rect 15485 7905 15519 7939
rect 15577 7905 15611 7939
rect 16129 7905 16163 7939
rect 16385 7905 16419 7939
rect 18613 7905 18647 7939
rect 19441 7905 19475 7939
rect 19533 7905 19567 7939
rect 19717 7905 19751 7939
rect 20545 7905 20579 7939
rect 20637 7905 20671 7939
rect 21005 7905 21039 7939
rect 21465 7905 21499 7939
rect 21649 7905 21683 7939
rect 21741 7905 21775 7939
rect 21833 7905 21867 7939
rect 22293 7905 22327 7939
rect 23029 7905 23063 7939
rect 23673 7905 23707 7939
rect 23857 7905 23891 7939
rect 24225 7905 24259 7939
rect 24409 7895 24443 7929
rect 24685 7905 24719 7939
rect 25145 7905 25179 7939
rect 25237 7905 25271 7939
rect 3249 7837 3283 7871
rect 6193 7837 6227 7871
rect 13737 7837 13771 7871
rect 15853 7837 15887 7871
rect 19257 7837 19291 7871
rect 19625 7837 19659 7871
rect 21097 7837 21131 7871
rect 22385 7837 22419 7871
rect 24133 7837 24167 7871
rect 21281 7769 21315 7803
rect 23949 7769 23983 7803
rect 3433 7701 3467 7735
rect 4261 7701 4295 7735
rect 7573 7701 7607 7735
rect 8125 7701 8159 7735
rect 10241 7701 10275 7735
rect 15117 7701 15151 7735
rect 17509 7701 17543 7735
rect 22017 7701 22051 7735
rect 23121 7701 23155 7735
rect 24961 7701 24995 7735
rect 3985 7497 4019 7531
rect 5365 7497 5399 7531
rect 5733 7497 5767 7531
rect 6469 7497 6503 7531
rect 11897 7497 11931 7531
rect 13369 7497 13403 7531
rect 13553 7497 13587 7531
rect 16681 7497 16715 7531
rect 18981 7497 19015 7531
rect 20269 7497 20303 7531
rect 23029 7497 23063 7531
rect 24409 7497 24443 7531
rect 26893 7497 26927 7531
rect 11161 7429 11195 7463
rect 20729 7429 20763 7463
rect 22845 7429 22879 7463
rect 3341 7361 3375 7395
rect 7021 7361 7055 7395
rect 7757 7361 7791 7395
rect 8861 7361 8895 7395
rect 17877 7361 17911 7395
rect 19349 7361 19383 7395
rect 24041 7361 24075 7395
rect 25513 7361 25547 7395
rect 2881 7293 2915 7327
rect 3065 7293 3099 7327
rect 3525 7293 3559 7327
rect 3617 7293 3651 7327
rect 3709 7293 3743 7327
rect 3801 7293 3835 7327
rect 4629 7293 4663 7327
rect 4997 7293 5031 7327
rect 6009 7293 6043 7327
rect 6101 7293 6135 7327
rect 6193 7293 6227 7327
rect 6377 7293 6411 7327
rect 9117 7293 9151 7327
rect 10609 7293 10643 7327
rect 10701 7293 10735 7327
rect 10885 7293 10919 7327
rect 10977 7293 11011 7327
rect 11253 7293 11287 7327
rect 11437 7293 11471 7327
rect 11529 7293 11563 7327
rect 11621 7293 11655 7327
rect 12725 7293 12759 7327
rect 12873 7293 12907 7327
rect 13093 7293 13127 7327
rect 13190 7293 13224 7327
rect 14666 7293 14700 7327
rect 14933 7293 14967 7327
rect 15117 7293 15151 7327
rect 16865 7293 16899 7327
rect 17601 7293 17635 7327
rect 18797 7293 18831 7327
rect 20637 7293 20671 7327
rect 20821 7293 20855 7327
rect 21465 7293 21499 7327
rect 21732 7293 21766 7327
rect 22937 7293 22971 7327
rect 23121 7293 23155 7327
rect 23949 7293 23983 7327
rect 24133 7293 24167 7327
rect 25421 7293 25455 7327
rect 25780 7293 25814 7327
rect 5365 7225 5399 7259
rect 13001 7225 13035 7259
rect 15384 7225 15418 7259
rect 20177 7225 20211 7259
rect 24393 7225 24427 7259
rect 24593 7225 24627 7259
rect 2973 7157 3007 7191
rect 5549 7157 5583 7191
rect 7205 7157 7239 7191
rect 10241 7157 10275 7191
rect 16497 7157 16531 7191
rect 19993 7157 20027 7191
rect 24225 7157 24259 7191
rect 24777 7157 24811 7191
rect 3893 6953 3927 6987
rect 8217 6953 8251 6987
rect 11529 6953 11563 6987
rect 12173 6953 12207 6987
rect 24041 6953 24075 6987
rect 25881 6953 25915 6987
rect 6193 6885 6227 6919
rect 8493 6885 8527 6919
rect 9749 6885 9783 6919
rect 9965 6885 9999 6919
rect 13001 6885 13035 6919
rect 20729 6885 20763 6919
rect 23857 6885 23891 6919
rect 2513 6817 2547 6851
rect 2780 6817 2814 6851
rect 4169 6817 4203 6851
rect 4436 6817 4470 6851
rect 7849 6817 7883 6851
rect 8396 6817 8430 6851
rect 8585 6817 8619 6851
rect 8713 6817 8747 6851
rect 8861 6817 8895 6851
rect 9137 6817 9171 6851
rect 9229 6817 9263 6851
rect 9413 6817 9447 6851
rect 9505 6817 9539 6851
rect 10057 6817 10091 6851
rect 10977 6817 11011 6851
rect 11069 6817 11103 6851
rect 11253 6817 11287 6851
rect 11345 6817 11379 6851
rect 12265 6817 12299 6851
rect 17868 6817 17902 6851
rect 19073 6817 19107 6851
rect 19809 6817 19843 6851
rect 19993 6817 20027 6851
rect 20269 6817 20303 6851
rect 20821 6817 20855 6851
rect 20913 6817 20947 6851
rect 21097 6817 21131 6851
rect 21741 6817 21775 6851
rect 24133 6817 24167 6851
rect 24225 6817 24259 6851
rect 24409 6817 24443 6851
rect 24501 6817 24535 6851
rect 24768 6817 24802 6851
rect 26157 6817 26191 6851
rect 26433 6817 26467 6851
rect 10333 6749 10367 6783
rect 12449 6749 12483 6783
rect 13093 6749 13127 6783
rect 13277 6749 13311 6783
rect 17601 6749 17635 6783
rect 19625 6749 19659 6783
rect 20177 6749 20211 6783
rect 26985 6749 27019 6783
rect 8953 6681 8987 6715
rect 9597 6681 9631 6715
rect 11805 6681 11839 6715
rect 20361 6681 20395 6715
rect 26065 6681 26099 6715
rect 5549 6613 5583 6647
rect 9781 6613 9815 6647
rect 10149 6613 10183 6647
rect 10241 6613 10275 6647
rect 12633 6613 12667 6647
rect 18981 6613 19015 6647
rect 20545 6613 20579 6647
rect 23029 6613 23063 6647
rect 4997 6409 5031 6443
rect 5825 6409 5859 6443
rect 9413 6409 9447 6443
rect 10333 6409 10367 6443
rect 11253 6409 11287 6443
rect 17693 6409 17727 6443
rect 18521 6409 18555 6443
rect 23489 6409 23523 6443
rect 23581 6409 23615 6443
rect 24133 6409 24167 6443
rect 25881 6409 25915 6443
rect 5549 6341 5583 6375
rect 10977 6341 11011 6375
rect 20729 6341 20763 6375
rect 6101 6273 6135 6307
rect 6285 6273 6319 6307
rect 6561 6273 6595 6307
rect 11069 6273 11103 6307
rect 18705 6273 18739 6307
rect 20637 6273 20671 6307
rect 23397 6273 23431 6307
rect 24501 6273 24535 6307
rect 5181 6205 5215 6239
rect 6009 6205 6043 6239
rect 6193 6205 6227 6239
rect 8033 6205 8067 6239
rect 8217 6205 8251 6239
rect 8493 6205 8527 6239
rect 8677 6205 8711 6239
rect 8861 6205 8895 6239
rect 9689 6205 9723 6239
rect 10425 6205 10459 6239
rect 11345 6205 11379 6239
rect 11437 6205 11471 6239
rect 11621 6205 11655 6239
rect 13737 6205 13771 6239
rect 14105 6205 14139 6239
rect 16129 6205 16163 6239
rect 18061 6205 18095 6239
rect 18429 6205 18463 6239
rect 18521 6205 18555 6239
rect 20453 6205 20487 6239
rect 20821 6205 20855 6239
rect 20913 6205 20947 6239
rect 22385 6205 22419 6239
rect 23673 6205 23707 6239
rect 24041 6205 24075 6239
rect 24317 6205 24351 6239
rect 6828 6137 6862 6171
rect 8125 6137 8159 6171
rect 10609 6137 10643 6171
rect 10701 6137 10735 6171
rect 11069 6137 11103 6171
rect 13921 6137 13955 6171
rect 14013 6137 14047 6171
rect 17509 6137 17543 6171
rect 17725 6137 17759 6171
rect 18153 6137 18187 6171
rect 18245 6137 18279 6171
rect 22140 6137 22174 6171
rect 23949 6137 23983 6171
rect 24409 6137 24443 6171
rect 24768 6137 24802 6171
rect 5273 6069 5307 6103
rect 5365 6069 5399 6103
rect 7941 6069 7975 6103
rect 8585 6069 8619 6103
rect 10793 6069 10827 6103
rect 11529 6069 11563 6103
rect 14289 6069 14323 6103
rect 15945 6069 15979 6103
rect 17877 6069 17911 6103
rect 21005 6069 21039 6103
rect 5825 5865 5859 5899
rect 7757 5865 7791 5899
rect 9505 5865 9539 5899
rect 11621 5865 11655 5899
rect 12081 5865 12115 5899
rect 12265 5865 12299 5899
rect 13093 5865 13127 5899
rect 13921 5865 13955 5899
rect 14749 5865 14783 5899
rect 15117 5865 15151 5899
rect 19257 5865 19291 5899
rect 20269 5865 20303 5899
rect 21373 5865 21407 5899
rect 22109 5865 22143 5899
rect 22753 5865 22787 5899
rect 25053 5865 25087 5899
rect 8585 5797 8619 5831
rect 10793 5797 10827 5831
rect 19625 5797 19659 5831
rect 20729 5797 20763 5831
rect 25697 5797 25731 5831
rect 3985 5729 4019 5763
rect 4077 5729 4111 5763
rect 4169 5729 4203 5763
rect 4353 5729 4387 5763
rect 5365 5729 5399 5763
rect 6009 5729 6043 5763
rect 7481 5729 7515 5763
rect 7849 5729 7883 5763
rect 8769 5729 8803 5763
rect 8953 5729 8987 5763
rect 10977 5729 11011 5763
rect 11897 5729 11931 5763
rect 12173 5729 12207 5763
rect 12633 5729 12667 5763
rect 13461 5729 13495 5763
rect 13553 5729 13587 5763
rect 14289 5729 14323 5763
rect 16313 5729 16347 5763
rect 16497 5729 16531 5763
rect 16589 5729 16623 5763
rect 18052 5729 18086 5763
rect 19441 5729 19475 5763
rect 19901 5729 19935 5763
rect 20085 5729 20119 5763
rect 20361 5729 20395 5763
rect 22937 5729 22971 5763
rect 24133 5729 24167 5763
rect 24409 5729 24443 5763
rect 25329 5729 25363 5763
rect 25513 5729 25547 5763
rect 25605 5729 25639 5763
rect 25789 5729 25823 5763
rect 4445 5661 4479 5695
rect 4997 5661 5031 5695
rect 7573 5661 7607 5695
rect 7757 5661 7791 5695
rect 8493 5661 8527 5695
rect 12725 5661 12759 5695
rect 12909 5661 12943 5695
rect 13737 5661 13771 5695
rect 14381 5661 14415 5695
rect 14473 5661 14507 5695
rect 15209 5661 15243 5695
rect 15301 5661 15335 5695
rect 16129 5661 16163 5695
rect 17785 5661 17819 5695
rect 21925 5661 21959 5695
rect 22293 5661 22327 5695
rect 22385 5661 22419 5695
rect 22477 5661 22511 5695
rect 22569 5661 22603 5695
rect 23949 5661 23983 5695
rect 19165 5593 19199 5627
rect 20913 5593 20947 5627
rect 3709 5525 3743 5559
rect 5549 5525 5583 5559
rect 11713 5525 11747 5559
rect 16773 5525 16807 5559
rect 20729 5525 20763 5559
rect 24317 5525 24351 5559
rect 25145 5525 25179 5559
rect 7021 5321 7055 5355
rect 9873 5321 9907 5355
rect 10057 5321 10091 5355
rect 13553 5321 13587 5355
rect 14565 5321 14599 5355
rect 15117 5321 15151 5355
rect 18245 5321 18279 5355
rect 21833 5321 21867 5355
rect 23581 5321 23615 5355
rect 25237 5321 25271 5355
rect 26709 5321 26743 5355
rect 4169 5185 4203 5219
rect 14197 5185 14231 5219
rect 15669 5185 15703 5219
rect 23397 5185 23431 5219
rect 23857 5185 23891 5219
rect 6193 5117 6227 5151
rect 7205 5117 7239 5151
rect 7389 5117 7423 5151
rect 7481 5117 7515 5151
rect 7757 5117 7791 5151
rect 8033 5117 8067 5151
rect 8493 5117 8527 5151
rect 11437 5117 11471 5151
rect 12725 5117 12759 5151
rect 14381 5117 14415 5151
rect 15485 5117 15519 5151
rect 15577 5117 15611 5151
rect 16589 5117 16623 5151
rect 16856 5117 16890 5151
rect 18429 5117 18463 5151
rect 19901 5117 19935 5151
rect 20085 5117 20119 5151
rect 20453 5117 20487 5151
rect 23121 5117 23155 5151
rect 23305 5117 23339 5151
rect 23673 5117 23707 5151
rect 25329 5117 25363 5151
rect 4436 5049 4470 5083
rect 7573 5049 7607 5083
rect 7941 5049 7975 5083
rect 8738 5049 8772 5083
rect 11192 5049 11226 5083
rect 14013 5049 14047 5083
rect 19993 5049 20027 5083
rect 20698 5049 20732 5083
rect 23397 5049 23431 5083
rect 24102 5049 24136 5083
rect 25574 5049 25608 5083
rect 5549 4981 5583 5015
rect 5641 4981 5675 5015
rect 12173 4981 12207 5015
rect 13921 4981 13955 5015
rect 17969 4981 18003 5015
rect 23213 4981 23247 5015
rect 4445 4777 4479 4811
rect 4721 4777 4755 4811
rect 7941 4777 7975 4811
rect 8493 4777 8527 4811
rect 12357 4777 12391 4811
rect 12817 4777 12851 4811
rect 13829 4777 13863 4811
rect 14657 4777 14691 4811
rect 23765 4777 23799 4811
rect 24793 4777 24827 4811
rect 24961 4777 24995 4811
rect 25237 4777 25271 4811
rect 15025 4709 15059 4743
rect 16405 4709 16439 4743
rect 17049 4709 17083 4743
rect 17141 4709 17175 4743
rect 24593 4709 24627 4743
rect 3065 4641 3099 4675
rect 3332 4641 3366 4675
rect 4997 4641 5031 4675
rect 5089 4641 5123 4675
rect 5181 4641 5215 4675
rect 5365 4641 5399 4675
rect 7757 4641 7791 4675
rect 8033 4641 8067 4675
rect 8309 4641 8343 4675
rect 8585 4641 8619 4675
rect 10425 4641 10459 4675
rect 10517 4641 10551 4675
rect 10609 4641 10643 4675
rect 10793 4641 10827 4675
rect 10977 4641 11011 4675
rect 11244 4641 11278 4675
rect 12633 4641 12667 4675
rect 12909 4641 12943 4675
rect 14197 4641 14231 4675
rect 15117 4641 15151 4675
rect 16221 4641 16255 4675
rect 16497 4641 16531 4675
rect 16589 4641 16623 4675
rect 16865 4641 16899 4675
rect 17233 4641 17267 4675
rect 18797 4641 18831 4675
rect 24409 4641 24443 4675
rect 25053 4641 25087 4675
rect 14289 4573 14323 4607
rect 14473 4573 14507 4607
rect 15209 4573 15243 4607
rect 18613 4573 18647 4607
rect 8125 4505 8159 4539
rect 17417 4505 17451 4539
rect 7573 4437 7607 4471
rect 10149 4437 10183 4471
rect 12449 4437 12483 4471
rect 16773 4437 16807 4471
rect 18981 4437 19015 4471
rect 24777 4437 24811 4471
rect 10057 4233 10091 4267
rect 12173 4233 12207 4267
rect 19625 4233 19659 4267
rect 3065 4165 3099 4199
rect 12265 4097 12299 4131
rect 13553 4097 13587 4131
rect 18705 4097 18739 4131
rect 21005 4097 21039 4131
rect 1685 4029 1719 4063
rect 3617 4029 3651 4063
rect 3801 4029 3835 4063
rect 4077 4029 4111 4063
rect 4445 4029 4479 4063
rect 4721 4029 4755 4063
rect 4813 4029 4847 4063
rect 4905 4029 4939 4063
rect 5089 4029 5123 4063
rect 6653 4029 6687 4063
rect 6745 4029 6779 4063
rect 6837 4029 6871 4063
rect 7021 4029 7055 4063
rect 7665 4029 7699 4063
rect 8401 4029 8435 4063
rect 8677 4029 8711 4063
rect 10701 4029 10735 4063
rect 10793 4029 10827 4063
rect 10977 4029 11011 4063
rect 11072 4029 11106 4063
rect 11207 4029 11241 4063
rect 11529 4029 11563 4063
rect 11713 4029 11747 4063
rect 11805 4029 11839 4063
rect 11897 4029 11931 4063
rect 12817 4029 12851 4063
rect 13737 4029 13771 4063
rect 14013 4029 14047 4063
rect 16681 4029 16715 4063
rect 16865 4029 16899 4063
rect 17049 4029 17083 4063
rect 17325 4029 17359 4063
rect 17509 4029 17543 4063
rect 17693 4029 17727 4063
rect 17877 4029 17911 4063
rect 18889 4029 18923 4063
rect 19349 4029 19383 4063
rect 23949 4029 23983 4063
rect 1952 3961 1986 3995
rect 4169 3961 4203 3995
rect 4261 3961 4295 3995
rect 5365 3961 5399 3995
rect 7113 3961 7147 3995
rect 8493 3961 8527 3995
rect 16957 3961 16991 3995
rect 20738 3961 20772 3995
rect 24133 3961 24167 3995
rect 3433 3893 3467 3927
rect 3893 3893 3927 3927
rect 4537 3893 4571 3927
rect 5273 3893 5307 3927
rect 6377 3893 6411 3927
rect 8861 3893 8895 3927
rect 11437 3893 11471 3927
rect 13921 3893 13955 3927
rect 17233 3893 17267 3927
rect 18061 3893 18095 3927
rect 19073 3893 19107 3927
rect 19533 3893 19567 3927
rect 2789 3689 2823 3723
rect 10793 3689 10827 3723
rect 12357 3689 12391 3723
rect 13185 3689 13219 3723
rect 13553 3689 13587 3723
rect 15209 3689 15243 3723
rect 16129 3689 16163 3723
rect 16497 3689 16531 3723
rect 19533 3689 19567 3723
rect 19625 3689 19659 3723
rect 6184 3621 6218 3655
rect 11244 3621 11278 3655
rect 14381 3621 14415 3655
rect 15577 3621 15611 3655
rect 18398 3621 18432 3655
rect 2973 3553 3007 3587
rect 3985 3553 4019 3587
rect 4261 3553 4295 3587
rect 4528 3553 4562 3587
rect 5917 3553 5951 3587
rect 8881 3553 8915 3587
rect 9137 3553 9171 3587
rect 9413 3553 9447 3587
rect 9680 3553 9714 3587
rect 10977 3553 11011 3587
rect 12633 3553 12667 3587
rect 12725 3553 12759 3587
rect 12817 3553 12851 3587
rect 13001 3553 13035 3587
rect 16957 3553 16991 3587
rect 17141 3553 17175 3587
rect 17233 3553 17267 3587
rect 17325 3553 17359 3587
rect 17877 3553 17911 3587
rect 20738 3553 20772 3587
rect 21005 3553 21039 3587
rect 4169 3485 4203 3519
rect 13645 3485 13679 3519
rect 13829 3485 13863 3519
rect 14197 3485 14231 3519
rect 14289 3485 14323 3519
rect 15669 3485 15703 3519
rect 15853 3485 15887 3519
rect 16589 3485 16623 3519
rect 16773 3485 16807 3519
rect 17693 3485 17727 3519
rect 18153 3485 18187 3519
rect 14749 3417 14783 3451
rect 17509 3417 17543 3451
rect 3801 3349 3835 3383
rect 5641 3349 5675 3383
rect 7297 3349 7331 3383
rect 7757 3349 7791 3383
rect 12449 3349 12483 3383
rect 18061 3349 18095 3383
rect 4629 3145 4663 3179
rect 6653 3145 6687 3179
rect 9137 3145 9171 3179
rect 12449 3145 12483 3179
rect 13553 3145 13587 3179
rect 20177 3145 20211 3179
rect 20453 3145 20487 3179
rect 7665 3077 7699 3111
rect 3249 3009 3283 3043
rect 5917 3009 5951 3043
rect 8401 3009 8435 3043
rect 10241 3009 10275 3043
rect 14197 3009 14231 3043
rect 18797 3009 18831 3043
rect 5365 2941 5399 2975
rect 5457 2941 5491 2975
rect 5733 2941 5767 2975
rect 6561 2941 6595 2975
rect 6929 2941 6963 2975
rect 7021 2941 7055 2975
rect 7113 2941 7147 2975
rect 7297 2941 7331 2975
rect 7849 2941 7883 2975
rect 7941 2941 7975 2975
rect 8217 2941 8251 2975
rect 9045 2941 9079 2975
rect 9413 2941 9447 2975
rect 9505 2941 9539 2975
rect 9597 2941 9631 2975
rect 9781 2941 9815 2975
rect 10057 2941 10091 2975
rect 10885 2941 10919 2975
rect 10977 2941 11011 2975
rect 11253 2941 11287 2975
rect 11897 2941 11931 2975
rect 12173 2941 12207 2975
rect 12289 2941 12323 2975
rect 13921 2941 13955 2975
rect 15853 2941 15887 2975
rect 16221 2941 16255 2975
rect 16497 2941 16531 2975
rect 16773 2941 16807 2975
rect 16865 2941 16899 2975
rect 18337 2941 18371 2975
rect 20269 2941 20303 2975
rect 3516 2873 3550 2907
rect 5549 2873 5583 2907
rect 8033 2873 8067 2907
rect 11069 2873 11103 2907
rect 12081 2873 12115 2907
rect 14013 2873 14047 2907
rect 14749 2873 14783 2907
rect 16037 2873 16071 2907
rect 16129 2873 16163 2907
rect 16681 2873 16715 2907
rect 19042 2873 19076 2907
rect 5181 2805 5215 2839
rect 9873 2805 9907 2839
rect 10701 2805 10735 2839
rect 14473 2805 14507 2839
rect 16405 2805 16439 2839
rect 17049 2805 17083 2839
rect 18521 2805 18555 2839
rect 3709 2601 3743 2635
rect 14197 2601 14231 2635
rect 14657 2601 14691 2635
rect 6469 2533 6503 2567
rect 6561 2533 6595 2567
rect 15669 2533 15703 2567
rect 16681 2533 16715 2567
rect 3893 2465 3927 2499
rect 5181 2465 5215 2499
rect 5365 2465 5399 2499
rect 6377 2465 6411 2499
rect 6745 2465 6779 2499
rect 7481 2465 7515 2499
rect 7849 2465 7883 2499
rect 8033 2465 8067 2499
rect 8677 2465 8711 2499
rect 10517 2465 10551 2499
rect 11621 2465 11655 2499
rect 12449 2465 12483 2499
rect 14289 2465 14323 2499
rect 16405 2465 16439 2499
rect 16497 2465 16531 2499
rect 16957 2465 16991 2499
rect 17141 2465 17175 2499
rect 17233 2465 17267 2499
rect 17509 2465 17543 2499
rect 19809 2465 19843 2499
rect 19993 2465 20027 2499
rect 20361 2465 20395 2499
rect 6837 2397 6871 2431
rect 7573 2397 7607 2431
rect 10701 2397 10735 2431
rect 11805 2397 11839 2431
rect 12265 2397 12299 2431
rect 12633 2397 12667 2431
rect 14105 2397 14139 2431
rect 16773 2397 16807 2431
rect 20545 2397 20579 2431
rect 21005 2397 21039 2431
rect 4997 2261 5031 2295
rect 6193 2261 6227 2295
rect 8493 2261 8527 2295
rect 10333 2261 10367 2295
rect 11437 2261 11471 2295
rect 15577 2261 15611 2295
rect 17417 2261 17451 2295
rect 17693 2261 17727 2295
rect 9781 2057 9815 2091
rect 5917 1989 5951 2023
rect 14381 1989 14415 2023
rect 16313 1989 16347 2023
rect 7665 1921 7699 1955
rect 19441 1921 19475 1955
rect 20729 1921 20763 1955
rect 4537 1853 4571 1887
rect 6193 1853 6227 1887
rect 6377 1853 6411 1887
rect 6561 1853 6595 1887
rect 6837 1853 6871 1887
rect 7573 1853 7607 1887
rect 7941 1853 7975 1887
rect 8125 1853 8159 1887
rect 8401 1853 8435 1887
rect 10425 1853 10459 1887
rect 11529 1853 11563 1887
rect 12633 1853 12667 1887
rect 13829 1853 13863 1887
rect 14013 1853 14047 1887
rect 14197 1853 14231 1887
rect 14473 1853 14507 1887
rect 14657 1853 14691 1887
rect 14841 1853 14875 1887
rect 14933 1853 14967 1887
rect 15761 1853 15795 1887
rect 15945 1853 15979 1887
rect 16134 1853 16168 1887
rect 17794 1853 17828 1887
rect 18061 1853 18095 1887
rect 18981 1853 19015 1887
rect 19165 1853 19199 1887
rect 19533 1853 19567 1887
rect 20269 1853 20303 1887
rect 20453 1853 20487 1887
rect 20821 1853 20855 1887
rect 4804 1785 4838 1819
rect 6929 1785 6963 1819
rect 8646 1785 8680 1819
rect 14105 1785 14139 1819
rect 16037 1785 16071 1819
rect 20177 1785 20211 1819
rect 6653 1717 6687 1751
rect 10241 1717 10275 1751
rect 11345 1717 11379 1751
rect 12817 1717 12851 1751
rect 15117 1717 15151 1751
rect 16681 1717 16715 1751
rect 21373 1717 21407 1751
rect 4905 1513 4939 1547
rect 7205 1513 7239 1547
rect 10793 1513 10827 1547
rect 12357 1513 12391 1547
rect 13921 1513 13955 1547
rect 16313 1513 16347 1547
rect 6092 1445 6126 1479
rect 9680 1445 9714 1479
rect 11244 1445 11278 1479
rect 12808 1445 12842 1479
rect 15126 1445 15160 1479
rect 17448 1445 17482 1479
rect 5089 1377 5123 1411
rect 7941 1377 7975 1411
rect 8585 1377 8619 1411
rect 8953 1377 8987 1411
rect 15485 1377 15519 1411
rect 17785 1377 17819 1411
rect 17969 1377 18003 1411
rect 18061 1377 18095 1411
rect 18158 1377 18192 1411
rect 19073 1377 19107 1411
rect 19257 1377 19291 1411
rect 19349 1377 19383 1411
rect 19493 1377 19527 1411
rect 19809 1377 19843 1411
rect 19993 1377 20027 1411
rect 20361 1377 20395 1411
rect 20545 1377 20579 1411
rect 21005 1377 21039 1411
rect 5825 1309 5859 1343
rect 8677 1309 8711 1343
rect 8861 1309 8895 1343
rect 9413 1309 9447 1343
rect 10977 1309 11011 1343
rect 12541 1309 12575 1343
rect 15393 1309 15427 1343
rect 17693 1309 17727 1343
rect 14013 1173 14047 1207
rect 15577 1173 15611 1207
rect 18337 1173 18371 1207
rect 19625 1173 19659 1207
rect 8493 901 8527 935
rect 9965 901 9999 935
rect 11345 901 11379 935
rect 13093 901 13127 935
rect 14841 901 14875 935
rect 7757 833 7791 867
rect 7665 765 7699 799
rect 8033 765 8067 799
rect 8217 765 8251 799
rect 8672 765 8706 799
rect 8769 765 8803 799
rect 9045 765 9079 799
rect 10144 765 10178 799
rect 10241 765 10275 799
rect 10517 765 10551 799
rect 11524 765 11558 799
rect 11621 765 11655 799
rect 11897 765 11931 799
rect 12541 765 12575 799
rect 12725 765 12759 799
rect 12817 765 12851 799
rect 12961 765 12995 799
rect 14289 765 14323 799
rect 14565 765 14599 799
rect 14709 765 14743 799
rect 7021 697 7055 731
rect 8861 697 8895 731
rect 10333 697 10367 731
rect 11713 697 11747 731
rect 14473 697 14507 731
<< metal1 >>
rect 17494 17484 17500 17536
rect 17552 17524 17558 17536
rect 17770 17524 17776 17536
rect 17552 17496 17776 17524
rect 17552 17484 17558 17496
rect 17770 17484 17776 17496
rect 17828 17484 17834 17536
rect 552 17434 27416 17456
rect 552 17382 3756 17434
rect 3808 17382 3820 17434
rect 3872 17382 3884 17434
rect 3936 17382 3948 17434
rect 4000 17382 4012 17434
rect 4064 17382 10472 17434
rect 10524 17382 10536 17434
rect 10588 17382 10600 17434
rect 10652 17382 10664 17434
rect 10716 17382 10728 17434
rect 10780 17382 17188 17434
rect 17240 17382 17252 17434
rect 17304 17382 17316 17434
rect 17368 17382 17380 17434
rect 17432 17382 17444 17434
rect 17496 17382 23904 17434
rect 23956 17382 23968 17434
rect 24020 17382 24032 17434
rect 24084 17382 24096 17434
rect 24148 17382 24160 17434
rect 24212 17382 27416 17434
rect 552 17360 27416 17382
rect 842 17280 848 17332
rect 900 17280 906 17332
rect 1486 17280 1492 17332
rect 1544 17280 1550 17332
rect 3602 17280 3608 17332
rect 3660 17320 3666 17332
rect 4065 17323 4123 17329
rect 4065 17320 4077 17323
rect 3660 17292 4077 17320
rect 3660 17280 3666 17292
rect 4065 17289 4077 17292
rect 4111 17289 4123 17323
rect 4065 17283 4123 17289
rect 5629 17323 5687 17329
rect 5629 17289 5641 17323
rect 5675 17320 5687 17323
rect 5902 17320 5908 17332
rect 5675 17292 5908 17320
rect 5675 17289 5687 17292
rect 5629 17283 5687 17289
rect 5902 17280 5908 17292
rect 5960 17280 5966 17332
rect 6546 17280 6552 17332
rect 6604 17320 6610 17332
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 6604 17292 6837 17320
rect 6604 17280 6610 17292
rect 6825 17289 6837 17292
rect 6871 17289 6883 17323
rect 6825 17283 6883 17289
rect 9122 17280 9128 17332
rect 9180 17320 9186 17332
rect 9217 17323 9275 17329
rect 9217 17320 9229 17323
rect 9180 17292 9229 17320
rect 9180 17280 9186 17292
rect 9217 17289 9229 17292
rect 9263 17289 9275 17323
rect 9217 17283 9275 17289
rect 12437 17323 12495 17329
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12986 17320 12992 17332
rect 12483 17292 12992 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12986 17280 12992 17292
rect 13044 17280 13050 17332
rect 13173 17323 13231 17329
rect 13173 17289 13185 17323
rect 13219 17320 13231 17323
rect 14274 17320 14280 17332
rect 13219 17292 14280 17320
rect 13219 17289 13231 17292
rect 13173 17283 13231 17289
rect 14274 17280 14280 17292
rect 14332 17280 14338 17332
rect 15562 17280 15568 17332
rect 15620 17320 15626 17332
rect 16301 17323 16359 17329
rect 16301 17320 16313 17323
rect 15620 17292 16313 17320
rect 15620 17280 15626 17292
rect 16301 17289 16313 17292
rect 16347 17289 16359 17323
rect 23385 17323 23443 17329
rect 23385 17320 23397 17323
rect 16301 17283 16359 17289
rect 19996 17292 23397 17320
rect 6641 17255 6699 17261
rect 6641 17221 6653 17255
rect 6687 17252 6699 17255
rect 7190 17252 7196 17264
rect 6687 17224 7196 17252
rect 6687 17221 6699 17224
rect 6641 17215 6699 17221
rect 7190 17212 7196 17224
rect 7248 17212 7254 17264
rect 12805 17255 12863 17261
rect 12805 17221 12817 17255
rect 12851 17252 12863 17255
rect 13630 17252 13636 17264
rect 12851 17224 13636 17252
rect 12851 17221 12863 17224
rect 12805 17215 12863 17221
rect 13630 17212 13636 17224
rect 13688 17212 13694 17264
rect 14918 17212 14924 17264
rect 14976 17252 14982 17264
rect 15657 17255 15715 17261
rect 15657 17252 15669 17255
rect 14976 17224 15669 17252
rect 14976 17212 14982 17224
rect 15657 17221 15669 17224
rect 15703 17221 15715 17255
rect 15657 17215 15715 17221
rect 16574 17212 16580 17264
rect 16632 17252 16638 17264
rect 19996 17261 20024 17292
rect 23385 17289 23397 17292
rect 23431 17289 23443 17323
rect 23385 17283 23443 17289
rect 17589 17255 17647 17261
rect 17589 17252 17601 17255
rect 16632 17224 17601 17252
rect 16632 17212 16638 17224
rect 17589 17221 17601 17224
rect 17635 17221 17647 17255
rect 17589 17215 17647 17221
rect 19981 17255 20039 17261
rect 19981 17221 19993 17255
rect 20027 17221 20039 17255
rect 19981 17215 20039 17221
rect 2682 17144 2688 17196
rect 2740 17184 2746 17196
rect 2777 17187 2835 17193
rect 2777 17184 2789 17187
rect 2740 17156 2789 17184
rect 2740 17144 2746 17156
rect 2777 17153 2789 17156
rect 2823 17153 2835 17187
rect 2777 17147 2835 17153
rect 3418 17144 3424 17196
rect 3476 17144 3482 17196
rect 4706 17144 4712 17196
rect 4764 17144 4770 17196
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 5353 17187 5411 17193
rect 5353 17184 5365 17187
rect 5316 17156 5365 17184
rect 5316 17144 5322 17156
rect 5353 17153 5365 17156
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 6273 17187 6331 17193
rect 6273 17153 6285 17187
rect 6319 17184 6331 17187
rect 8478 17184 8484 17196
rect 6319 17156 8484 17184
rect 6319 17153 6331 17156
rect 6273 17147 6331 17153
rect 8478 17144 8484 17156
rect 8536 17144 8542 17196
rect 9858 17144 9864 17196
rect 9916 17184 9922 17196
rect 9916 17156 10456 17184
rect 9916 17144 9922 17156
rect 5902 17076 5908 17128
rect 5960 17116 5966 17128
rect 6457 17119 6515 17125
rect 6457 17116 6469 17119
rect 5960 17088 6469 17116
rect 5960 17076 5966 17088
rect 6457 17085 6469 17088
rect 6503 17085 6515 17119
rect 6457 17079 6515 17085
rect 10045 17119 10103 17125
rect 10045 17085 10057 17119
rect 10091 17085 10103 17119
rect 10045 17079 10103 17085
rect 5994 17008 6000 17060
rect 6052 17008 6058 17060
rect 10060 17048 10088 17079
rect 10134 17076 10140 17128
rect 10192 17076 10198 17128
rect 10226 17076 10232 17128
rect 10284 17076 10290 17128
rect 10428 17125 10456 17156
rect 25222 17144 25228 17196
rect 25280 17184 25286 17196
rect 25280 17156 26188 17184
rect 25280 17144 25286 17156
rect 10413 17119 10471 17125
rect 10413 17085 10425 17119
rect 10459 17085 10471 17119
rect 10413 17079 10471 17085
rect 10686 17076 10692 17128
rect 10744 17116 10750 17128
rect 11517 17119 11575 17125
rect 11517 17116 11529 17119
rect 10744 17088 11529 17116
rect 10744 17076 10750 17088
rect 11517 17085 11529 17088
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 12621 17119 12679 17125
rect 12621 17085 12633 17119
rect 12667 17116 12679 17119
rect 12894 17116 12900 17128
rect 12667 17088 12900 17116
rect 12667 17085 12679 17088
rect 12621 17079 12679 17085
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 12989 17119 13047 17125
rect 12989 17085 13001 17119
rect 13035 17116 13047 17119
rect 13078 17116 13084 17128
rect 13035 17088 13084 17116
rect 13035 17085 13047 17088
rect 12989 17079 13047 17085
rect 13078 17076 13084 17088
rect 13136 17076 13142 17128
rect 13357 17119 13415 17125
rect 13357 17085 13369 17119
rect 13403 17116 13415 17119
rect 13538 17116 13544 17128
rect 13403 17088 13544 17116
rect 13403 17085 13415 17088
rect 13357 17079 13415 17085
rect 13538 17076 13544 17088
rect 13596 17076 13602 17128
rect 14366 17076 14372 17128
rect 14424 17076 14430 17128
rect 14550 17076 14556 17128
rect 14608 17116 14614 17128
rect 15289 17119 15347 17125
rect 15289 17116 15301 17119
rect 14608 17088 15301 17116
rect 14608 17076 14614 17088
rect 15289 17085 15301 17088
rect 15335 17085 15347 17119
rect 15289 17079 15347 17085
rect 15473 17119 15531 17125
rect 15473 17085 15485 17119
rect 15519 17116 15531 17119
rect 15838 17116 15844 17128
rect 15519 17088 15844 17116
rect 15519 17085 15531 17088
rect 15473 17079 15531 17085
rect 15838 17076 15844 17088
rect 15896 17076 15902 17128
rect 16117 17119 16175 17125
rect 16117 17085 16129 17119
rect 16163 17085 16175 17119
rect 16117 17079 16175 17085
rect 10965 17051 11023 17057
rect 10965 17048 10977 17051
rect 10060 17020 10977 17048
rect 10965 17017 10977 17020
rect 11011 17017 11023 17051
rect 10965 17011 11023 17017
rect 15562 17008 15568 17060
rect 15620 17048 15626 17060
rect 16132 17048 16160 17079
rect 16206 17076 16212 17128
rect 16264 17116 16270 17128
rect 16485 17119 16543 17125
rect 16485 17116 16497 17119
rect 16264 17088 16497 17116
rect 16264 17076 16270 17088
rect 16485 17085 16497 17088
rect 16531 17085 16543 17119
rect 16485 17079 16543 17085
rect 16850 17076 16856 17128
rect 16908 17116 16914 17128
rect 16945 17119 17003 17125
rect 16945 17116 16957 17119
rect 16908 17088 16957 17116
rect 16908 17076 16914 17088
rect 16945 17085 16957 17088
rect 16991 17085 17003 17119
rect 16945 17079 17003 17085
rect 17770 17076 17776 17128
rect 17828 17076 17834 17128
rect 19426 17076 19432 17128
rect 19484 17116 19490 17128
rect 20441 17119 20499 17125
rect 20441 17116 20453 17119
rect 19484 17088 20453 17116
rect 19484 17076 19490 17088
rect 20441 17085 20453 17088
rect 20487 17085 20499 17119
rect 20441 17079 20499 17085
rect 21634 17076 21640 17128
rect 21692 17076 21698 17128
rect 22002 17076 22008 17128
rect 22060 17116 22066 17128
rect 22281 17119 22339 17125
rect 22281 17116 22293 17119
rect 22060 17088 22293 17116
rect 22060 17076 22066 17088
rect 22281 17085 22293 17088
rect 22327 17085 22339 17119
rect 22281 17079 22339 17085
rect 22646 17076 22652 17128
rect 22704 17116 22710 17128
rect 22925 17119 22983 17125
rect 22925 17116 22937 17119
rect 22704 17088 22937 17116
rect 22704 17076 22710 17088
rect 22925 17085 22937 17088
rect 22971 17085 22983 17119
rect 22925 17079 22983 17085
rect 23290 17076 23296 17128
rect 23348 17116 23354 17128
rect 23569 17119 23627 17125
rect 23569 17116 23581 17119
rect 23348 17088 23581 17116
rect 23348 17076 23354 17088
rect 23569 17085 23581 17088
rect 23615 17085 23627 17119
rect 23569 17079 23627 17085
rect 23750 17076 23756 17128
rect 23808 17116 23814 17128
rect 24213 17119 24271 17125
rect 24213 17116 24225 17119
rect 23808 17088 24225 17116
rect 23808 17076 23814 17088
rect 24213 17085 24225 17088
rect 24259 17085 24271 17119
rect 24213 17079 24271 17085
rect 24578 17076 24584 17128
rect 24636 17116 24642 17128
rect 24857 17119 24915 17125
rect 24857 17116 24869 17119
rect 24636 17088 24869 17116
rect 24636 17076 24642 17088
rect 24857 17085 24869 17088
rect 24903 17085 24915 17119
rect 24857 17079 24915 17085
rect 25774 17076 25780 17128
rect 25832 17076 25838 17128
rect 26160 17125 26188 17156
rect 26145 17119 26203 17125
rect 26145 17085 26157 17119
rect 26191 17085 26203 17119
rect 26145 17079 26203 17085
rect 26510 17076 26516 17128
rect 26568 17116 26574 17128
rect 26605 17119 26663 17125
rect 26605 17116 26617 17119
rect 26568 17088 26617 17116
rect 26568 17076 26574 17088
rect 26605 17085 26617 17088
rect 26651 17085 26663 17119
rect 26605 17079 26663 17085
rect 15620 17020 16160 17048
rect 15620 17008 15626 17020
rect 19518 17008 19524 17060
rect 19576 17048 19582 17060
rect 19613 17051 19671 17057
rect 19613 17048 19625 17051
rect 19576 17020 19625 17048
rect 19576 17008 19582 17020
rect 19613 17017 19625 17020
rect 19659 17017 19671 17051
rect 19613 17011 19671 17017
rect 9766 16940 9772 16992
rect 9824 16940 9830 16992
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 13725 16983 13783 16989
rect 13725 16980 13737 16983
rect 12584 16952 13737 16980
rect 12584 16940 12590 16952
rect 13725 16949 13737 16952
rect 13771 16949 13783 16983
rect 13725 16943 13783 16949
rect 14734 16940 14740 16992
rect 14792 16940 14798 16992
rect 16666 16940 16672 16992
rect 16724 16940 16730 16992
rect 17034 16940 17040 16992
rect 17092 16980 17098 16992
rect 17129 16983 17187 16989
rect 17129 16980 17141 16983
rect 17092 16952 17141 16980
rect 17092 16940 17098 16952
rect 17129 16949 17141 16952
rect 17175 16949 17187 16983
rect 17129 16943 17187 16949
rect 19794 16940 19800 16992
rect 19852 16980 19858 16992
rect 20073 16983 20131 16989
rect 20073 16980 20085 16983
rect 19852 16952 20085 16980
rect 19852 16940 19858 16952
rect 20073 16949 20085 16952
rect 20119 16949 20131 16983
rect 20073 16943 20131 16949
rect 20257 16983 20315 16989
rect 20257 16949 20269 16983
rect 20303 16980 20315 16983
rect 20346 16980 20352 16992
rect 20303 16952 20352 16980
rect 20303 16949 20315 16952
rect 20257 16943 20315 16949
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 21450 16940 21456 16992
rect 21508 16940 21514 16992
rect 21726 16940 21732 16992
rect 21784 16980 21790 16992
rect 22097 16983 22155 16989
rect 22097 16980 22109 16983
rect 21784 16952 22109 16980
rect 21784 16940 21790 16952
rect 22097 16949 22109 16952
rect 22143 16949 22155 16983
rect 22097 16943 22155 16949
rect 22738 16940 22744 16992
rect 22796 16940 22802 16992
rect 24026 16940 24032 16992
rect 24084 16940 24090 16992
rect 24670 16940 24676 16992
rect 24728 16940 24734 16992
rect 24854 16940 24860 16992
rect 24912 16980 24918 16992
rect 25225 16983 25283 16989
rect 25225 16980 25237 16983
rect 24912 16952 25237 16980
rect 24912 16940 24918 16952
rect 25225 16949 25237 16952
rect 25271 16949 25283 16983
rect 25225 16943 25283 16949
rect 25958 16940 25964 16992
rect 26016 16940 26022 16992
rect 26786 16940 26792 16992
rect 26844 16940 26850 16992
rect 552 16890 27576 16912
rect 552 16838 7114 16890
rect 7166 16838 7178 16890
rect 7230 16838 7242 16890
rect 7294 16838 7306 16890
rect 7358 16838 7370 16890
rect 7422 16838 13830 16890
rect 13882 16838 13894 16890
rect 13946 16838 13958 16890
rect 14010 16838 14022 16890
rect 14074 16838 14086 16890
rect 14138 16838 20546 16890
rect 20598 16838 20610 16890
rect 20662 16838 20674 16890
rect 20726 16838 20738 16890
rect 20790 16838 20802 16890
rect 20854 16838 27262 16890
rect 27314 16838 27326 16890
rect 27378 16838 27390 16890
rect 27442 16838 27454 16890
rect 27506 16838 27518 16890
rect 27570 16838 27576 16890
rect 552 16816 27576 16838
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 10965 16779 11023 16785
rect 10965 16776 10977 16779
rect 10192 16748 10977 16776
rect 10192 16736 10198 16748
rect 10965 16745 10977 16748
rect 11011 16745 11023 16779
rect 10965 16739 11023 16745
rect 11698 16736 11704 16788
rect 11756 16776 11762 16788
rect 12161 16779 12219 16785
rect 12161 16776 12173 16779
rect 11756 16748 12173 16776
rect 11756 16736 11762 16748
rect 12161 16745 12173 16748
rect 12207 16745 12219 16779
rect 12161 16739 12219 16745
rect 12342 16736 12348 16788
rect 12400 16776 12406 16788
rect 12621 16779 12679 16785
rect 12621 16776 12633 16779
rect 12400 16748 12633 16776
rect 12400 16736 12406 16748
rect 12621 16745 12633 16748
rect 12667 16745 12679 16779
rect 12621 16739 12679 16745
rect 14185 16779 14243 16785
rect 14185 16745 14197 16779
rect 14231 16776 14243 16779
rect 14366 16776 14372 16788
rect 14231 16748 14372 16776
rect 14231 16745 14243 16748
rect 14185 16739 14243 16745
rect 14366 16736 14372 16748
rect 14424 16776 14430 16788
rect 15378 16776 15384 16788
rect 14424 16748 15384 16776
rect 14424 16736 14430 16748
rect 15378 16736 15384 16748
rect 15436 16736 15442 16788
rect 17126 16736 17132 16788
rect 17184 16736 17190 16788
rect 17957 16779 18015 16785
rect 17957 16745 17969 16779
rect 18003 16776 18015 16779
rect 18506 16776 18512 16788
rect 18003 16748 18512 16776
rect 18003 16745 18015 16748
rect 17957 16739 18015 16745
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 19061 16779 19119 16785
rect 19061 16745 19073 16779
rect 19107 16776 19119 16779
rect 19150 16776 19156 16788
rect 19107 16748 19156 16776
rect 19107 16745 19119 16748
rect 19061 16739 19119 16745
rect 19150 16736 19156 16748
rect 19208 16736 19214 16788
rect 19978 16736 19984 16788
rect 20036 16776 20042 16788
rect 20073 16779 20131 16785
rect 20073 16776 20085 16779
rect 20036 16748 20085 16776
rect 20036 16736 20042 16748
rect 20073 16745 20085 16748
rect 20119 16745 20131 16779
rect 20349 16779 20407 16785
rect 20349 16776 20361 16779
rect 20073 16739 20131 16745
rect 20180 16748 20361 16776
rect 9576 16711 9634 16717
rect 6104 16680 7788 16708
rect 4525 16643 4583 16649
rect 4525 16609 4537 16643
rect 4571 16640 4583 16643
rect 4614 16640 4620 16652
rect 4571 16612 4620 16640
rect 4571 16609 4583 16612
rect 4525 16603 4583 16609
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 4893 16643 4951 16649
rect 4893 16609 4905 16643
rect 4939 16640 4951 16643
rect 5258 16640 5264 16652
rect 4939 16612 5264 16640
rect 4939 16609 4951 16612
rect 4893 16603 4951 16609
rect 5258 16600 5264 16612
rect 5316 16600 5322 16652
rect 6104 16649 6132 16680
rect 7760 16652 7788 16680
rect 9576 16677 9588 16711
rect 9622 16708 9634 16711
rect 9766 16708 9772 16720
rect 9622 16680 9772 16708
rect 9622 16677 9634 16680
rect 9576 16671 9634 16677
rect 9766 16668 9772 16680
rect 9824 16668 9830 16720
rect 11146 16668 11152 16720
rect 11204 16708 11210 16720
rect 11241 16711 11299 16717
rect 11241 16708 11253 16711
rect 11204 16680 11253 16708
rect 11204 16668 11210 16680
rect 11241 16677 11253 16680
rect 11287 16708 11299 16711
rect 14550 16708 14556 16720
rect 11287 16680 14556 16708
rect 11287 16677 11299 16680
rect 11241 16671 11299 16677
rect 14550 16668 14556 16680
rect 14608 16668 14614 16720
rect 15286 16668 15292 16720
rect 15344 16708 15350 16720
rect 15344 16680 15976 16708
rect 15344 16668 15350 16680
rect 6362 16649 6368 16652
rect 6089 16643 6147 16649
rect 6089 16609 6101 16643
rect 6135 16609 6147 16643
rect 6089 16603 6147 16609
rect 6356 16603 6368 16649
rect 6362 16600 6368 16603
rect 6420 16600 6426 16652
rect 7742 16600 7748 16652
rect 7800 16600 7806 16652
rect 8012 16643 8070 16649
rect 8012 16609 8024 16643
rect 8058 16640 8070 16643
rect 8478 16640 8484 16652
rect 8058 16612 8484 16640
rect 8058 16609 8070 16612
rect 8012 16603 8070 16609
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 8570 16600 8576 16652
rect 8628 16640 8634 16652
rect 9309 16643 9367 16649
rect 9309 16640 9321 16643
rect 8628 16612 9321 16640
rect 8628 16600 8634 16612
rect 9309 16609 9321 16612
rect 9355 16609 9367 16643
rect 9309 16603 9367 16609
rect 10870 16600 10876 16652
rect 10928 16640 10934 16652
rect 10965 16643 11023 16649
rect 10965 16640 10977 16643
rect 10928 16612 10977 16640
rect 10928 16600 10934 16612
rect 10965 16609 10977 16612
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 11112 16612 11836 16640
rect 11112 16600 11118 16612
rect 2038 16464 2044 16516
rect 2096 16504 2102 16516
rect 5902 16504 5908 16516
rect 2096 16476 5908 16504
rect 2096 16464 2102 16476
rect 5902 16464 5908 16476
rect 5960 16464 5966 16516
rect 10686 16464 10692 16516
rect 10744 16504 10750 16516
rect 10962 16504 10968 16516
rect 10744 16476 10968 16504
rect 10744 16464 10750 16476
rect 10962 16464 10968 16476
rect 11020 16464 11026 16516
rect 11057 16507 11115 16513
rect 11057 16473 11069 16507
rect 11103 16504 11115 16507
rect 11238 16504 11244 16516
rect 11103 16476 11244 16504
rect 11103 16473 11115 16476
rect 11057 16467 11115 16473
rect 11238 16464 11244 16476
rect 11296 16464 11302 16516
rect 11808 16513 11836 16612
rect 11882 16600 11888 16652
rect 11940 16640 11946 16652
rect 11977 16643 12035 16649
rect 11977 16640 11989 16643
rect 11940 16612 11989 16640
rect 11940 16600 11946 16612
rect 11977 16609 11989 16612
rect 12023 16609 12035 16643
rect 11977 16603 12035 16609
rect 12342 16600 12348 16652
rect 12400 16600 12406 16652
rect 12434 16600 12440 16652
rect 12492 16600 12498 16652
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 13061 16643 13119 16649
rect 13061 16640 13073 16643
rect 12676 16612 13073 16640
rect 12676 16600 12682 16612
rect 13061 16609 13073 16612
rect 13107 16609 13119 16643
rect 13061 16603 13119 16609
rect 14461 16643 14519 16649
rect 14461 16609 14473 16643
rect 14507 16640 14519 16643
rect 14568 16640 14596 16668
rect 14507 16612 14596 16640
rect 14507 16609 14519 16612
rect 14461 16603 14519 16609
rect 12802 16532 12808 16584
rect 12860 16532 12866 16584
rect 14568 16513 14596 16612
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15948 16649 15976 16680
rect 16022 16668 16028 16720
rect 16080 16708 16086 16720
rect 16209 16711 16267 16717
rect 16209 16708 16221 16711
rect 16080 16680 16221 16708
rect 16080 16668 16086 16680
rect 16209 16677 16221 16680
rect 16255 16708 16267 16711
rect 16666 16708 16672 16720
rect 16255 16680 16672 16708
rect 16255 16677 16267 16680
rect 16209 16671 16267 16677
rect 16666 16668 16672 16680
rect 16724 16668 16730 16720
rect 19610 16668 19616 16720
rect 19668 16708 19674 16720
rect 20180 16708 20208 16748
rect 20349 16745 20361 16748
rect 20395 16745 20407 16779
rect 20349 16739 20407 16745
rect 21542 16736 21548 16788
rect 21600 16776 21606 16788
rect 21729 16779 21787 16785
rect 21729 16776 21741 16779
rect 21600 16748 21741 16776
rect 21600 16736 21606 16748
rect 21729 16745 21741 16748
rect 21775 16745 21787 16779
rect 21729 16739 21787 16745
rect 25774 16736 25780 16788
rect 25832 16776 25838 16788
rect 25832 16748 26556 16776
rect 25832 16736 25838 16748
rect 20809 16711 20867 16717
rect 20809 16708 20821 16711
rect 19668 16680 20208 16708
rect 20272 16680 20821 16708
rect 19668 16668 19674 16680
rect 15666 16643 15724 16649
rect 15666 16640 15678 16643
rect 15252 16612 15678 16640
rect 15252 16600 15258 16612
rect 15666 16609 15678 16612
rect 15712 16609 15724 16643
rect 15666 16603 15724 16609
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16609 15991 16643
rect 15933 16603 15991 16609
rect 16393 16643 16451 16649
rect 16393 16609 16405 16643
rect 16439 16640 16451 16643
rect 16850 16640 16856 16652
rect 16439 16612 16856 16640
rect 16439 16609 16451 16612
rect 16393 16603 16451 16609
rect 16850 16600 16856 16612
rect 16908 16640 16914 16652
rect 17589 16643 17647 16649
rect 17589 16640 17601 16643
rect 16908 16612 17601 16640
rect 16908 16600 16914 16612
rect 17589 16609 17601 16612
rect 17635 16640 17647 16643
rect 18417 16643 18475 16649
rect 18417 16640 18429 16643
rect 17635 16612 18429 16640
rect 17635 16609 17647 16612
rect 17589 16603 17647 16609
rect 18417 16609 18429 16612
rect 18463 16640 18475 16643
rect 19518 16640 19524 16652
rect 18463 16612 19524 16640
rect 18463 16609 18475 16612
rect 18417 16603 18475 16609
rect 19518 16600 19524 16612
rect 19576 16640 19582 16652
rect 20272 16640 20300 16680
rect 20809 16677 20821 16680
rect 20855 16708 20867 16711
rect 21269 16711 21327 16717
rect 21269 16708 21281 16711
rect 20855 16680 21281 16708
rect 20855 16677 20867 16680
rect 20809 16671 20867 16677
rect 21269 16677 21281 16680
rect 21315 16677 21327 16711
rect 25133 16711 25191 16717
rect 21269 16671 21327 16677
rect 24688 16680 25084 16708
rect 24688 16649 24716 16680
rect 19576 16612 20300 16640
rect 24489 16643 24547 16649
rect 19576 16600 19582 16612
rect 19628 16581 19656 16612
rect 24489 16609 24501 16643
rect 24535 16640 24547 16643
rect 24673 16643 24731 16649
rect 24535 16612 24624 16640
rect 24535 16609 24547 16612
rect 24489 16603 24547 16609
rect 19613 16575 19671 16581
rect 19613 16541 19625 16575
rect 19659 16541 19671 16575
rect 21726 16572 21732 16584
rect 19613 16535 19671 16541
rect 19996 16544 21732 16572
rect 11793 16507 11851 16513
rect 11793 16473 11805 16507
rect 11839 16473 11851 16507
rect 11793 16467 11851 16473
rect 14553 16507 14611 16513
rect 14553 16473 14565 16507
rect 14599 16473 14611 16507
rect 14553 16467 14611 16473
rect 17313 16507 17371 16513
rect 17313 16473 17325 16507
rect 17359 16504 17371 16507
rect 17678 16504 17684 16516
rect 17359 16476 17684 16504
rect 17359 16473 17371 16476
rect 17313 16467 17371 16473
rect 17678 16464 17684 16476
rect 17736 16464 17742 16516
rect 18138 16464 18144 16516
rect 18196 16464 18202 16516
rect 19996 16513 20024 16544
rect 21726 16532 21732 16544
rect 21784 16532 21790 16584
rect 24596 16572 24624 16612
rect 24673 16609 24685 16643
rect 24719 16609 24731 16643
rect 24673 16603 24731 16609
rect 24762 16600 24768 16652
rect 24820 16600 24826 16652
rect 24854 16600 24860 16652
rect 24912 16600 24918 16652
rect 25056 16640 25084 16680
rect 25133 16677 25145 16711
rect 25179 16708 25191 16711
rect 25179 16680 25820 16708
rect 25179 16677 25191 16680
rect 25133 16671 25191 16677
rect 25792 16649 25820 16680
rect 25777 16643 25835 16649
rect 25056 16612 25728 16640
rect 25314 16572 25320 16584
rect 24596 16544 25320 16572
rect 25314 16532 25320 16544
rect 25372 16532 25378 16584
rect 25700 16572 25728 16612
rect 25777 16609 25789 16643
rect 25823 16609 25835 16643
rect 25777 16603 25835 16609
rect 25866 16600 25872 16652
rect 25924 16640 25930 16652
rect 26145 16643 26203 16649
rect 26145 16640 26157 16643
rect 25924 16612 26157 16640
rect 25924 16600 25930 16612
rect 26145 16609 26157 16612
rect 26191 16609 26203 16643
rect 26145 16603 26203 16609
rect 26418 16600 26424 16652
rect 26476 16600 26482 16652
rect 26528 16649 26556 16748
rect 26789 16711 26847 16717
rect 26789 16677 26801 16711
rect 26835 16708 26847 16711
rect 27062 16708 27068 16720
rect 26835 16680 27068 16708
rect 26835 16677 26847 16680
rect 26789 16671 26847 16677
rect 27062 16668 27068 16680
rect 27120 16668 27126 16720
rect 26514 16643 26572 16649
rect 26514 16609 26526 16643
rect 26560 16609 26572 16643
rect 26514 16603 26572 16609
rect 26694 16600 26700 16652
rect 26752 16600 26758 16652
rect 26878 16600 26884 16652
rect 26936 16649 26942 16652
rect 26936 16603 26944 16649
rect 26936 16600 26942 16603
rect 26234 16572 26240 16584
rect 25700 16544 26240 16572
rect 26234 16532 26240 16544
rect 26292 16532 26298 16584
rect 19245 16507 19303 16513
rect 19245 16473 19257 16507
rect 19291 16473 19303 16507
rect 19245 16467 19303 16473
rect 19981 16507 20039 16513
rect 19981 16473 19993 16507
rect 20027 16473 20039 16507
rect 19981 16467 20039 16473
rect 20533 16507 20591 16513
rect 20533 16473 20545 16507
rect 20579 16504 20591 16507
rect 21450 16504 21456 16516
rect 20579 16476 21456 16504
rect 20579 16473 20591 16476
rect 20533 16467 20591 16473
rect 7469 16439 7527 16445
rect 7469 16405 7481 16439
rect 7515 16436 7527 16439
rect 8018 16436 8024 16448
rect 7515 16408 8024 16436
rect 7515 16405 7527 16408
rect 7469 16399 7527 16405
rect 8018 16396 8024 16408
rect 8076 16396 8082 16448
rect 9125 16439 9183 16445
rect 9125 16405 9137 16439
rect 9171 16436 9183 16439
rect 9490 16436 9496 16448
rect 9171 16408 9496 16436
rect 9171 16405 9183 16408
rect 9125 16399 9183 16405
rect 9490 16396 9496 16408
rect 9548 16396 9554 16448
rect 13722 16396 13728 16448
rect 13780 16436 13786 16448
rect 14369 16439 14427 16445
rect 14369 16436 14381 16439
rect 13780 16408 14381 16436
rect 13780 16396 13786 16408
rect 14369 16405 14381 16408
rect 14415 16405 14427 16439
rect 19260 16436 19288 16467
rect 21450 16464 21456 16476
rect 21508 16464 21514 16516
rect 21637 16507 21695 16513
rect 21637 16473 21649 16507
rect 21683 16504 21695 16507
rect 22738 16504 22744 16516
rect 21683 16476 22744 16504
rect 21683 16473 21695 16476
rect 21637 16467 21695 16473
rect 22738 16464 22744 16476
rect 22796 16464 22802 16516
rect 24026 16436 24032 16448
rect 19260 16408 24032 16436
rect 14369 16399 14427 16405
rect 24026 16396 24032 16408
rect 24084 16396 24090 16448
rect 25222 16396 25228 16448
rect 25280 16396 25286 16448
rect 25406 16396 25412 16448
rect 25464 16436 25470 16448
rect 25961 16439 26019 16445
rect 25961 16436 25973 16439
rect 25464 16408 25973 16436
rect 25464 16396 25470 16408
rect 25961 16405 25973 16408
rect 26007 16405 26019 16439
rect 25961 16399 26019 16405
rect 26970 16396 26976 16448
rect 27028 16436 27034 16448
rect 27065 16439 27123 16445
rect 27065 16436 27077 16439
rect 27028 16408 27077 16436
rect 27028 16396 27034 16408
rect 27065 16405 27077 16408
rect 27111 16405 27123 16439
rect 27065 16399 27123 16405
rect 552 16346 27416 16368
rect 552 16294 3756 16346
rect 3808 16294 3820 16346
rect 3872 16294 3884 16346
rect 3936 16294 3948 16346
rect 4000 16294 4012 16346
rect 4064 16294 10472 16346
rect 10524 16294 10536 16346
rect 10588 16294 10600 16346
rect 10652 16294 10664 16346
rect 10716 16294 10728 16346
rect 10780 16294 17188 16346
rect 17240 16294 17252 16346
rect 17304 16294 17316 16346
rect 17368 16294 17380 16346
rect 17432 16294 17444 16346
rect 17496 16294 23904 16346
rect 23956 16294 23968 16346
rect 24020 16294 24032 16346
rect 24084 16294 24096 16346
rect 24148 16294 24160 16346
rect 24212 16294 27416 16346
rect 552 16272 27416 16294
rect 5902 16192 5908 16244
rect 5960 16232 5966 16244
rect 5997 16235 6055 16241
rect 5997 16232 6009 16235
rect 5960 16204 6009 16232
rect 5960 16192 5966 16204
rect 5997 16201 6009 16204
rect 6043 16201 6055 16235
rect 5997 16195 6055 16201
rect 6362 16192 6368 16244
rect 6420 16192 6426 16244
rect 8478 16192 8484 16244
rect 8536 16232 8542 16244
rect 8941 16235 8999 16241
rect 8941 16232 8953 16235
rect 8536 16204 8953 16232
rect 8536 16192 8542 16204
rect 8941 16201 8953 16204
rect 8987 16201 8999 16235
rect 8941 16195 8999 16201
rect 9769 16235 9827 16241
rect 9769 16201 9781 16235
rect 9815 16201 9827 16235
rect 9769 16195 9827 16201
rect 10045 16235 10103 16241
rect 10045 16201 10057 16235
rect 10091 16232 10103 16235
rect 10226 16232 10232 16244
rect 10091 16204 10232 16232
rect 10091 16201 10103 16204
rect 10045 16195 10103 16201
rect 8757 16167 8815 16173
rect 7024 16136 8708 16164
rect 7024 16040 7052 16136
rect 8018 16056 8024 16108
rect 8076 16056 8082 16108
rect 8680 16096 8708 16136
rect 8757 16133 8769 16167
rect 8803 16164 8815 16167
rect 9674 16164 9680 16176
rect 8803 16136 9680 16164
rect 8803 16133 8815 16136
rect 8757 16127 8815 16133
rect 9674 16124 9680 16136
rect 9732 16124 9738 16176
rect 9784 16164 9812 16195
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 10870 16192 10876 16244
rect 10928 16232 10934 16244
rect 10928 16204 11100 16232
rect 10928 16192 10934 16204
rect 10962 16164 10968 16176
rect 9784 16136 10968 16164
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 11072 16164 11100 16204
rect 11146 16192 11152 16244
rect 11204 16192 11210 16244
rect 11793 16235 11851 16241
rect 11793 16201 11805 16235
rect 11839 16232 11851 16235
rect 12618 16232 12624 16244
rect 11839 16204 12624 16232
rect 11839 16201 11851 16204
rect 11793 16195 11851 16201
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 12713 16235 12771 16241
rect 12713 16201 12725 16235
rect 12759 16232 12771 16235
rect 12759 16204 12940 16232
rect 12759 16201 12771 16204
rect 12713 16195 12771 16201
rect 11701 16167 11759 16173
rect 11072 16136 11661 16164
rect 9766 16096 9772 16108
rect 8680 16068 9772 16096
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 9876 16068 10548 16096
rect 6638 15988 6644 16040
rect 6696 15988 6702 16040
rect 6733 16031 6791 16037
rect 6733 15997 6745 16031
rect 6779 15997 6791 16031
rect 6733 15991 6791 15997
rect 5902 15920 5908 15972
rect 5960 15920 5966 15972
rect 6748 15960 6776 15991
rect 6822 15988 6828 16040
rect 6880 15988 6886 16040
rect 7006 15988 7012 16040
rect 7064 15988 7070 16040
rect 8036 16028 8064 16056
rect 8481 16031 8539 16037
rect 8481 16028 8493 16031
rect 8036 16000 8493 16028
rect 8481 15997 8493 16000
rect 8527 15997 8539 16031
rect 8481 15991 8539 15997
rect 8846 15988 8852 16040
rect 8904 16028 8910 16040
rect 9125 16031 9183 16037
rect 9125 16028 9137 16031
rect 8904 16000 9137 16028
rect 8904 15988 8910 16000
rect 9125 15997 9137 16000
rect 9171 15997 9183 16031
rect 9125 15991 9183 15997
rect 9490 15988 9496 16040
rect 9548 15988 9554 16040
rect 9876 15960 9904 16068
rect 10134 15988 10140 16040
rect 10192 16037 10198 16040
rect 10192 16031 10228 16037
rect 10216 15997 10228 16031
rect 10192 15991 10228 15997
rect 10192 15988 10198 15991
rect 10520 15960 10548 16068
rect 10686 16056 10692 16108
rect 10744 16096 10750 16108
rect 10744 16068 11468 16096
rect 10744 16056 10750 16068
rect 10594 15988 10600 16040
rect 10652 16028 10658 16040
rect 10870 16028 10876 16040
rect 10652 16000 10876 16028
rect 10652 15988 10658 16000
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 10962 15988 10968 16040
rect 11020 15988 11026 16040
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 16028 11207 16031
rect 11238 16028 11244 16040
rect 11195 16000 11244 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 11054 15960 11060 15972
rect 6748 15932 9904 15960
rect 9968 15932 10272 15960
rect 10520 15932 11060 15960
rect 7466 15852 7472 15904
rect 7524 15852 7530 15904
rect 9968 15901 9996 15932
rect 10244 15901 10272 15932
rect 11054 15920 11060 15932
rect 11112 15920 11118 15972
rect 11164 15960 11192 15991
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 11440 16037 11468 16068
rect 11425 16031 11483 16037
rect 11425 15997 11437 16031
rect 11471 15997 11483 16031
rect 11633 16028 11661 16136
rect 11701 16133 11713 16167
rect 11747 16164 11759 16167
rect 12158 16164 12164 16176
rect 11747 16136 12164 16164
rect 11747 16133 11759 16136
rect 11701 16127 11759 16133
rect 12158 16124 12164 16136
rect 12216 16124 12222 16176
rect 12805 16099 12863 16105
rect 12805 16065 12817 16099
rect 12851 16065 12863 16099
rect 12805 16059 12863 16065
rect 11701 16031 11759 16037
rect 11701 16028 11713 16031
rect 11633 16000 11713 16028
rect 11425 15991 11483 15997
rect 11701 15997 11713 16000
rect 11747 15997 11759 16031
rect 11701 15991 11759 15997
rect 11716 15960 11744 15991
rect 11974 15988 11980 16040
rect 12032 15988 12038 16040
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 16028 12311 16031
rect 12345 16031 12403 16037
rect 12345 16028 12357 16031
rect 12299 16000 12357 16028
rect 12299 15997 12311 16000
rect 12253 15991 12311 15997
rect 12345 15997 12357 16000
rect 12391 15997 12403 16031
rect 12345 15991 12403 15997
rect 12526 15988 12532 16040
rect 12584 15988 12590 16040
rect 12710 15988 12716 16040
rect 12768 16028 12774 16040
rect 12820 16028 12848 16059
rect 12768 16000 12848 16028
rect 12768 15988 12774 16000
rect 12158 15960 12164 15972
rect 11164 15932 11560 15960
rect 11716 15932 12164 15960
rect 9953 15895 10011 15901
rect 9953 15861 9965 15895
rect 9999 15861 10011 15895
rect 9953 15855 10011 15861
rect 10229 15895 10287 15901
rect 10229 15861 10241 15895
rect 10275 15861 10287 15895
rect 10229 15855 10287 15861
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 11532 15901 11560 15932
rect 12158 15920 12164 15932
rect 12216 15960 12222 15972
rect 12912 15969 12940 16204
rect 13170 16192 13176 16244
rect 13228 16192 13234 16244
rect 15013 16235 15071 16241
rect 15013 16201 15025 16235
rect 15059 16232 15071 16235
rect 15194 16232 15200 16244
rect 15059 16204 15200 16232
rect 15059 16201 15071 16204
rect 15013 16195 15071 16201
rect 15194 16192 15200 16204
rect 15252 16192 15258 16244
rect 18138 16192 18144 16244
rect 18196 16232 18202 16244
rect 24670 16232 24676 16244
rect 18196 16204 24676 16232
rect 18196 16192 18202 16204
rect 24670 16192 24676 16204
rect 24728 16192 24734 16244
rect 13357 16167 13415 16173
rect 13357 16133 13369 16167
rect 13403 16133 13415 16167
rect 13357 16127 13415 16133
rect 12986 16056 12992 16108
rect 13044 16056 13050 16108
rect 13372 16096 13400 16127
rect 13446 16124 13452 16176
rect 13504 16164 13510 16176
rect 15473 16167 15531 16173
rect 15473 16164 15485 16167
rect 13504 16136 15485 16164
rect 13504 16124 13510 16136
rect 15473 16133 15485 16136
rect 15519 16133 15531 16167
rect 15473 16127 15531 16133
rect 17678 16124 17684 16176
rect 17736 16164 17742 16176
rect 25958 16164 25964 16176
rect 17736 16136 25964 16164
rect 17736 16124 17742 16136
rect 25958 16124 25964 16136
rect 26016 16124 26022 16176
rect 13372 16068 14596 16096
rect 13213 16031 13271 16037
rect 13213 15997 13225 16031
rect 13259 16028 13271 16031
rect 13722 16028 13728 16040
rect 13259 16000 13728 16028
rect 13259 15997 13271 16000
rect 13213 15991 13271 15997
rect 13722 15988 13728 16000
rect 13780 15988 13786 16040
rect 14182 15988 14188 16040
rect 14240 15988 14246 16040
rect 14366 15988 14372 16040
rect 14424 15988 14430 16040
rect 14568 16037 14596 16068
rect 23934 16056 23940 16108
rect 23992 16096 23998 16108
rect 26786 16096 26792 16108
rect 23992 16068 26792 16096
rect 23992 16056 23998 16068
rect 26786 16056 26792 16068
rect 26844 16056 26850 16108
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 15997 14611 16031
rect 14553 15991 14611 15997
rect 14642 15988 14648 16040
rect 14700 15988 14706 16040
rect 14734 15988 14740 16040
rect 14792 15988 14798 16040
rect 15289 16031 15347 16037
rect 15289 15997 15301 16031
rect 15335 16028 15347 16031
rect 15378 16028 15384 16040
rect 15335 16000 15384 16028
rect 15335 15997 15347 16000
rect 15289 15991 15347 15997
rect 15378 15988 15384 16000
rect 15436 15988 15442 16040
rect 18782 15988 18788 16040
rect 18840 15988 18846 16040
rect 20070 15988 20076 16040
rect 20128 15988 20134 16040
rect 20254 15988 20260 16040
rect 20312 15988 20318 16040
rect 21726 15988 21732 16040
rect 21784 15988 21790 16040
rect 24486 15988 24492 16040
rect 24544 16028 24550 16040
rect 24949 16031 25007 16037
rect 24949 16028 24961 16031
rect 24544 16000 24961 16028
rect 24544 15988 24550 16000
rect 24949 15997 24961 16000
rect 24995 15997 25007 16031
rect 24949 15991 25007 15997
rect 25314 15988 25320 16040
rect 25372 15988 25378 16040
rect 25498 15988 25504 16040
rect 25556 15988 25562 16040
rect 25593 16031 25651 16037
rect 25593 15997 25605 16031
rect 25639 15997 25651 16031
rect 25593 15991 25651 15997
rect 25685 16031 25743 16037
rect 25685 15997 25697 16031
rect 25731 16028 25743 16031
rect 26329 16031 26387 16037
rect 26329 16028 26341 16031
rect 25731 16000 26341 16028
rect 25731 15997 25743 16000
rect 25685 15991 25743 15997
rect 26329 15997 26341 16000
rect 26375 15997 26387 16031
rect 26329 15991 26387 15997
rect 12897 15963 12955 15969
rect 12897 15960 12909 15963
rect 12216 15932 12909 15960
rect 12216 15920 12222 15932
rect 12897 15929 12909 15932
rect 12943 15929 12955 15963
rect 12897 15923 12955 15929
rect 15105 15963 15163 15969
rect 15105 15929 15117 15963
rect 15151 15929 15163 15963
rect 25608 15960 25636 15991
rect 26602 15988 26608 16040
rect 26660 16028 26666 16040
rect 26881 16031 26939 16037
rect 26881 16028 26893 16031
rect 26660 16000 26893 16028
rect 26660 15988 26666 16000
rect 26881 15997 26893 16000
rect 26927 15997 26939 16031
rect 26881 15991 26939 15997
rect 15105 15923 15163 15929
rect 24964 15932 25636 15960
rect 10781 15895 10839 15901
rect 10781 15892 10793 15895
rect 10560 15864 10793 15892
rect 10560 15852 10566 15864
rect 10781 15861 10793 15864
rect 10827 15861 10839 15895
rect 10781 15855 10839 15861
rect 11517 15895 11575 15901
rect 11517 15861 11529 15895
rect 11563 15892 11575 15895
rect 13170 15892 13176 15904
rect 11563 15864 13176 15892
rect 11563 15861 11575 15864
rect 11517 15855 11575 15861
rect 13170 15852 13176 15864
rect 13228 15852 13234 15904
rect 13630 15852 13636 15904
rect 13688 15852 13694 15904
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 15120 15892 15148 15923
rect 24964 15904 24992 15932
rect 14240 15864 15148 15892
rect 14240 15852 14246 15864
rect 19334 15852 19340 15904
rect 19392 15852 19398 15904
rect 19426 15852 19432 15904
rect 19484 15852 19490 15904
rect 20809 15895 20867 15901
rect 20809 15861 20821 15895
rect 20855 15892 20867 15895
rect 20898 15892 20904 15904
rect 20855 15864 20904 15892
rect 20855 15861 20867 15864
rect 20809 15855 20867 15861
rect 20898 15852 20904 15864
rect 20956 15852 20962 15904
rect 21082 15852 21088 15904
rect 21140 15852 21146 15904
rect 24394 15852 24400 15904
rect 24452 15852 24458 15904
rect 24946 15852 24952 15904
rect 25004 15852 25010 15904
rect 25961 15895 26019 15901
rect 25961 15861 25973 15895
rect 26007 15892 26019 15895
rect 26050 15892 26056 15904
rect 26007 15864 26056 15892
rect 26007 15861 26019 15864
rect 25961 15855 26019 15861
rect 26050 15852 26056 15864
rect 26108 15852 26114 15904
rect 552 15802 27576 15824
rect 552 15750 7114 15802
rect 7166 15750 7178 15802
rect 7230 15750 7242 15802
rect 7294 15750 7306 15802
rect 7358 15750 7370 15802
rect 7422 15750 13830 15802
rect 13882 15750 13894 15802
rect 13946 15750 13958 15802
rect 14010 15750 14022 15802
rect 14074 15750 14086 15802
rect 14138 15750 20546 15802
rect 20598 15750 20610 15802
rect 20662 15750 20674 15802
rect 20726 15750 20738 15802
rect 20790 15750 20802 15802
rect 20854 15750 27262 15802
rect 27314 15750 27326 15802
rect 27378 15750 27390 15802
rect 27442 15750 27454 15802
rect 27506 15750 27518 15802
rect 27570 15750 27576 15802
rect 552 15728 27576 15750
rect 4525 15691 4583 15697
rect 4525 15657 4537 15691
rect 4571 15688 4583 15691
rect 4571 15660 5120 15688
rect 4571 15657 4583 15660
rect 4525 15651 4583 15657
rect 5092 15629 5120 15660
rect 6638 15648 6644 15700
rect 6696 15648 6702 15700
rect 6822 15648 6828 15700
rect 6880 15688 6886 15700
rect 7101 15691 7159 15697
rect 7101 15688 7113 15691
rect 6880 15660 7113 15688
rect 6880 15648 6886 15660
rect 7101 15657 7113 15660
rect 7147 15657 7159 15691
rect 7101 15651 7159 15657
rect 8846 15648 8852 15700
rect 8904 15648 8910 15700
rect 10502 15688 10508 15700
rect 9508 15660 10508 15688
rect 5077 15623 5135 15629
rect 5077 15589 5089 15623
rect 5123 15620 5135 15623
rect 5994 15620 6000 15632
rect 5123 15592 6000 15620
rect 5123 15589 5135 15592
rect 5077 15583 5135 15589
rect 5994 15580 6000 15592
rect 6052 15580 6058 15632
rect 7469 15623 7527 15629
rect 7469 15620 7481 15623
rect 6656 15592 7481 15620
rect 6656 15564 6684 15592
rect 7469 15589 7481 15592
rect 7515 15620 7527 15623
rect 8294 15620 8300 15632
rect 7515 15592 8300 15620
rect 7515 15589 7527 15592
rect 7469 15583 7527 15589
rect 8294 15580 8300 15592
rect 8352 15580 8358 15632
rect 9401 15623 9459 15629
rect 9401 15620 9413 15623
rect 8680 15592 9413 15620
rect 3418 15561 3424 15564
rect 3412 15515 3424 15561
rect 3418 15512 3424 15515
rect 3476 15512 3482 15564
rect 6457 15555 6515 15561
rect 6457 15521 6469 15555
rect 6503 15521 6515 15555
rect 6457 15515 6515 15521
rect 1394 15444 1400 15496
rect 1452 15484 1458 15496
rect 3145 15487 3203 15493
rect 3145 15484 3157 15487
rect 1452 15456 3157 15484
rect 1452 15444 1458 15456
rect 3145 15453 3157 15456
rect 3191 15453 3203 15487
rect 6472 15484 6500 15515
rect 6638 15512 6644 15564
rect 6696 15512 6702 15564
rect 7285 15555 7343 15561
rect 7285 15521 7297 15555
rect 7331 15550 7343 15555
rect 7374 15550 7380 15564
rect 7331 15522 7380 15550
rect 7331 15521 7343 15522
rect 7285 15515 7343 15521
rect 7374 15512 7380 15522
rect 7432 15512 7438 15564
rect 7561 15555 7619 15561
rect 7561 15521 7573 15555
rect 7607 15521 7619 15555
rect 7561 15515 7619 15521
rect 6822 15484 6828 15496
rect 6472 15456 6828 15484
rect 3145 15447 3203 15453
rect 6822 15444 6828 15456
rect 6880 15484 6886 15496
rect 7576 15484 7604 15515
rect 8478 15512 8484 15564
rect 8536 15512 8542 15564
rect 8680 15561 8708 15592
rect 9401 15589 9413 15592
rect 9447 15589 9459 15623
rect 9401 15583 9459 15589
rect 8665 15555 8723 15561
rect 8665 15521 8677 15555
rect 8711 15521 8723 15555
rect 8665 15515 8723 15521
rect 9125 15555 9183 15561
rect 9125 15521 9137 15555
rect 9171 15521 9183 15555
rect 9125 15515 9183 15521
rect 6880 15456 7604 15484
rect 9140 15484 9168 15515
rect 9306 15512 9312 15564
rect 9364 15552 9370 15564
rect 9508 15552 9536 15660
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 11974 15648 11980 15700
rect 12032 15688 12038 15700
rect 12032 15660 13483 15688
rect 12032 15648 12038 15660
rect 9600 15592 11468 15620
rect 9600 15561 9628 15592
rect 9364 15524 9536 15552
rect 9585 15555 9643 15561
rect 9364 15512 9370 15524
rect 9585 15521 9597 15555
rect 9631 15521 9643 15555
rect 9585 15515 9643 15521
rect 9674 15512 9680 15564
rect 9732 15512 9738 15564
rect 9766 15512 9772 15564
rect 9824 15512 9830 15564
rect 9907 15555 9965 15561
rect 9907 15521 9919 15555
rect 9953 15552 9965 15555
rect 10137 15555 10195 15561
rect 10137 15552 10149 15555
rect 9953 15524 10149 15552
rect 9953 15521 9965 15524
rect 9907 15515 9965 15521
rect 10137 15521 10149 15524
rect 10183 15521 10195 15555
rect 10321 15555 10379 15561
rect 10321 15552 10333 15555
rect 10137 15515 10195 15521
rect 10244 15524 10333 15552
rect 9490 15484 9496 15496
rect 9140 15456 9496 15484
rect 6880 15444 6886 15456
rect 7576 15416 7604 15456
rect 9490 15444 9496 15456
rect 9548 15484 9554 15496
rect 10045 15487 10103 15493
rect 10045 15484 10057 15487
rect 9548 15456 10057 15484
rect 9548 15444 9554 15456
rect 10045 15453 10057 15456
rect 10091 15453 10103 15487
rect 10045 15447 10103 15453
rect 9674 15416 9680 15428
rect 7576 15388 9680 15416
rect 9674 15376 9680 15388
rect 9732 15376 9738 15428
rect 9858 15376 9864 15428
rect 9916 15416 9922 15428
rect 10244 15416 10272 15524
rect 10321 15521 10333 15524
rect 10367 15552 10379 15555
rect 10502 15552 10508 15564
rect 10367 15524 10508 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 10502 15512 10508 15524
rect 10560 15512 10566 15564
rect 10597 15555 10655 15561
rect 10597 15521 10609 15555
rect 10643 15552 10655 15555
rect 10686 15552 10692 15564
rect 10643 15524 10692 15552
rect 10643 15521 10655 15524
rect 10597 15515 10655 15521
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 11440 15484 11468 15592
rect 12250 15512 12256 15564
rect 12308 15512 12314 15564
rect 12345 15555 12403 15561
rect 12345 15521 12357 15555
rect 12391 15552 12403 15555
rect 12452 15552 12480 15660
rect 12989 15623 13047 15629
rect 12989 15589 13001 15623
rect 13035 15620 13047 15623
rect 13326 15623 13384 15629
rect 13326 15620 13338 15623
rect 13035 15592 13338 15620
rect 13035 15589 13047 15592
rect 12989 15583 13047 15589
rect 13326 15589 13338 15592
rect 13372 15589 13384 15623
rect 13455 15620 13483 15660
rect 14182 15648 14188 15700
rect 14240 15688 14246 15700
rect 14461 15691 14519 15697
rect 14461 15688 14473 15691
rect 14240 15660 14473 15688
rect 14240 15648 14246 15660
rect 14461 15657 14473 15660
rect 14507 15657 14519 15691
rect 14461 15651 14519 15657
rect 18782 15648 18788 15700
rect 18840 15648 18846 15700
rect 20254 15648 20260 15700
rect 20312 15648 20318 15700
rect 20993 15691 21051 15697
rect 20993 15657 21005 15691
rect 21039 15688 21051 15691
rect 21039 15660 22094 15688
rect 21039 15657 21051 15660
rect 20993 15651 21051 15657
rect 14366 15620 14372 15632
rect 13455 15592 14372 15620
rect 13326 15583 13384 15589
rect 14366 15580 14372 15592
rect 14424 15620 14430 15632
rect 18874 15620 18880 15632
rect 14424 15592 18880 15620
rect 14424 15580 14430 15592
rect 18874 15580 18880 15592
rect 18932 15580 18938 15632
rect 19144 15623 19202 15629
rect 19144 15589 19156 15623
rect 19190 15620 19202 15623
rect 19426 15620 19432 15632
rect 19190 15592 19432 15620
rect 19190 15589 19202 15592
rect 19144 15583 19202 15589
rect 19426 15580 19432 15592
rect 19484 15580 19490 15632
rect 22066 15620 22094 15660
rect 22830 15648 22836 15700
rect 22888 15688 22894 15700
rect 23661 15691 23719 15697
rect 23661 15688 23673 15691
rect 22888 15660 23673 15688
rect 22888 15648 22894 15660
rect 23661 15657 23673 15660
rect 23707 15657 23719 15691
rect 23661 15651 23719 15657
rect 24486 15648 24492 15700
rect 24544 15648 24550 15700
rect 25685 15691 25743 15697
rect 25685 15657 25697 15691
rect 25731 15688 25743 15691
rect 25774 15688 25780 15700
rect 25731 15660 25780 15688
rect 25731 15657 25743 15660
rect 25685 15651 25743 15657
rect 25774 15648 25780 15660
rect 25832 15648 25838 15700
rect 22382 15623 22440 15629
rect 22382 15620 22394 15623
rect 20548 15592 21312 15620
rect 22066 15592 22394 15620
rect 12391 15524 12480 15552
rect 12391 15521 12403 15524
rect 12345 15515 12403 15521
rect 12526 15512 12532 15564
rect 12584 15512 12590 15564
rect 12621 15555 12679 15561
rect 12621 15521 12633 15555
rect 12667 15521 12679 15555
rect 12621 15515 12679 15521
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 13630 15552 13636 15564
rect 12759 15524 13636 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 12161 15487 12219 15493
rect 12161 15484 12173 15487
rect 11440 15456 12173 15484
rect 12161 15453 12173 15456
rect 12207 15453 12219 15487
rect 12161 15447 12219 15453
rect 9916 15388 10272 15416
rect 12176 15416 12204 15447
rect 12636 15416 12664 15515
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 16206 15512 16212 15564
rect 16264 15561 16270 15564
rect 16264 15555 16313 15561
rect 16264 15521 16267 15555
rect 16301 15521 16313 15555
rect 16264 15515 16313 15521
rect 16264 15512 16270 15515
rect 16390 15512 16396 15564
rect 16448 15512 16454 15564
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15521 16543 15555
rect 16666 15552 16672 15564
rect 16627 15524 16672 15552
rect 16485 15515 16543 15521
rect 12802 15444 12808 15496
rect 12860 15484 12866 15496
rect 13081 15487 13139 15493
rect 13081 15484 13093 15487
rect 12860 15456 13093 15484
rect 12860 15444 12866 15456
rect 13081 15453 13093 15456
rect 13127 15453 13139 15487
rect 16500 15484 16528 15515
rect 16666 15512 16672 15524
rect 16724 15512 16730 15564
rect 16758 15512 16764 15564
rect 16816 15512 16822 15564
rect 17672 15555 17730 15561
rect 17672 15521 17684 15555
rect 17718 15552 17730 15555
rect 18690 15552 18696 15564
rect 17718 15524 18696 15552
rect 17718 15521 17730 15524
rect 17672 15515 17730 15521
rect 18690 15512 18696 15524
rect 18748 15512 18754 15564
rect 19886 15512 19892 15564
rect 19944 15552 19950 15564
rect 20162 15552 20168 15564
rect 19944 15524 20168 15552
rect 19944 15512 19950 15524
rect 20162 15512 20168 15524
rect 20220 15552 20226 15564
rect 20548 15561 20576 15592
rect 20349 15555 20407 15561
rect 20349 15552 20361 15555
rect 20220 15524 20361 15552
rect 20220 15512 20226 15524
rect 20349 15521 20361 15524
rect 20395 15521 20407 15555
rect 20349 15515 20407 15521
rect 20533 15555 20591 15561
rect 20533 15521 20545 15555
rect 20579 15521 20591 15555
rect 20533 15515 20591 15521
rect 20625 15555 20683 15561
rect 20625 15521 20637 15555
rect 20671 15521 20683 15555
rect 20625 15515 20683 15521
rect 20717 15555 20775 15561
rect 20717 15521 20729 15555
rect 20763 15552 20775 15555
rect 21082 15552 21088 15564
rect 20763 15524 21088 15552
rect 20763 15521 20775 15524
rect 20717 15515 20775 15521
rect 16942 15484 16948 15496
rect 16500 15456 16948 15484
rect 13081 15447 13139 15453
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15453 17463 15487
rect 17405 15447 17463 15453
rect 18877 15487 18935 15493
rect 18877 15453 18889 15487
rect 18923 15453 18935 15487
rect 18877 15447 18935 15453
rect 12176 15388 12664 15416
rect 9916 15376 9922 15388
rect 4246 15308 4252 15360
rect 4304 15348 4310 15360
rect 5169 15351 5227 15357
rect 5169 15348 5181 15351
rect 4304 15320 5181 15348
rect 4304 15308 4310 15320
rect 5169 15317 5181 15320
rect 5215 15348 5227 15351
rect 6638 15348 6644 15360
rect 5215 15320 6644 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 9309 15351 9367 15357
rect 9309 15348 9321 15351
rect 8996 15320 9321 15348
rect 8996 15308 9002 15320
rect 9309 15317 9321 15320
rect 9355 15348 9367 15351
rect 9766 15348 9772 15360
rect 9355 15320 9772 15348
rect 9355 15317 9367 15320
rect 9309 15311 9367 15317
rect 9766 15308 9772 15320
rect 9824 15308 9830 15360
rect 15194 15308 15200 15360
rect 15252 15348 15258 15360
rect 16117 15351 16175 15357
rect 16117 15348 16129 15351
rect 15252 15320 16129 15348
rect 15252 15308 15258 15320
rect 16117 15317 16129 15320
rect 16163 15317 16175 15351
rect 17420 15348 17448 15447
rect 18892 15416 18920 15447
rect 20438 15444 20444 15496
rect 20496 15484 20502 15496
rect 20640 15484 20668 15515
rect 21082 15512 21088 15524
rect 21140 15512 21146 15564
rect 21284 15552 21312 15592
rect 22382 15589 22394 15592
rect 22428 15589 22440 15623
rect 22382 15583 22440 15589
rect 22646 15580 22652 15632
rect 22704 15620 22710 15632
rect 23017 15623 23075 15629
rect 23017 15620 23029 15623
rect 22704 15592 23029 15620
rect 22704 15580 22710 15592
rect 23017 15589 23029 15592
rect 23063 15589 23075 15623
rect 24504 15620 24532 15648
rect 23017 15583 23075 15589
rect 23308 15592 24532 15620
rect 24572 15623 24630 15629
rect 22554 15552 22560 15564
rect 21284 15524 22560 15552
rect 22554 15512 22560 15524
rect 22612 15512 22618 15564
rect 22922 15561 22928 15564
rect 22920 15552 22928 15561
rect 22883 15524 22928 15552
rect 22920 15515 22928 15524
rect 22922 15512 22928 15515
rect 22980 15512 22986 15564
rect 23106 15512 23112 15564
rect 23164 15512 23170 15564
rect 23308 15561 23336 15592
rect 24572 15589 24584 15623
rect 24618 15620 24630 15623
rect 25222 15620 25228 15632
rect 24618 15592 25228 15620
rect 24618 15589 24630 15592
rect 24572 15583 24630 15589
rect 25222 15580 25228 15592
rect 25280 15580 25286 15632
rect 23292 15555 23350 15561
rect 23292 15521 23304 15555
rect 23338 15521 23350 15555
rect 23292 15515 23350 15521
rect 23382 15512 23388 15564
rect 23440 15512 23446 15564
rect 23566 15512 23572 15564
rect 23624 15552 23630 15564
rect 23934 15552 23940 15564
rect 23624 15524 23940 15552
rect 23624 15512 23630 15524
rect 23934 15512 23940 15524
rect 23992 15512 23998 15564
rect 24854 15512 24860 15564
rect 24912 15552 24918 15564
rect 26973 15555 27031 15561
rect 26973 15552 26985 15555
rect 24912 15524 26985 15552
rect 24912 15512 24918 15524
rect 26973 15521 26985 15524
rect 27019 15521 27031 15555
rect 26973 15515 27031 15521
rect 20496 15456 20668 15484
rect 22649 15487 22707 15493
rect 20496 15444 20502 15456
rect 22649 15453 22661 15487
rect 22695 15484 22707 15487
rect 23474 15484 23480 15496
rect 22695 15456 23480 15484
rect 22695 15453 22707 15456
rect 22649 15447 22707 15453
rect 23474 15444 23480 15456
rect 23532 15484 23538 15496
rect 24305 15487 24363 15493
rect 24305 15484 24317 15487
rect 23532 15456 24317 15484
rect 23532 15444 23538 15456
rect 24305 15453 24317 15456
rect 24351 15453 24363 15487
rect 24305 15447 24363 15453
rect 18340 15388 18920 15416
rect 17770 15348 17776 15360
rect 17420 15320 17776 15348
rect 16117 15311 16175 15317
rect 17770 15308 17776 15320
rect 17828 15348 17834 15360
rect 18340 15348 18368 15388
rect 17828 15320 18368 15348
rect 21269 15351 21327 15357
rect 17828 15308 17834 15320
rect 21269 15317 21281 15351
rect 21315 15348 21327 15351
rect 21726 15348 21732 15360
rect 21315 15320 21732 15348
rect 21315 15317 21327 15320
rect 21269 15311 21327 15317
rect 21726 15308 21732 15320
rect 21784 15308 21790 15360
rect 22738 15308 22744 15360
rect 22796 15308 22802 15360
rect 24320 15348 24348 15447
rect 24670 15348 24676 15360
rect 24320 15320 24676 15348
rect 24670 15308 24676 15320
rect 24728 15308 24734 15360
rect 25774 15308 25780 15360
rect 25832 15348 25838 15360
rect 26421 15351 26479 15357
rect 26421 15348 26433 15351
rect 25832 15320 26433 15348
rect 25832 15308 25838 15320
rect 26421 15317 26433 15320
rect 26467 15317 26479 15351
rect 26421 15311 26479 15317
rect 552 15258 27416 15280
rect 552 15206 3756 15258
rect 3808 15206 3820 15258
rect 3872 15206 3884 15258
rect 3936 15206 3948 15258
rect 4000 15206 4012 15258
rect 4064 15206 10472 15258
rect 10524 15206 10536 15258
rect 10588 15206 10600 15258
rect 10652 15206 10664 15258
rect 10716 15206 10728 15258
rect 10780 15206 17188 15258
rect 17240 15206 17252 15258
rect 17304 15206 17316 15258
rect 17368 15206 17380 15258
rect 17432 15206 17444 15258
rect 17496 15206 23904 15258
rect 23956 15206 23968 15258
rect 24020 15206 24032 15258
rect 24084 15206 24096 15258
rect 24148 15206 24160 15258
rect 24212 15206 27416 15258
rect 552 15184 27416 15206
rect 4798 15104 4804 15156
rect 4856 15144 4862 15156
rect 4893 15147 4951 15153
rect 4893 15144 4905 15147
rect 4856 15116 4905 15144
rect 4856 15104 4862 15116
rect 4893 15113 4905 15116
rect 4939 15144 4951 15147
rect 5169 15147 5227 15153
rect 5169 15144 5181 15147
rect 4939 15116 5181 15144
rect 4939 15113 4951 15116
rect 4893 15107 4951 15113
rect 5169 15113 5181 15116
rect 5215 15113 5227 15147
rect 5169 15107 5227 15113
rect 5258 15104 5264 15156
rect 5316 15144 5322 15156
rect 5316 15116 5948 15144
rect 5316 15104 5322 15116
rect 4709 15079 4767 15085
rect 4709 15076 4721 15079
rect 4540 15048 4721 15076
rect 1394 14900 1400 14952
rect 1452 14940 1458 14952
rect 1673 14943 1731 14949
rect 1673 14940 1685 14943
rect 1452 14912 1685 14940
rect 1452 14900 1458 14912
rect 1673 14909 1685 14912
rect 1719 14909 1731 14943
rect 1673 14903 1731 14909
rect 4246 14900 4252 14952
rect 4304 14940 4310 14952
rect 4433 14943 4491 14949
rect 4433 14940 4445 14943
rect 4304 14912 4445 14940
rect 4304 14900 4310 14912
rect 4433 14909 4445 14912
rect 4479 14909 4491 14943
rect 4433 14903 4491 14909
rect 1940 14875 1998 14881
rect 1940 14841 1952 14875
rect 1986 14872 1998 14875
rect 4338 14872 4344 14884
rect 1986 14844 4344 14872
rect 1986 14841 1998 14844
rect 1940 14835 1998 14841
rect 4338 14832 4344 14844
rect 4396 14832 4402 14884
rect 3053 14807 3111 14813
rect 3053 14773 3065 14807
rect 3099 14804 3111 14807
rect 3786 14804 3792 14816
rect 3099 14776 3792 14804
rect 3099 14773 3111 14776
rect 3053 14767 3111 14773
rect 3786 14764 3792 14776
rect 3844 14804 3850 14816
rect 4540 14804 4568 15048
rect 4709 15045 4721 15048
rect 4755 15045 4767 15079
rect 5813 15079 5871 15085
rect 5813 15076 5825 15079
rect 4709 15039 4767 15045
rect 5552 15048 5825 15076
rect 5552 14952 5580 15048
rect 5813 15045 5825 15048
rect 5859 15045 5871 15079
rect 5920 15076 5948 15116
rect 5994 15104 6000 15156
rect 6052 15104 6058 15156
rect 6104 15116 9260 15144
rect 6104 15076 6132 15116
rect 5920 15048 6132 15076
rect 9125 15079 9183 15085
rect 5813 15039 5871 15045
rect 9125 15045 9137 15079
rect 9171 15045 9183 15079
rect 9232 15076 9260 15116
rect 9306 15104 9312 15156
rect 9364 15144 9370 15156
rect 9493 15147 9551 15153
rect 9493 15144 9505 15147
rect 9364 15116 9505 15144
rect 9364 15104 9370 15116
rect 9493 15113 9505 15116
rect 9539 15113 9551 15147
rect 9493 15107 9551 15113
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 10229 15147 10287 15153
rect 10229 15144 10241 15147
rect 9732 15116 10241 15144
rect 9732 15104 9738 15116
rect 10229 15113 10241 15116
rect 10275 15144 10287 15147
rect 10781 15147 10839 15153
rect 10275 15116 10456 15144
rect 10275 15113 10287 15116
rect 10229 15107 10287 15113
rect 10318 15076 10324 15088
rect 9232 15048 10324 15076
rect 9125 15039 9183 15045
rect 9140 15008 9168 15039
rect 10318 15036 10324 15048
rect 10376 15036 10382 15088
rect 9140 14980 9720 15008
rect 5350 14900 5356 14952
rect 5408 14900 5414 14952
rect 5534 14900 5540 14952
rect 5592 14900 5598 14952
rect 6365 14943 6423 14949
rect 6365 14940 6377 14943
rect 5736 14912 6377 14940
rect 5074 14832 5080 14884
rect 5132 14832 5138 14884
rect 5736 14813 5764 14912
rect 6365 14909 6377 14912
rect 6411 14909 6423 14943
rect 6365 14903 6423 14909
rect 6638 14900 6644 14952
rect 6696 14900 6702 14952
rect 6822 14900 6828 14952
rect 6880 14900 6886 14952
rect 9401 14943 9459 14949
rect 8220 14912 9352 14940
rect 8220 14884 8248 14912
rect 6181 14875 6239 14881
rect 6181 14841 6193 14875
rect 6227 14872 6239 14875
rect 8202 14872 8208 14884
rect 6227 14844 8208 14872
rect 6227 14841 6239 14844
rect 6181 14835 6239 14841
rect 8202 14832 8208 14844
rect 8260 14832 8266 14884
rect 8294 14832 8300 14884
rect 8352 14872 8358 14884
rect 8757 14875 8815 14881
rect 8757 14872 8769 14875
rect 8352 14844 8769 14872
rect 8352 14832 8358 14844
rect 8757 14841 8769 14844
rect 8803 14841 8815 14875
rect 9324 14872 9352 14912
rect 9401 14909 9413 14943
rect 9447 14940 9459 14943
rect 9490 14940 9496 14952
rect 9447 14912 9496 14940
rect 9447 14909 9459 14912
rect 9401 14903 9459 14909
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 9692 14949 9720 14980
rect 9677 14943 9735 14949
rect 9677 14909 9689 14943
rect 9723 14940 9735 14943
rect 9950 14940 9956 14952
rect 9723 14912 9956 14940
rect 9723 14909 9735 14912
rect 9677 14903 9735 14909
rect 9950 14900 9956 14912
rect 10008 14900 10014 14952
rect 10428 14949 10456 15116
rect 10781 15113 10793 15147
rect 10827 15144 10839 15147
rect 10870 15144 10876 15156
rect 10827 15116 10876 15144
rect 10827 15113 10839 15116
rect 10781 15107 10839 15113
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 12526 15104 12532 15156
rect 12584 15144 12590 15156
rect 13541 15147 13599 15153
rect 13541 15144 13553 15147
rect 12584 15116 13553 15144
rect 12584 15104 12590 15116
rect 13541 15113 13553 15116
rect 13587 15113 13599 15147
rect 13541 15107 13599 15113
rect 13725 15147 13783 15153
rect 13725 15113 13737 15147
rect 13771 15113 13783 15147
rect 13725 15107 13783 15113
rect 12250 15036 12256 15088
rect 12308 15076 12314 15088
rect 13740 15076 13768 15107
rect 16758 15104 16764 15156
rect 16816 15144 16822 15156
rect 18598 15144 18604 15156
rect 16816 15116 18604 15144
rect 16816 15104 16822 15116
rect 18598 15104 18604 15116
rect 18656 15104 18662 15156
rect 18690 15104 18696 15156
rect 18748 15104 18754 15156
rect 19260 15116 20484 15144
rect 12308 15048 13768 15076
rect 16301 15079 16359 15085
rect 12308 15036 12314 15048
rect 16301 15045 16313 15079
rect 16347 15076 16359 15079
rect 19260 15076 19288 15116
rect 16347 15048 17724 15076
rect 16347 15045 16359 15048
rect 16301 15039 16359 15045
rect 16206 14968 16212 15020
rect 16264 15008 16270 15020
rect 17696 15017 17724 15048
rect 18248 15048 19288 15076
rect 17681 15011 17739 15017
rect 16264 14980 17632 15008
rect 16264 14968 16270 14980
rect 10413 14943 10471 14949
rect 10413 14909 10425 14943
rect 10459 14909 10471 14943
rect 10413 14903 10471 14909
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 12986 14940 12992 14952
rect 12492 14912 12992 14940
rect 12492 14900 12498 14912
rect 12986 14900 12992 14912
rect 13044 14940 13050 14952
rect 13817 14943 13875 14949
rect 13817 14940 13829 14943
rect 13044 14912 13829 14940
rect 13044 14900 13050 14912
rect 13817 14909 13829 14912
rect 13863 14909 13875 14943
rect 13817 14903 13875 14909
rect 14093 14943 14151 14949
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 14182 14940 14188 14952
rect 14139 14912 14188 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 14182 14900 14188 14912
rect 14240 14900 14246 14952
rect 14921 14943 14979 14949
rect 14921 14909 14933 14943
rect 14967 14940 14979 14943
rect 14967 14912 15332 14940
rect 14967 14909 14979 14912
rect 14921 14903 14979 14909
rect 15304 14884 15332 14912
rect 15930 14900 15936 14952
rect 15988 14940 15994 14952
rect 16945 14943 17003 14949
rect 16945 14940 16957 14943
rect 15988 14912 16957 14940
rect 15988 14900 15994 14912
rect 16945 14909 16957 14912
rect 16991 14909 17003 14943
rect 17604 14940 17632 14980
rect 17681 14977 17693 15011
rect 17727 14977 17739 15011
rect 17681 14971 17739 14977
rect 18046 14949 18052 14952
rect 18003 14943 18052 14949
rect 18003 14940 18015 14943
rect 17604 14912 18015 14940
rect 16945 14903 17003 14909
rect 18003 14909 18015 14912
rect 18049 14909 18052 14943
rect 18003 14903 18052 14909
rect 18046 14900 18052 14903
rect 18104 14900 18110 14952
rect 10137 14875 10195 14881
rect 10137 14872 10149 14875
rect 9324 14844 10149 14872
rect 8757 14835 8815 14841
rect 10137 14841 10149 14844
rect 10183 14841 10195 14875
rect 10137 14835 10195 14841
rect 10318 14832 10324 14884
rect 10376 14872 10382 14884
rect 10597 14875 10655 14881
rect 10597 14872 10609 14875
rect 10376 14844 10609 14872
rect 10376 14832 10382 14844
rect 10597 14841 10609 14844
rect 10643 14841 10655 14875
rect 10597 14835 10655 14841
rect 15188 14875 15246 14881
rect 15188 14841 15200 14875
rect 15234 14841 15246 14875
rect 15188 14835 15246 14841
rect 3844 14776 4568 14804
rect 5721 14807 5779 14813
rect 3844 14764 3850 14776
rect 5721 14773 5733 14807
rect 5767 14773 5779 14807
rect 5721 14767 5779 14773
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 5971 14807 6029 14813
rect 5971 14804 5983 14807
rect 5868 14776 5983 14804
rect 5868 14764 5874 14776
rect 5971 14773 5983 14776
rect 6017 14773 6029 14807
rect 5971 14767 6029 14773
rect 6454 14764 6460 14816
rect 6512 14764 6518 14816
rect 6730 14764 6736 14816
rect 6788 14764 6794 14816
rect 8570 14764 8576 14816
rect 8628 14804 8634 14816
rect 9122 14804 9128 14816
rect 8628 14776 9128 14804
rect 8628 14764 8634 14776
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 9214 14764 9220 14816
rect 9272 14764 9278 14816
rect 9582 14764 9588 14816
rect 9640 14804 9646 14816
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9640 14776 9873 14804
rect 9640 14764 9646 14776
rect 9861 14773 9873 14776
rect 9907 14773 9919 14807
rect 15212 14804 15240 14835
rect 15286 14832 15292 14884
rect 15344 14832 15350 14884
rect 16393 14875 16451 14881
rect 16393 14872 16405 14875
rect 15396 14844 16405 14872
rect 15396 14804 15424 14844
rect 16393 14841 16405 14844
rect 16439 14841 16451 14875
rect 16393 14835 16451 14841
rect 17678 14832 17684 14884
rect 17736 14872 17742 14884
rect 17736 14844 18092 14872
rect 17736 14832 17742 14844
rect 15212 14776 15424 14804
rect 9861 14767 9919 14773
rect 15654 14764 15660 14816
rect 15712 14804 15718 14816
rect 16666 14804 16672 14816
rect 15712 14776 16672 14804
rect 15712 14764 15718 14776
rect 16666 14764 16672 14776
rect 16724 14804 16730 14816
rect 17129 14807 17187 14813
rect 17129 14804 17141 14807
rect 16724 14776 17141 14804
rect 16724 14764 16730 14776
rect 17129 14773 17141 14776
rect 17175 14773 17187 14807
rect 17129 14767 17187 14773
rect 17218 14764 17224 14816
rect 17276 14804 17282 14816
rect 17865 14807 17923 14813
rect 17865 14804 17877 14807
rect 17276 14776 17877 14804
rect 17276 14764 17282 14776
rect 17865 14773 17877 14776
rect 17911 14773 17923 14807
rect 18064 14804 18092 14844
rect 18138 14832 18144 14884
rect 18196 14832 18202 14884
rect 18248 14881 18276 15048
rect 19334 15036 19340 15088
rect 19392 15036 19398 15088
rect 20165 15079 20223 15085
rect 20165 15045 20177 15079
rect 20211 15045 20223 15079
rect 20165 15039 20223 15045
rect 18782 15008 18788 15020
rect 18432 14980 18788 15008
rect 18432 14949 18460 14980
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 19352 15008 19380 15036
rect 18984 14980 19380 15008
rect 18416 14943 18474 14949
rect 18416 14909 18428 14943
rect 18462 14909 18474 14943
rect 18416 14903 18474 14909
rect 18509 14943 18567 14949
rect 18509 14909 18521 14943
rect 18555 14940 18567 14943
rect 18598 14940 18604 14952
rect 18555 14912 18604 14940
rect 18555 14909 18567 14912
rect 18509 14903 18567 14909
rect 18598 14900 18604 14912
rect 18656 14900 18662 14952
rect 18984 14949 19012 14980
rect 19518 14968 19524 15020
rect 19576 14968 19582 15020
rect 20180 15008 20208 15039
rect 19996 14980 20208 15008
rect 18969 14943 19027 14949
rect 18969 14909 18981 14943
rect 19015 14909 19027 14943
rect 18969 14903 19027 14909
rect 19058 14900 19064 14952
rect 19116 14900 19122 14952
rect 19153 14943 19211 14949
rect 19153 14909 19165 14943
rect 19199 14909 19211 14943
rect 19153 14903 19211 14909
rect 19337 14943 19395 14949
rect 19337 14909 19349 14943
rect 19383 14940 19395 14943
rect 19886 14940 19892 14952
rect 19383 14912 19892 14940
rect 19383 14909 19395 14912
rect 19337 14903 19395 14909
rect 18233 14875 18291 14881
rect 18233 14841 18245 14875
rect 18279 14841 18291 14875
rect 19168 14872 19196 14903
rect 19886 14900 19892 14912
rect 19944 14900 19950 14952
rect 19996 14872 20024 14980
rect 20254 14900 20260 14952
rect 20312 14949 20318 14952
rect 20312 14943 20361 14949
rect 20312 14909 20315 14943
rect 20349 14909 20361 14943
rect 20456 14940 20484 15116
rect 24486 15104 24492 15156
rect 24544 15104 24550 15156
rect 26970 15144 26976 15156
rect 24596 15116 26976 15144
rect 24026 15036 24032 15088
rect 24084 15076 24090 15088
rect 24596 15076 24624 15116
rect 26970 15104 26976 15116
rect 27028 15104 27034 15156
rect 24084 15048 24624 15076
rect 24084 15036 24090 15048
rect 20898 15008 20904 15020
rect 20732 14980 20904 15008
rect 20732 14949 20760 14980
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 23474 15008 23480 15020
rect 22480 14980 23480 15008
rect 20533 14943 20591 14949
rect 20533 14940 20545 14943
rect 20456 14912 20545 14940
rect 20312 14903 20361 14909
rect 20533 14909 20545 14912
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 20716 14943 20774 14949
rect 20716 14909 20728 14943
rect 20762 14909 20774 14943
rect 20716 14903 20774 14909
rect 20312 14900 20318 14903
rect 19168 14844 20024 14872
rect 20441 14875 20499 14881
rect 18233 14835 18291 14841
rect 20441 14841 20453 14875
rect 20487 14841 20499 14875
rect 20548 14872 20576 14903
rect 20806 14900 20812 14952
rect 20864 14900 20870 14952
rect 21085 14943 21143 14949
rect 21085 14909 21097 14943
rect 21131 14940 21143 14943
rect 22480 14940 22508 14980
rect 23474 14968 23480 14980
rect 23532 14968 23538 15020
rect 21131 14912 22508 14940
rect 22557 14943 22615 14949
rect 21131 14909 21143 14912
rect 21085 14903 21143 14909
rect 22557 14909 22569 14943
rect 22603 14909 22615 14943
rect 22557 14903 22615 14909
rect 21174 14872 21180 14884
rect 20548 14844 21180 14872
rect 20441 14835 20499 14841
rect 18248 14804 18276 14835
rect 18064 14776 18276 14804
rect 17865 14767 17923 14773
rect 19334 14764 19340 14816
rect 19392 14804 19398 14816
rect 20073 14807 20131 14813
rect 20073 14804 20085 14807
rect 19392 14776 20085 14804
rect 19392 14764 19398 14776
rect 20073 14773 20085 14776
rect 20119 14804 20131 14807
rect 20456 14804 20484 14835
rect 21174 14832 21180 14844
rect 21232 14832 21238 14884
rect 21352 14875 21410 14881
rect 21352 14841 21364 14875
rect 21398 14872 21410 14875
rect 22002 14872 22008 14884
rect 21398 14844 22008 14872
rect 21398 14841 21410 14844
rect 21352 14835 21410 14841
rect 22002 14832 22008 14844
rect 22060 14832 22066 14884
rect 22572 14872 22600 14903
rect 24670 14900 24676 14952
rect 24728 14940 24734 14952
rect 25869 14943 25927 14949
rect 25869 14940 25881 14943
rect 24728 14912 25881 14940
rect 24728 14900 24734 14912
rect 25869 14909 25881 14912
rect 25915 14909 25927 14943
rect 25869 14903 25927 14909
rect 25958 14900 25964 14952
rect 26016 14940 26022 14952
rect 26513 14943 26571 14949
rect 26513 14940 26525 14943
rect 26016 14912 26525 14940
rect 26016 14900 26022 14912
rect 26513 14909 26525 14912
rect 26559 14909 26571 14943
rect 26513 14903 26571 14909
rect 22480 14844 22600 14872
rect 25624 14875 25682 14881
rect 22480 14813 22508 14844
rect 25624 14841 25636 14875
rect 25670 14872 25682 14875
rect 25774 14872 25780 14884
rect 25670 14844 25780 14872
rect 25670 14841 25682 14844
rect 25624 14835 25682 14841
rect 25774 14832 25780 14844
rect 25832 14832 25838 14884
rect 20119 14776 20484 14804
rect 22465 14807 22523 14813
rect 20119 14773 20131 14776
rect 20073 14767 20131 14773
rect 22465 14773 22477 14807
rect 22511 14773 22523 14807
rect 22465 14767 22523 14773
rect 23198 14764 23204 14816
rect 23256 14764 23262 14816
rect 25130 14764 25136 14816
rect 25188 14804 25194 14816
rect 25866 14804 25872 14816
rect 25188 14776 25872 14804
rect 25188 14764 25194 14776
rect 25866 14764 25872 14776
rect 25924 14804 25930 14816
rect 25961 14807 26019 14813
rect 25961 14804 25973 14807
rect 25924 14776 25973 14804
rect 25924 14764 25930 14776
rect 25961 14773 25973 14776
rect 26007 14773 26019 14807
rect 25961 14767 26019 14773
rect 552 14714 27576 14736
rect 552 14662 7114 14714
rect 7166 14662 7178 14714
rect 7230 14662 7242 14714
rect 7294 14662 7306 14714
rect 7358 14662 7370 14714
rect 7422 14662 13830 14714
rect 13882 14662 13894 14714
rect 13946 14662 13958 14714
rect 14010 14662 14022 14714
rect 14074 14662 14086 14714
rect 14138 14662 20546 14714
rect 20598 14662 20610 14714
rect 20662 14662 20674 14714
rect 20726 14662 20738 14714
rect 20790 14662 20802 14714
rect 20854 14662 27262 14714
rect 27314 14662 27326 14714
rect 27378 14662 27390 14714
rect 27442 14662 27454 14714
rect 27506 14662 27518 14714
rect 27570 14662 27576 14714
rect 552 14640 27576 14662
rect 3418 14560 3424 14612
rect 3476 14600 3482 14612
rect 3973 14603 4031 14609
rect 3973 14600 3985 14603
rect 3476 14572 3985 14600
rect 3476 14560 3482 14572
rect 3973 14569 3985 14572
rect 4019 14569 4031 14603
rect 3973 14563 4031 14569
rect 4338 14560 4344 14612
rect 4396 14600 4402 14612
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 4396 14572 4445 14600
rect 4396 14560 4402 14572
rect 4433 14569 4445 14572
rect 4479 14569 4491 14603
rect 5258 14600 5264 14612
rect 4433 14563 4491 14569
rect 4632 14572 5264 14600
rect 1940 14467 1998 14473
rect 1940 14433 1952 14467
rect 1986 14464 1998 14467
rect 3234 14464 3240 14476
rect 1986 14436 3240 14464
rect 1986 14433 1998 14436
rect 1940 14427 1998 14433
rect 3234 14424 3240 14436
rect 3292 14424 3298 14476
rect 3786 14424 3792 14476
rect 3844 14424 3850 14476
rect 4154 14424 4160 14476
rect 4212 14424 4218 14476
rect 4632 14473 4660 14572
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 5350 14560 5356 14612
rect 5408 14560 5414 14612
rect 6454 14560 6460 14612
rect 6512 14600 6518 14612
rect 9858 14600 9864 14612
rect 6512 14572 9864 14600
rect 6512 14560 6518 14572
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 9950 14560 9956 14612
rect 10008 14560 10014 14612
rect 11054 14560 11060 14612
rect 11112 14600 11118 14612
rect 11241 14603 11299 14609
rect 11241 14600 11253 14603
rect 11112 14572 11253 14600
rect 11112 14560 11118 14572
rect 11241 14569 11253 14572
rect 11287 14569 11299 14603
rect 11241 14563 11299 14569
rect 11348 14572 15884 14600
rect 5534 14532 5540 14544
rect 4908 14504 5540 14532
rect 4617 14467 4675 14473
rect 4617 14433 4629 14467
rect 4663 14433 4675 14467
rect 4617 14427 4675 14433
rect 4798 14424 4804 14476
rect 4856 14424 4862 14476
rect 4908 14473 4936 14504
rect 5534 14492 5540 14504
rect 5592 14492 5598 14544
rect 5994 14492 6000 14544
rect 6052 14532 6058 14544
rect 6822 14532 6828 14544
rect 6052 14504 6828 14532
rect 6052 14492 6058 14504
rect 6822 14492 6828 14504
rect 6880 14492 6886 14544
rect 7558 14492 7564 14544
rect 7616 14532 7622 14544
rect 8021 14535 8079 14541
rect 8021 14532 8033 14535
rect 7616 14504 8033 14532
rect 7616 14492 7622 14504
rect 8021 14501 8033 14504
rect 8067 14501 8079 14535
rect 8021 14495 8079 14501
rect 8237 14535 8295 14541
rect 8237 14501 8249 14535
rect 8283 14532 8295 14535
rect 8478 14532 8484 14544
rect 8283 14504 8484 14532
rect 8283 14501 8295 14504
rect 8237 14495 8295 14501
rect 8478 14492 8484 14504
rect 8536 14492 8542 14544
rect 8846 14541 8852 14544
rect 8840 14495 8852 14541
rect 8846 14492 8852 14495
rect 8904 14492 8910 14544
rect 4893 14467 4951 14473
rect 4893 14433 4905 14467
rect 4939 14433 4951 14467
rect 4893 14427 4951 14433
rect 5261 14467 5319 14473
rect 5261 14433 5273 14467
rect 5307 14433 5319 14467
rect 5261 14427 5319 14433
rect 5445 14467 5503 14473
rect 5445 14433 5457 14467
rect 5491 14464 5503 14467
rect 6270 14464 6276 14476
rect 5491 14436 6276 14464
rect 5491 14433 5503 14436
rect 5445 14427 5503 14433
rect 1394 14356 1400 14408
rect 1452 14396 1458 14408
rect 1673 14399 1731 14405
rect 1673 14396 1685 14399
rect 1452 14368 1685 14396
rect 1452 14356 1458 14368
rect 1673 14365 1685 14368
rect 1719 14365 1731 14399
rect 3804 14396 3832 14424
rect 5276 14396 5304 14427
rect 6270 14424 6276 14436
rect 6328 14424 6334 14476
rect 8570 14424 8576 14476
rect 8628 14424 8634 14476
rect 9858 14464 9864 14476
rect 8680 14436 9864 14464
rect 3804 14368 5304 14396
rect 1673 14359 1731 14365
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 7006 14396 7012 14408
rect 5408 14368 7012 14396
rect 5408 14356 5414 14368
rect 7006 14356 7012 14368
rect 7064 14356 7070 14408
rect 7466 14356 7472 14408
rect 7524 14396 7530 14408
rect 8680 14396 8708 14436
rect 9858 14424 9864 14436
rect 9916 14424 9922 14476
rect 9968 14464 9996 14560
rect 10042 14492 10048 14544
rect 10100 14532 10106 14544
rect 11348 14532 11376 14572
rect 10100 14504 11376 14532
rect 11609 14535 11667 14541
rect 10100 14492 10106 14504
rect 11609 14501 11621 14535
rect 11655 14532 11667 14535
rect 13262 14532 13268 14544
rect 11655 14504 13268 14532
rect 11655 14501 11667 14504
rect 11609 14495 11667 14501
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 10229 14467 10287 14473
rect 10229 14464 10241 14467
rect 9968 14436 10241 14464
rect 10229 14433 10241 14436
rect 10275 14433 10287 14467
rect 10229 14427 10287 14433
rect 10413 14467 10471 14473
rect 10413 14433 10425 14467
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 11701 14467 11759 14473
rect 11701 14433 11713 14467
rect 11747 14464 11759 14467
rect 12158 14464 12164 14476
rect 11747 14436 12164 14464
rect 11747 14433 11759 14436
rect 11701 14427 11759 14433
rect 10428 14396 10456 14427
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 14200 14473 14228 14572
rect 15194 14532 15200 14544
rect 14292 14504 15200 14532
rect 14292 14473 14320 14504
rect 15194 14492 15200 14504
rect 15252 14492 15258 14544
rect 15396 14504 15608 14532
rect 14093 14467 14151 14473
rect 14093 14433 14105 14467
rect 14139 14433 14151 14467
rect 14093 14427 14151 14433
rect 14185 14467 14243 14473
rect 14185 14433 14197 14467
rect 14231 14433 14243 14467
rect 14185 14427 14243 14433
rect 14277 14467 14335 14473
rect 14277 14433 14289 14467
rect 14323 14433 14335 14467
rect 14277 14427 14335 14433
rect 7524 14368 8708 14396
rect 9968 14368 10456 14396
rect 7524 14356 7530 14368
rect 7024 14328 7052 14356
rect 7024 14300 8616 14328
rect 3050 14220 3056 14272
rect 3108 14220 3114 14272
rect 3237 14263 3295 14269
rect 3237 14229 3249 14263
rect 3283 14260 3295 14263
rect 3418 14260 3424 14272
rect 3283 14232 3424 14260
rect 3283 14229 3295 14232
rect 3237 14223 3295 14229
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 8202 14220 8208 14272
rect 8260 14220 8266 14272
rect 8386 14220 8392 14272
rect 8444 14220 8450 14272
rect 8588 14260 8616 14300
rect 8754 14260 8760 14272
rect 8588 14232 8760 14260
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 8938 14220 8944 14272
rect 8996 14260 9002 14272
rect 9968 14260 9996 14368
rect 11330 14356 11336 14408
rect 11388 14396 11394 14408
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 11388 14368 11805 14396
rect 11388 14356 11394 14368
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 11882 14356 11888 14408
rect 11940 14396 11946 14408
rect 12805 14399 12863 14405
rect 12805 14396 12817 14399
rect 11940 14368 12817 14396
rect 11940 14356 11946 14368
rect 12805 14365 12817 14368
rect 12851 14365 12863 14399
rect 14108 14396 14136 14427
rect 14458 14424 14464 14476
rect 14516 14464 14522 14476
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 14516 14436 15301 14464
rect 14516 14424 14522 14436
rect 15289 14433 15301 14436
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 14108 14368 14565 14396
rect 12805 14359 12863 14365
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 15102 14356 15108 14408
rect 15160 14356 15166 14408
rect 8996 14232 9996 14260
rect 8996 14220 9002 14232
rect 10226 14220 10232 14272
rect 10284 14260 10290 14272
rect 10597 14263 10655 14269
rect 10597 14260 10609 14263
rect 10284 14232 10609 14260
rect 10284 14220 10290 14232
rect 10597 14229 10609 14232
rect 10643 14229 10655 14263
rect 10597 14223 10655 14229
rect 12250 14220 12256 14272
rect 12308 14220 12314 14272
rect 13814 14220 13820 14272
rect 13872 14220 13878 14272
rect 15396 14260 15424 14504
rect 15580 14473 15608 14504
rect 15473 14467 15531 14473
rect 15473 14433 15485 14467
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 15565 14467 15623 14473
rect 15565 14433 15577 14467
rect 15611 14433 15623 14467
rect 15565 14427 15623 14433
rect 15488 14396 15516 14427
rect 15654 14424 15660 14476
rect 15712 14424 15718 14476
rect 15856 14464 15884 14572
rect 15930 14560 15936 14612
rect 15988 14560 15994 14612
rect 16390 14560 16396 14612
rect 16448 14600 16454 14612
rect 16485 14603 16543 14609
rect 16485 14600 16497 14603
rect 16448 14572 16497 14600
rect 16448 14560 16454 14572
rect 16485 14569 16497 14572
rect 16531 14569 16543 14603
rect 16485 14563 16543 14569
rect 19245 14603 19303 14609
rect 19245 14569 19257 14603
rect 19291 14600 19303 14603
rect 19518 14600 19524 14612
rect 19291 14572 19524 14600
rect 19291 14569 19303 14572
rect 19245 14563 19303 14569
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 20070 14560 20076 14612
rect 20128 14560 20134 14612
rect 20162 14560 20168 14612
rect 20220 14600 20226 14612
rect 20714 14600 20720 14612
rect 20220 14572 20720 14600
rect 20220 14560 20226 14572
rect 20714 14560 20720 14572
rect 20772 14560 20778 14612
rect 21652 14572 22508 14600
rect 18046 14492 18052 14544
rect 18104 14532 18110 14544
rect 20898 14532 20904 14544
rect 18104 14504 20208 14532
rect 18104 14492 18110 14504
rect 20180 14476 20208 14504
rect 20364 14504 20904 14532
rect 16117 14467 16175 14473
rect 16117 14464 16129 14467
rect 15856 14436 16129 14464
rect 16117 14433 16129 14436
rect 16163 14433 16175 14467
rect 17218 14464 17224 14476
rect 16117 14427 16175 14433
rect 16224 14436 17224 14464
rect 16224 14396 16252 14436
rect 17218 14424 17224 14436
rect 17276 14424 17282 14476
rect 18132 14467 18190 14473
rect 18132 14433 18144 14467
rect 18178 14464 18190 14467
rect 19337 14467 19395 14473
rect 19337 14464 19349 14467
rect 18178 14436 19349 14464
rect 18178 14433 18190 14436
rect 18132 14427 18190 14433
rect 19337 14433 19349 14436
rect 19383 14433 19395 14467
rect 19337 14427 19395 14433
rect 20162 14424 20168 14476
rect 20220 14424 20226 14476
rect 20364 14473 20392 14504
rect 20898 14492 20904 14504
rect 20956 14492 20962 14544
rect 21174 14492 21180 14544
rect 21232 14532 21238 14544
rect 21652 14541 21680 14572
rect 21637 14535 21695 14541
rect 21637 14532 21649 14535
rect 21232 14504 21649 14532
rect 21232 14492 21238 14504
rect 21637 14501 21649 14504
rect 21683 14501 21695 14535
rect 22480 14532 22508 14572
rect 22554 14560 22560 14612
rect 22612 14600 22618 14612
rect 22741 14603 22799 14609
rect 22741 14600 22753 14603
rect 22612 14572 22753 14600
rect 22612 14560 22618 14572
rect 22741 14569 22753 14572
rect 22787 14569 22799 14603
rect 22741 14563 22799 14569
rect 24489 14603 24547 14609
rect 24489 14569 24501 14603
rect 24535 14600 24547 14603
rect 24854 14600 24860 14612
rect 24535 14572 24860 14600
rect 24535 14569 24547 14572
rect 24489 14563 24547 14569
rect 24854 14560 24860 14572
rect 24912 14560 24918 14612
rect 25317 14603 25375 14609
rect 25317 14569 25329 14603
rect 25363 14600 25375 14603
rect 25498 14600 25504 14612
rect 25363 14572 25504 14600
rect 25363 14569 25375 14572
rect 25317 14563 25375 14569
rect 25498 14560 25504 14572
rect 25556 14560 25562 14612
rect 25608 14572 26188 14600
rect 23106 14532 23112 14544
rect 21637 14495 21695 14501
rect 21744 14504 22140 14532
rect 22480 14504 23112 14532
rect 20349 14467 20407 14473
rect 20349 14433 20361 14467
rect 20395 14433 20407 14467
rect 20349 14427 20407 14433
rect 20438 14424 20444 14476
rect 20496 14424 20502 14476
rect 20533 14467 20591 14473
rect 20533 14433 20545 14467
rect 20579 14433 20591 14467
rect 20533 14427 20591 14433
rect 15488 14368 16252 14396
rect 16482 14356 16488 14408
rect 16540 14396 16546 14408
rect 17037 14399 17095 14405
rect 17037 14396 17049 14399
rect 16540 14368 17049 14396
rect 16540 14356 16546 14368
rect 17037 14365 17049 14368
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 17862 14356 17868 14408
rect 17920 14356 17926 14408
rect 19886 14356 19892 14408
rect 19944 14356 19950 14408
rect 20456 14328 20484 14424
rect 20548 14396 20576 14427
rect 20714 14424 20720 14476
rect 20772 14464 20778 14476
rect 20990 14464 20996 14476
rect 20772 14436 20996 14464
rect 20772 14424 20778 14436
rect 20990 14424 20996 14436
rect 21048 14424 21054 14476
rect 21448 14467 21506 14473
rect 21448 14433 21460 14467
rect 21494 14433 21506 14467
rect 21448 14427 21506 14433
rect 21463 14396 21491 14427
rect 21542 14424 21548 14476
rect 21600 14424 21606 14476
rect 21634 14396 21640 14408
rect 20548 14368 21312 14396
rect 21463 14368 21640 14396
rect 21284 14337 21312 14368
rect 21634 14356 21640 14368
rect 21692 14396 21698 14408
rect 21744 14396 21772 14504
rect 21818 14424 21824 14476
rect 21876 14424 21882 14476
rect 21910 14424 21916 14476
rect 21968 14424 21974 14476
rect 22112 14464 22140 14504
rect 23106 14492 23112 14504
rect 23164 14532 23170 14544
rect 23658 14532 23664 14544
rect 23164 14504 23664 14532
rect 23164 14492 23170 14504
rect 23658 14492 23664 14504
rect 23716 14492 23722 14544
rect 25608 14541 25636 14572
rect 25593 14535 25651 14541
rect 23860 14504 25268 14532
rect 22922 14473 22928 14476
rect 22920 14464 22928 14473
rect 22112 14436 22928 14464
rect 22920 14427 22928 14436
rect 22922 14424 22928 14427
rect 22980 14424 22986 14476
rect 23014 14424 23020 14476
rect 23072 14424 23078 14476
rect 23198 14424 23204 14476
rect 23256 14473 23262 14476
rect 23256 14467 23295 14473
rect 23283 14433 23295 14467
rect 23256 14427 23295 14433
rect 23256 14424 23262 14427
rect 23382 14424 23388 14476
rect 23440 14424 23446 14476
rect 23750 14424 23756 14476
rect 23808 14464 23814 14476
rect 23860 14473 23888 14504
rect 23845 14467 23903 14473
rect 23845 14464 23857 14467
rect 23808 14436 23857 14464
rect 23808 14424 23814 14436
rect 23845 14433 23857 14436
rect 23891 14433 23903 14467
rect 23845 14427 23903 14433
rect 24026 14424 24032 14476
rect 24084 14424 24090 14476
rect 24121 14467 24179 14473
rect 24121 14433 24133 14467
rect 24167 14433 24179 14467
rect 24121 14427 24179 14433
rect 24213 14467 24271 14473
rect 24213 14433 24225 14467
rect 24259 14464 24271 14467
rect 24394 14464 24400 14476
rect 24259 14436 24400 14464
rect 24259 14433 24271 14436
rect 24213 14427 24271 14433
rect 21692 14368 21772 14396
rect 21692 14356 21698 14368
rect 19076 14300 20484 14328
rect 19076 14272 19104 14300
rect 16301 14263 16359 14269
rect 16301 14260 16313 14263
rect 15396 14232 16313 14260
rect 16301 14229 16313 14232
rect 16347 14260 16359 14263
rect 19058 14260 19064 14272
rect 16347 14232 19064 14260
rect 16347 14229 16359 14232
rect 16301 14223 16359 14229
rect 19058 14220 19064 14232
rect 19116 14220 19122 14272
rect 20456 14260 20484 14300
rect 21269 14331 21327 14337
rect 21269 14297 21281 14331
rect 21315 14297 21327 14331
rect 21928 14328 21956 14424
rect 22002 14356 22008 14408
rect 22060 14356 22066 14408
rect 22278 14356 22284 14408
rect 22336 14396 22342 14408
rect 22557 14399 22615 14405
rect 22557 14396 22569 14399
rect 22336 14368 22569 14396
rect 22336 14356 22342 14368
rect 22557 14365 22569 14368
rect 22603 14365 22615 14399
rect 22557 14359 22615 14365
rect 23400 14328 23428 14424
rect 24136 14396 24164 14427
rect 24394 14424 24400 14436
rect 24452 14424 24458 14476
rect 24857 14467 24915 14473
rect 24857 14433 24869 14467
rect 24903 14433 24915 14467
rect 24857 14427 24915 14433
rect 24762 14396 24768 14408
rect 21928 14300 23428 14328
rect 23584 14368 24768 14396
rect 21269 14291 21327 14297
rect 22830 14260 22836 14272
rect 20456 14232 22836 14260
rect 22830 14220 22836 14232
rect 22888 14260 22894 14272
rect 23584 14260 23612 14368
rect 24762 14356 24768 14368
rect 24820 14356 24826 14408
rect 24872 14396 24900 14427
rect 24946 14424 24952 14476
rect 25004 14424 25010 14476
rect 25038 14424 25044 14476
rect 25096 14424 25102 14476
rect 25240 14473 25268 14504
rect 25593 14501 25605 14535
rect 25639 14501 25651 14535
rect 26160 14532 26188 14572
rect 26234 14560 26240 14612
rect 26292 14600 26298 14612
rect 27065 14603 27123 14609
rect 27065 14600 27077 14603
rect 26292 14572 27077 14600
rect 26292 14560 26298 14572
rect 27065 14569 27077 14572
rect 27111 14569 27123 14603
rect 27065 14563 27123 14569
rect 26326 14532 26332 14544
rect 26160 14504 26332 14532
rect 25593 14495 25651 14501
rect 26326 14492 26332 14504
rect 26384 14492 26390 14544
rect 25225 14467 25283 14473
rect 25225 14433 25237 14467
rect 25271 14464 25283 14467
rect 25314 14464 25320 14476
rect 25271 14436 25320 14464
rect 25271 14433 25283 14436
rect 25225 14427 25283 14433
rect 25314 14424 25320 14436
rect 25372 14424 25378 14476
rect 25498 14473 25504 14476
rect 25496 14464 25504 14473
rect 25459 14436 25504 14464
rect 25496 14427 25504 14436
rect 25498 14424 25504 14427
rect 25556 14424 25562 14476
rect 25685 14467 25743 14473
rect 25840 14467 25898 14473
rect 25972 14467 26030 14473
rect 25685 14464 25697 14467
rect 25608 14436 25697 14464
rect 25130 14396 25136 14408
rect 24872 14368 25136 14396
rect 25130 14356 25136 14368
rect 25188 14356 25194 14408
rect 23658 14288 23664 14340
rect 23716 14328 23722 14340
rect 25608 14328 25636 14436
rect 25685 14433 25697 14436
rect 25731 14433 25743 14467
rect 25685 14427 25743 14433
rect 25783 14439 25852 14467
rect 23716 14300 25636 14328
rect 25783 14328 25811 14439
rect 25840 14433 25852 14439
rect 25886 14436 25911 14467
rect 25886 14433 25898 14436
rect 25840 14427 25898 14433
rect 25972 14433 25984 14467
rect 26018 14464 26030 14467
rect 26418 14464 26424 14476
rect 26018 14436 26424 14464
rect 26018 14433 26030 14436
rect 25972 14427 26030 14433
rect 26418 14424 26424 14436
rect 26476 14424 26482 14476
rect 26602 14473 26608 14476
rect 26569 14467 26608 14473
rect 26569 14433 26581 14467
rect 26569 14427 26608 14433
rect 26602 14424 26608 14427
rect 26660 14424 26666 14476
rect 26694 14424 26700 14476
rect 26752 14424 26758 14476
rect 26786 14424 26792 14476
rect 26844 14424 26850 14476
rect 26878 14424 26884 14476
rect 26936 14473 26942 14476
rect 26936 14464 26944 14473
rect 26936 14436 26981 14464
rect 26936 14427 26944 14436
rect 26936 14424 26942 14427
rect 26712 14396 26740 14424
rect 26620 14368 26740 14396
rect 25866 14328 25872 14340
rect 25783 14300 25872 14328
rect 23716 14288 23722 14300
rect 22888 14232 23612 14260
rect 22888 14220 22894 14232
rect 24578 14220 24584 14272
rect 24636 14220 24642 14272
rect 25608 14260 25636 14300
rect 25866 14288 25872 14300
rect 25924 14288 25930 14340
rect 26510 14260 26516 14272
rect 25608 14232 26516 14260
rect 26510 14220 26516 14232
rect 26568 14260 26574 14272
rect 26620 14260 26648 14368
rect 26568 14232 26648 14260
rect 26568 14220 26574 14232
rect 552 14170 27416 14192
rect 552 14118 3756 14170
rect 3808 14118 3820 14170
rect 3872 14118 3884 14170
rect 3936 14118 3948 14170
rect 4000 14118 4012 14170
rect 4064 14118 10472 14170
rect 10524 14118 10536 14170
rect 10588 14118 10600 14170
rect 10652 14118 10664 14170
rect 10716 14118 10728 14170
rect 10780 14118 17188 14170
rect 17240 14118 17252 14170
rect 17304 14118 17316 14170
rect 17368 14118 17380 14170
rect 17432 14118 17444 14170
rect 17496 14118 23904 14170
rect 23956 14118 23968 14170
rect 24020 14118 24032 14170
rect 24084 14118 24096 14170
rect 24148 14118 24160 14170
rect 24212 14118 27416 14170
rect 552 14096 27416 14118
rect 3234 14016 3240 14068
rect 3292 14016 3298 14068
rect 4065 14059 4123 14065
rect 4065 14025 4077 14059
rect 4111 14056 4123 14059
rect 4430 14056 4436 14068
rect 4111 14028 4436 14056
rect 4111 14025 4123 14028
rect 4065 14019 4123 14025
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 4525 14059 4583 14065
rect 4525 14025 4537 14059
rect 4571 14056 4583 14059
rect 5810 14056 5816 14068
rect 4571 14028 5816 14056
rect 4571 14025 4583 14028
rect 4525 14019 4583 14025
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 9769 14059 9827 14065
rect 9769 14056 9781 14059
rect 8260 14028 9781 14056
rect 8260 14016 8266 14028
rect 9769 14025 9781 14028
rect 9815 14056 9827 14059
rect 9861 14059 9919 14065
rect 9861 14056 9873 14059
rect 9815 14028 9873 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 9861 14025 9873 14028
rect 9907 14056 9919 14059
rect 11330 14056 11336 14068
rect 9907 14028 11336 14056
rect 9907 14025 9919 14028
rect 9861 14019 9919 14025
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 12802 14056 12808 14068
rect 11440 14028 12808 14056
rect 3326 13948 3332 14000
rect 3384 13988 3390 14000
rect 4249 13991 4307 13997
rect 3384 13960 3556 13988
rect 3384 13948 3390 13960
rect 3418 13880 3424 13932
rect 3476 13880 3482 13932
rect 3528 13920 3556 13960
rect 4249 13957 4261 13991
rect 4295 13957 4307 13991
rect 4249 13951 4307 13957
rect 3605 13923 3663 13929
rect 3605 13920 3617 13923
rect 3528 13892 3617 13920
rect 3605 13889 3617 13892
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 3697 13923 3755 13929
rect 3697 13889 3709 13923
rect 3743 13920 3755 13923
rect 4264 13920 4292 13951
rect 4338 13948 4344 14000
rect 4396 13948 4402 14000
rect 5445 13991 5503 13997
rect 5445 13957 5457 13991
rect 5491 13988 5503 13991
rect 5905 13991 5963 13997
rect 5905 13988 5917 13991
rect 5491 13960 5917 13988
rect 5491 13957 5503 13960
rect 5445 13951 5503 13957
rect 5905 13957 5917 13960
rect 5951 13957 5963 13991
rect 5905 13951 5963 13957
rect 4522 13920 4528 13932
rect 3743 13892 4528 13920
rect 3743 13889 3755 13892
rect 3697 13883 3755 13889
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 6089 13923 6147 13929
rect 6089 13920 6101 13923
rect 5132 13892 6101 13920
rect 5132 13880 5138 13892
rect 6089 13889 6101 13892
rect 6135 13889 6147 13923
rect 6089 13883 6147 13889
rect 6457 13923 6515 13929
rect 6457 13889 6469 13923
rect 6503 13920 6515 13923
rect 7193 13923 7251 13929
rect 7193 13920 7205 13923
rect 6503 13892 7205 13920
rect 6503 13889 6515 13892
rect 6457 13883 6515 13889
rect 7193 13889 7205 13892
rect 7239 13889 7251 13923
rect 7193 13883 7251 13889
rect 3510 13812 3516 13864
rect 3568 13852 3574 13864
rect 4246 13852 4252 13864
rect 3568 13824 4252 13852
rect 3568 13812 3574 13824
rect 4246 13812 4252 13824
rect 4304 13852 4310 13864
rect 4304 13824 4752 13852
rect 4304 13812 4310 13824
rect 3050 13744 3056 13796
rect 3108 13784 3114 13796
rect 4522 13793 4528 13796
rect 3881 13787 3939 13793
rect 3881 13784 3893 13787
rect 3108 13756 3893 13784
rect 3108 13744 3114 13756
rect 3881 13753 3893 13756
rect 3927 13784 3939 13787
rect 4493 13787 4528 13793
rect 3927 13756 4384 13784
rect 3927 13753 3939 13756
rect 3881 13747 3939 13753
rect 4062 13676 4068 13728
rect 4120 13725 4126 13728
rect 4120 13719 4139 13725
rect 4127 13685 4139 13719
rect 4356 13716 4384 13756
rect 4493 13753 4505 13787
rect 4493 13747 4528 13753
rect 4522 13744 4528 13747
rect 4580 13744 4586 13796
rect 4724 13793 4752 13824
rect 5258 13812 5264 13864
rect 5316 13812 5322 13864
rect 5537 13855 5595 13861
rect 5537 13821 5549 13855
rect 5583 13821 5595 13855
rect 5537 13815 5595 13821
rect 4709 13787 4767 13793
rect 4709 13753 4721 13787
rect 4755 13784 4767 13787
rect 5552 13784 5580 13815
rect 5626 13812 5632 13864
rect 5684 13812 5690 13864
rect 5905 13855 5963 13861
rect 5905 13821 5917 13855
rect 5951 13852 5963 13855
rect 5994 13852 6000 13864
rect 5951 13824 6000 13852
rect 5951 13821 5963 13824
rect 5905 13815 5963 13821
rect 5994 13812 6000 13824
rect 6052 13812 6058 13864
rect 6104 13852 6132 13883
rect 7466 13880 7472 13932
rect 7524 13880 7530 13932
rect 7742 13880 7748 13932
rect 7800 13920 7806 13932
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 7800 13892 8401 13920
rect 7800 13880 7806 13892
rect 8389 13889 8401 13892
rect 8435 13889 8447 13923
rect 8389 13883 8447 13889
rect 9398 13880 9404 13932
rect 9456 13920 9462 13932
rect 11440 13929 11468 14028
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 14921 14059 14979 14065
rect 14921 14025 14933 14059
rect 14967 14056 14979 14059
rect 15102 14056 15108 14068
rect 14967 14028 15108 14056
rect 14967 14025 14979 14028
rect 14921 14019 14979 14025
rect 15102 14016 15108 14028
rect 15160 14016 15166 14068
rect 16482 14016 16488 14068
rect 16540 14016 16546 14068
rect 17494 14016 17500 14068
rect 17552 14056 17558 14068
rect 18693 14059 18751 14065
rect 18693 14056 18705 14059
rect 17552 14028 18705 14056
rect 17552 14016 17558 14028
rect 18693 14025 18705 14028
rect 18739 14025 18751 14059
rect 18693 14019 18751 14025
rect 18782 14016 18788 14068
rect 18840 14056 18846 14068
rect 20349 14059 20407 14065
rect 20349 14056 20361 14059
rect 18840 14028 20361 14056
rect 18840 14016 18846 14028
rect 20349 14025 20361 14028
rect 20395 14056 20407 14059
rect 21634 14056 21640 14068
rect 20395 14028 21640 14056
rect 20395 14025 20407 14028
rect 20349 14019 20407 14025
rect 21634 14016 21640 14028
rect 21692 14016 21698 14068
rect 22278 14016 22284 14068
rect 22336 14016 22342 14068
rect 23198 14056 23204 14068
rect 22572 14028 23204 14056
rect 18138 13948 18144 14000
rect 18196 13988 18202 14000
rect 18509 13991 18567 13997
rect 18509 13988 18521 13991
rect 18196 13960 18521 13988
rect 18196 13948 18202 13960
rect 18509 13957 18521 13960
rect 18555 13988 18567 13991
rect 21542 13988 21548 14000
rect 18555 13960 19555 13988
rect 18555 13957 18567 13960
rect 18509 13951 18567 13957
rect 11425 13923 11483 13929
rect 11425 13920 11437 13923
rect 9456 13892 11437 13920
rect 9456 13880 9462 13892
rect 11425 13889 11437 13892
rect 11471 13889 11483 13923
rect 11425 13883 11483 13889
rect 12802 13880 12808 13932
rect 12860 13920 12866 13932
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 12860 13892 13553 13920
rect 12860 13880 12866 13892
rect 13541 13889 13553 13892
rect 13587 13889 13599 13923
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 13541 13883 13599 13889
rect 18432 13892 19441 13920
rect 6104 13824 6224 13852
rect 4755 13756 5580 13784
rect 6196 13784 6224 13824
rect 6270 13812 6276 13864
rect 6328 13852 6334 13864
rect 8662 13861 8668 13864
rect 6549 13855 6607 13861
rect 6549 13852 6561 13855
rect 6328 13824 6561 13852
rect 6328 13812 6334 13824
rect 6549 13821 6561 13824
rect 6595 13821 6607 13855
rect 6733 13855 6791 13861
rect 6733 13852 6745 13855
rect 6549 13815 6607 13821
rect 6656 13824 6745 13852
rect 6656 13784 6684 13824
rect 6733 13821 6745 13824
rect 6779 13821 6791 13855
rect 6733 13815 6791 13821
rect 8656 13815 8668 13861
rect 8662 13812 8668 13815
rect 8720 13812 8726 13864
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 9640 13824 9873 13852
rect 9640 13812 9646 13824
rect 9861 13821 9873 13824
rect 9907 13821 9919 13855
rect 9861 13815 9919 13821
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13852 10103 13855
rect 10318 13852 10324 13864
rect 10091 13824 10324 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 6196 13756 6684 13784
rect 6917 13787 6975 13793
rect 4755 13753 4767 13756
rect 4709 13747 4767 13753
rect 6917 13753 6929 13787
rect 6963 13784 6975 13787
rect 8202 13784 8208 13796
rect 6963 13756 8208 13784
rect 6963 13753 6975 13756
rect 6917 13747 6975 13753
rect 8202 13744 8208 13756
rect 8260 13744 8266 13796
rect 10060 13784 10088 13815
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 11692 13855 11750 13861
rect 11692 13821 11704 13855
rect 11738 13852 11750 13855
rect 12250 13852 12256 13864
rect 11738 13824 12256 13852
rect 11738 13821 11750 13824
rect 11692 13815 11750 13821
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 13814 13861 13820 13864
rect 13808 13852 13820 13861
rect 13775 13824 13820 13852
rect 13808 13815 13820 13824
rect 13814 13812 13820 13815
rect 13872 13812 13878 13864
rect 15105 13855 15163 13861
rect 15105 13821 15117 13855
rect 15151 13852 15163 13855
rect 15194 13852 15200 13864
rect 15151 13824 15200 13852
rect 15151 13821 15163 13824
rect 15105 13815 15163 13821
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17862 13852 17868 13864
rect 17175 13824 17868 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 18432 13852 18460 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 17972 13824 18460 13852
rect 19337 13855 19395 13861
rect 14366 13784 14372 13796
rect 8680 13756 10088 13784
rect 10244 13756 14372 13784
rect 5721 13719 5779 13725
rect 5721 13716 5733 13719
rect 4356 13688 5733 13716
rect 4120 13679 4139 13685
rect 5721 13685 5733 13688
rect 5767 13716 5779 13719
rect 6638 13716 6644 13728
rect 5767 13688 6644 13716
rect 5767 13685 5779 13688
rect 5721 13679 5779 13685
rect 4120 13676 4126 13679
rect 6638 13676 6644 13688
rect 6696 13716 6702 13728
rect 8680 13716 8708 13756
rect 6696 13688 8708 13716
rect 6696 13676 6702 13688
rect 8754 13676 8760 13728
rect 8812 13716 8818 13728
rect 9398 13716 9404 13728
rect 8812 13688 9404 13716
rect 8812 13676 8818 13688
rect 9398 13676 9404 13688
rect 9456 13676 9462 13728
rect 9490 13676 9496 13728
rect 9548 13716 9554 13728
rect 10244 13725 10272 13756
rect 14366 13744 14372 13756
rect 14424 13744 14430 13796
rect 15372 13787 15430 13793
rect 15372 13753 15384 13787
rect 15418 13784 15430 13787
rect 16114 13784 16120 13796
rect 15418 13756 16120 13784
rect 15418 13753 15430 13756
rect 15372 13747 15430 13753
rect 16114 13744 16120 13756
rect 16172 13744 16178 13796
rect 17396 13787 17454 13793
rect 17396 13753 17408 13787
rect 17442 13784 17454 13787
rect 17972 13784 18000 13824
rect 19337 13821 19349 13855
rect 19383 13852 19395 13855
rect 19527 13852 19555 13960
rect 21468 13960 21548 13988
rect 21468 13929 21496 13960
rect 21542 13948 21548 13960
rect 21600 13948 21606 14000
rect 21453 13923 21511 13929
rect 21453 13889 21465 13923
rect 21499 13889 21511 13923
rect 21453 13883 21511 13889
rect 19383 13824 19555 13852
rect 19383 13821 19395 13824
rect 19337 13815 19395 13821
rect 19702 13812 19708 13864
rect 19760 13852 19766 13864
rect 19981 13855 20039 13861
rect 19981 13852 19993 13855
rect 19760 13824 19993 13852
rect 19760 13812 19766 13824
rect 19981 13821 19993 13824
rect 20027 13821 20039 13855
rect 19981 13815 20039 13821
rect 20162 13812 20168 13864
rect 20220 13812 20226 13864
rect 21082 13812 21088 13864
rect 21140 13852 21146 13864
rect 22572 13861 22600 14028
rect 23198 14016 23204 14028
rect 23256 14016 23262 14068
rect 23382 14016 23388 14068
rect 23440 14056 23446 14068
rect 26418 14056 26424 14068
rect 23440 14028 26424 14056
rect 23440 14016 23446 14028
rect 26418 14016 26424 14028
rect 26476 14016 26482 14068
rect 26602 14016 26608 14068
rect 26660 14056 26666 14068
rect 26881 14059 26939 14065
rect 26881 14056 26893 14059
rect 26660 14028 26893 14056
rect 26660 14016 26666 14028
rect 26881 14025 26893 14028
rect 26927 14025 26939 14059
rect 26881 14019 26939 14025
rect 24578 13988 24584 14000
rect 23124 13960 24584 13988
rect 22830 13920 22836 13932
rect 22664 13892 22836 13920
rect 22664 13861 22692 13892
rect 22830 13880 22836 13892
rect 22888 13880 22894 13932
rect 23124 13929 23152 13960
rect 24578 13948 24584 13960
rect 24636 13948 24642 14000
rect 23109 13923 23167 13929
rect 23109 13889 23121 13923
rect 23155 13889 23167 13923
rect 23109 13883 23167 13889
rect 23661 13923 23719 13929
rect 23661 13889 23673 13923
rect 23707 13920 23719 13923
rect 24854 13920 24860 13932
rect 23707 13892 24860 13920
rect 23707 13889 23719 13892
rect 23661 13883 23719 13889
rect 24854 13880 24860 13892
rect 24912 13880 24918 13932
rect 21545 13855 21603 13861
rect 21545 13852 21557 13855
rect 21140 13824 21557 13852
rect 21140 13812 21146 13824
rect 21545 13821 21557 13824
rect 21591 13821 21603 13855
rect 21545 13815 21603 13821
rect 22557 13855 22615 13861
rect 22557 13821 22569 13855
rect 22603 13821 22615 13855
rect 22557 13815 22615 13821
rect 22649 13855 22707 13861
rect 22649 13821 22661 13855
rect 22695 13821 22707 13855
rect 22649 13815 22707 13821
rect 22738 13812 22744 13864
rect 22796 13812 22802 13864
rect 22925 13855 22983 13861
rect 22925 13852 22937 13855
rect 22848 13824 22937 13852
rect 17442 13756 18000 13784
rect 17442 13753 17454 13756
rect 17396 13747 17454 13753
rect 18230 13744 18236 13796
rect 18288 13784 18294 13796
rect 19426 13784 19432 13796
rect 18288 13756 19432 13784
rect 18288 13744 18294 13756
rect 19426 13744 19432 13756
rect 19484 13744 19490 13796
rect 20990 13744 20996 13796
rect 21048 13784 21054 13796
rect 22848 13784 22876 13824
rect 22925 13821 22937 13824
rect 22971 13852 22983 13855
rect 23750 13852 23756 13864
rect 22971 13824 23756 13852
rect 22971 13821 22983 13824
rect 22925 13815 22983 13821
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 24489 13855 24547 13861
rect 24489 13821 24501 13855
rect 24535 13821 24547 13855
rect 24489 13815 24547 13821
rect 21048 13756 22876 13784
rect 24504 13784 24532 13815
rect 24578 13812 24584 13864
rect 24636 13812 24642 13864
rect 24670 13812 24676 13864
rect 24728 13852 24734 13864
rect 25501 13855 25559 13861
rect 25501 13852 25513 13855
rect 24728 13824 25513 13852
rect 24728 13812 24734 13824
rect 25501 13821 25513 13824
rect 25547 13821 25559 13855
rect 25501 13815 25559 13821
rect 25768 13855 25826 13861
rect 25768 13821 25780 13855
rect 25814 13852 25826 13855
rect 26050 13852 26056 13864
rect 25814 13824 26056 13852
rect 25814 13821 25826 13824
rect 25768 13815 25826 13821
rect 26050 13812 26056 13824
rect 26108 13812 26114 13864
rect 25866 13784 25872 13796
rect 24504 13756 25872 13784
rect 21048 13744 21054 13756
rect 25866 13744 25872 13756
rect 25924 13744 25930 13796
rect 10229 13719 10287 13725
rect 10229 13716 10241 13719
rect 9548 13688 10241 13716
rect 9548 13676 9554 13688
rect 10229 13685 10241 13688
rect 10275 13685 10287 13719
rect 10229 13679 10287 13685
rect 12805 13719 12863 13725
rect 12805 13685 12817 13719
rect 12851 13716 12863 13719
rect 13170 13716 13176 13728
rect 12851 13688 13176 13716
rect 12851 13685 12863 13688
rect 12805 13679 12863 13685
rect 13170 13676 13176 13688
rect 13228 13676 13234 13728
rect 14274 13676 14280 13728
rect 14332 13716 14338 13728
rect 16206 13716 16212 13728
rect 14332 13688 16212 13716
rect 14332 13676 14338 13688
rect 16206 13676 16212 13688
rect 16264 13676 16270 13728
rect 18782 13676 18788 13728
rect 18840 13716 18846 13728
rect 19702 13716 19708 13728
rect 18840 13688 19708 13716
rect 18840 13676 18846 13688
rect 19702 13676 19708 13688
rect 19760 13676 19766 13728
rect 20809 13719 20867 13725
rect 20809 13685 20821 13719
rect 20855 13716 20867 13719
rect 20898 13716 20904 13728
rect 20855 13688 20904 13716
rect 20855 13685 20867 13688
rect 20809 13679 20867 13685
rect 20898 13676 20904 13688
rect 20956 13676 20962 13728
rect 22186 13676 22192 13728
rect 22244 13676 22250 13728
rect 23842 13676 23848 13728
rect 23900 13676 23906 13728
rect 25225 13719 25283 13725
rect 25225 13685 25237 13719
rect 25271 13716 25283 13719
rect 25682 13716 25688 13728
rect 25271 13688 25688 13716
rect 25271 13685 25283 13688
rect 25225 13679 25283 13685
rect 25682 13676 25688 13688
rect 25740 13676 25746 13728
rect 552 13626 27576 13648
rect 552 13574 7114 13626
rect 7166 13574 7178 13626
rect 7230 13574 7242 13626
rect 7294 13574 7306 13626
rect 7358 13574 7370 13626
rect 7422 13574 13830 13626
rect 13882 13574 13894 13626
rect 13946 13574 13958 13626
rect 14010 13574 14022 13626
rect 14074 13574 14086 13626
rect 14138 13574 20546 13626
rect 20598 13574 20610 13626
rect 20662 13574 20674 13626
rect 20726 13574 20738 13626
rect 20790 13574 20802 13626
rect 20854 13574 27262 13626
rect 27314 13574 27326 13626
rect 27378 13574 27390 13626
rect 27442 13574 27454 13626
rect 27506 13574 27518 13626
rect 27570 13574 27576 13626
rect 552 13552 27576 13574
rect 4065 13515 4123 13521
rect 4065 13481 4077 13515
rect 4111 13512 4123 13515
rect 4154 13512 4160 13524
rect 4111 13484 4160 13512
rect 4111 13481 4123 13484
rect 4065 13475 4123 13481
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 4246 13472 4252 13524
rect 4304 13512 4310 13524
rect 4617 13515 4675 13521
rect 4304 13484 4568 13512
rect 4304 13472 4310 13484
rect 3421 13447 3479 13453
rect 3421 13413 3433 13447
rect 3467 13444 3479 13447
rect 3510 13444 3516 13456
rect 3467 13416 3516 13444
rect 3467 13413 3479 13416
rect 3421 13407 3479 13413
rect 3510 13404 3516 13416
rect 3568 13404 3574 13456
rect 4540 13444 4568 13484
rect 4617 13481 4629 13515
rect 4663 13512 4675 13515
rect 4706 13512 4712 13524
rect 4663 13484 4712 13512
rect 4663 13481 4675 13484
rect 4617 13475 4675 13481
rect 4706 13472 4712 13484
rect 4764 13512 4770 13524
rect 5258 13512 5264 13524
rect 4764 13484 5264 13512
rect 4764 13472 4770 13484
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 6270 13472 6276 13524
rect 6328 13472 6334 13524
rect 8478 13472 8484 13524
rect 8536 13472 8542 13524
rect 8573 13515 8631 13521
rect 8573 13481 8585 13515
rect 8619 13512 8631 13515
rect 8662 13512 8668 13524
rect 8619 13484 8668 13512
rect 8619 13481 8631 13484
rect 8573 13475 8631 13481
rect 8662 13472 8668 13484
rect 8720 13472 8726 13524
rect 8846 13472 8852 13524
rect 8904 13512 8910 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8904 13484 8953 13512
rect 8904 13472 8910 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 8941 13475 8999 13481
rect 11609 13515 11667 13521
rect 11609 13481 11621 13515
rect 11655 13481 11667 13515
rect 11609 13475 11667 13481
rect 4540 13416 4752 13444
rect 3786 13336 3792 13388
rect 3844 13336 3850 13388
rect 3881 13379 3939 13385
rect 3881 13345 3893 13379
rect 3927 13345 3939 13379
rect 3881 13339 3939 13345
rect 4157 13379 4215 13385
rect 4157 13345 4169 13379
rect 4203 13374 4215 13379
rect 4338 13376 4344 13388
rect 4264 13374 4344 13376
rect 4203 13348 4344 13374
rect 4203 13346 4292 13348
rect 4203 13345 4215 13346
rect 4157 13339 4215 13345
rect 3234 13268 3240 13320
rect 3292 13268 3298 13320
rect 3896 13240 3924 13339
rect 4338 13336 4344 13348
rect 4396 13336 4402 13388
rect 4724 13385 4752 13416
rect 4798 13404 4804 13456
rect 4856 13404 4862 13456
rect 5626 13444 5632 13456
rect 4908 13416 5632 13444
rect 4908 13385 4936 13416
rect 5626 13404 5632 13416
rect 5684 13444 5690 13456
rect 6546 13444 6552 13456
rect 5684 13416 6552 13444
rect 5684 13404 5690 13416
rect 6546 13404 6552 13416
rect 6604 13404 6610 13456
rect 8386 13404 8392 13456
rect 8444 13404 8450 13456
rect 8496 13444 8524 13472
rect 8757 13447 8815 13453
rect 8757 13444 8769 13447
rect 8496 13416 8769 13444
rect 8757 13413 8769 13416
rect 8803 13413 8815 13447
rect 9582 13444 9588 13456
rect 8757 13407 8815 13413
rect 9140 13416 9588 13444
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13345 4491 13379
rect 4433 13339 4491 13345
rect 4715 13379 4773 13385
rect 4715 13345 4727 13379
rect 4761 13345 4773 13379
rect 4715 13339 4773 13345
rect 4893 13379 4951 13385
rect 4893 13345 4905 13379
rect 4939 13345 4951 13379
rect 4893 13339 4951 13345
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4448 13308 4476 13339
rect 4908 13308 4936 13339
rect 4120 13280 4936 13308
rect 6196 13308 6224 13339
rect 6270 13336 6276 13388
rect 6328 13336 6334 13388
rect 6457 13379 6515 13385
rect 6457 13345 6469 13379
rect 6503 13376 6515 13379
rect 6730 13376 6736 13388
rect 6503 13348 6736 13376
rect 6503 13345 6515 13348
rect 6457 13339 6515 13345
rect 6730 13336 6736 13348
rect 6788 13336 6794 13388
rect 6825 13379 6883 13385
rect 6825 13345 6837 13379
rect 6871 13376 6883 13379
rect 7558 13376 7564 13388
rect 6871 13348 7564 13376
rect 6871 13345 6883 13348
rect 6825 13339 6883 13345
rect 7006 13308 7012 13320
rect 6196 13280 7012 13308
rect 4120 13268 4126 13280
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 4154 13240 4160 13252
rect 3896 13212 4160 13240
rect 4154 13200 4160 13212
rect 4212 13200 4218 13252
rect 4338 13200 4344 13252
rect 4396 13240 4402 13252
rect 4396 13212 5304 13240
rect 4396 13200 4402 13212
rect 2038 13132 2044 13184
rect 2096 13172 2102 13184
rect 2685 13175 2743 13181
rect 2685 13172 2697 13175
rect 2096 13144 2697 13172
rect 2096 13132 2102 13144
rect 2685 13141 2697 13144
rect 2731 13141 2743 13175
rect 2685 13135 2743 13141
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 4982 13172 4988 13184
rect 3927 13144 4988 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 5276 13172 5304 13212
rect 5810 13200 5816 13252
rect 5868 13240 5874 13252
rect 7116 13240 7144 13348
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 8113 13379 8171 13385
rect 8113 13345 8125 13379
rect 8159 13376 8171 13379
rect 8404 13376 8432 13404
rect 8159 13348 8432 13376
rect 8159 13345 8171 13348
rect 8113 13339 8171 13345
rect 8570 13336 8576 13388
rect 8628 13376 8634 13388
rect 8665 13379 8723 13385
rect 8665 13376 8677 13379
rect 8628 13348 8677 13376
rect 8628 13336 8634 13348
rect 8665 13345 8677 13348
rect 8711 13345 8723 13379
rect 8665 13339 8723 13345
rect 8846 13336 8852 13388
rect 8904 13336 8910 13388
rect 9140 13385 9168 13416
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 11624 13444 11652 13475
rect 11882 13472 11888 13524
rect 11940 13472 11946 13524
rect 14274 13512 14280 13524
rect 12084 13484 14280 13512
rect 11974 13444 11980 13456
rect 9784 13416 11980 13444
rect 9125 13379 9183 13385
rect 9125 13345 9137 13379
rect 9171 13345 9183 13379
rect 9125 13339 9183 13345
rect 9214 13336 9220 13388
rect 9272 13336 9278 13388
rect 9398 13336 9404 13388
rect 9456 13336 9462 13388
rect 7926 13268 7932 13320
rect 7984 13308 7990 13320
rect 8205 13311 8263 13317
rect 8205 13308 8217 13311
rect 7984 13280 8217 13308
rect 7984 13268 7990 13280
rect 8205 13277 8217 13280
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 8294 13268 8300 13320
rect 8352 13268 8358 13320
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 8754 13308 8760 13320
rect 8435 13280 8760 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 8754 13268 8760 13280
rect 8812 13308 8818 13320
rect 9784 13308 9812 13416
rect 11974 13404 11980 13416
rect 12032 13404 12038 13456
rect 9858 13336 9864 13388
rect 9916 13376 9922 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9916 13348 10057 13376
rect 9916 13336 9922 13348
rect 10045 13345 10057 13348
rect 10091 13345 10103 13379
rect 10045 13339 10103 13345
rect 8812 13280 9812 13308
rect 10060 13308 10088 13339
rect 10226 13336 10232 13388
rect 10284 13376 10290 13388
rect 11793 13379 11851 13385
rect 11793 13376 11805 13379
rect 10284 13348 11805 13376
rect 10284 13336 10290 13348
rect 11793 13345 11805 13348
rect 11839 13376 11851 13379
rect 12084 13376 12112 13484
rect 12621 13447 12679 13453
rect 12621 13444 12633 13447
rect 12176 13416 12633 13444
rect 12176 13388 12204 13416
rect 12621 13413 12633 13416
rect 12667 13413 12679 13447
rect 12621 13407 12679 13413
rect 11839 13348 12112 13376
rect 11839 13345 11851 13348
rect 11793 13339 11851 13345
rect 12158 13336 12164 13388
rect 12216 13336 12222 13388
rect 12253 13379 12311 13385
rect 12253 13345 12265 13379
rect 12299 13345 12311 13379
rect 12253 13339 12311 13345
rect 12345 13379 12403 13385
rect 12345 13345 12357 13379
rect 12391 13345 12403 13379
rect 12345 13339 12403 13345
rect 12529 13379 12587 13385
rect 12529 13345 12541 13379
rect 12575 13345 12587 13379
rect 12529 13339 12587 13345
rect 12268 13308 12296 13339
rect 10060 13280 12296 13308
rect 8812 13268 8818 13280
rect 5868 13212 7144 13240
rect 9309 13243 9367 13249
rect 5868 13200 5874 13212
rect 9309 13209 9321 13243
rect 9355 13240 9367 13243
rect 9398 13240 9404 13252
rect 9355 13212 9404 13240
rect 9355 13209 9367 13212
rect 9309 13203 9367 13209
rect 9398 13200 9404 13212
rect 9456 13200 9462 13252
rect 12360 13240 12388 13339
rect 12544 13308 12572 13339
rect 13170 13336 13176 13388
rect 13228 13336 13234 13388
rect 14108 13376 14136 13484
rect 14274 13472 14280 13484
rect 14332 13472 14338 13524
rect 14476 13484 15231 13512
rect 14366 13404 14372 13456
rect 14424 13444 14430 13456
rect 14476 13444 14504 13484
rect 15102 13444 15108 13456
rect 14424 13416 14504 13444
rect 14568 13416 15108 13444
rect 14424 13404 14430 13416
rect 14180 13379 14238 13385
rect 14180 13376 14192 13379
rect 14108 13348 14192 13376
rect 14180 13345 14192 13348
rect 14226 13345 14238 13379
rect 14180 13339 14238 13345
rect 14274 13336 14280 13388
rect 14332 13336 14338 13388
rect 14568 13385 14596 13416
rect 15102 13404 15108 13416
rect 15160 13404 15166 13456
rect 15203 13444 15231 13484
rect 16114 13472 16120 13524
rect 16172 13472 16178 13524
rect 16942 13512 16948 13524
rect 16868 13484 16948 13512
rect 16868 13444 16896 13484
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 17037 13515 17095 13521
rect 17037 13481 17049 13515
rect 17083 13512 17095 13515
rect 17678 13512 17684 13524
rect 17083 13484 17684 13512
rect 17083 13481 17095 13484
rect 17037 13475 17095 13481
rect 17678 13472 17684 13484
rect 17736 13472 17742 13524
rect 17770 13472 17776 13524
rect 17828 13472 17834 13524
rect 18141 13515 18199 13521
rect 18141 13481 18153 13515
rect 18187 13512 18199 13515
rect 19613 13515 19671 13521
rect 18187 13484 18368 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 17788 13444 17816 13472
rect 15203 13416 16896 13444
rect 14552 13379 14610 13385
rect 14552 13345 14564 13379
rect 14598 13345 14610 13379
rect 14552 13339 14610 13345
rect 14645 13379 14703 13385
rect 14645 13345 14657 13379
rect 14691 13345 14703 13379
rect 14645 13339 14703 13345
rect 12710 13308 12716 13320
rect 12544 13280 12716 13308
rect 12710 13268 12716 13280
rect 12768 13308 12774 13320
rect 14458 13308 14464 13320
rect 12768 13280 14464 13308
rect 12768 13268 12774 13280
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 14001 13243 14059 13249
rect 14001 13240 14013 13243
rect 9508 13212 11744 13240
rect 12360 13212 14013 13240
rect 6089 13175 6147 13181
rect 6089 13172 6101 13175
rect 5276 13144 6101 13172
rect 6089 13141 6101 13144
rect 6135 13172 6147 13175
rect 6270 13172 6276 13184
rect 6135 13144 6276 13172
rect 6135 13141 6147 13144
rect 6089 13135 6147 13141
rect 6270 13132 6276 13144
rect 6328 13132 6334 13184
rect 7009 13175 7067 13181
rect 7009 13141 7021 13175
rect 7055 13172 7067 13175
rect 8018 13172 8024 13184
rect 7055 13144 8024 13172
rect 7055 13141 7067 13144
rect 7009 13135 7067 13141
rect 8018 13132 8024 13144
rect 8076 13132 8082 13184
rect 8202 13132 8208 13184
rect 8260 13172 8266 13184
rect 9508 13172 9536 13212
rect 8260 13144 9536 13172
rect 8260 13132 8266 13144
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 9861 13175 9919 13181
rect 9861 13172 9873 13175
rect 9824 13144 9873 13172
rect 9824 13132 9830 13144
rect 9861 13141 9873 13144
rect 9907 13141 9919 13175
rect 11716 13172 11744 13212
rect 14001 13209 14013 13212
rect 14047 13209 14059 13243
rect 14001 13203 14059 13209
rect 14660 13240 14688 13339
rect 16390 13336 16396 13388
rect 16448 13336 16454 13388
rect 16485 13379 16543 13385
rect 16485 13345 16497 13379
rect 16531 13345 16543 13379
rect 16485 13339 16543 13345
rect 14734 13268 14740 13320
rect 14792 13268 14798 13320
rect 14918 13268 14924 13320
rect 14976 13308 14982 13320
rect 16500 13308 16528 13339
rect 16574 13336 16580 13388
rect 16632 13336 16638 13388
rect 16758 13336 16764 13388
rect 16816 13336 16822 13388
rect 16868 13385 16896 13416
rect 16960 13416 17816 13444
rect 18340 13444 18368 13484
rect 19613 13481 19625 13515
rect 19659 13512 19671 13515
rect 19886 13512 19892 13524
rect 19659 13484 19892 13512
rect 19659 13481 19671 13484
rect 19613 13475 19671 13481
rect 19886 13472 19892 13484
rect 19944 13472 19950 13524
rect 20533 13515 20591 13521
rect 20533 13481 20545 13515
rect 20579 13512 20591 13515
rect 21082 13512 21088 13524
rect 20579 13484 21088 13512
rect 20579 13481 20591 13484
rect 20533 13475 20591 13481
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 21269 13515 21327 13521
rect 21269 13481 21281 13515
rect 21315 13512 21327 13515
rect 21542 13512 21548 13524
rect 21315 13484 21548 13512
rect 21315 13481 21327 13484
rect 21269 13475 21327 13481
rect 21542 13472 21548 13484
rect 21600 13472 21606 13524
rect 22922 13472 22928 13524
rect 22980 13512 22986 13524
rect 23566 13512 23572 13524
rect 22980 13484 23572 13512
rect 22980 13472 22986 13484
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 24397 13515 24455 13521
rect 24397 13481 24409 13515
rect 24443 13512 24455 13515
rect 24578 13512 24584 13524
rect 24443 13484 24584 13512
rect 24443 13481 24455 13484
rect 24397 13475 24455 13481
rect 24578 13472 24584 13484
rect 24636 13472 24642 13524
rect 25958 13472 25964 13524
rect 26016 13472 26022 13524
rect 18782 13444 18788 13456
rect 18340 13416 18788 13444
rect 16853 13379 16911 13385
rect 16853 13345 16865 13379
rect 16899 13345 16911 13379
rect 16853 13339 16911 13345
rect 16960 13320 16988 13416
rect 17497 13379 17555 13385
rect 17497 13345 17509 13379
rect 17543 13345 17555 13379
rect 17497 13339 17555 13345
rect 16942 13308 16948 13320
rect 14976 13280 16948 13308
rect 14976 13268 14982 13280
rect 16942 13268 16948 13280
rect 17000 13268 17006 13320
rect 16666 13240 16672 13252
rect 14660 13212 16672 13240
rect 14660 13172 14688 13212
rect 16666 13200 16672 13212
rect 16724 13200 16730 13252
rect 16758 13200 16764 13252
rect 16816 13240 16822 13252
rect 17512 13240 17540 13339
rect 17678 13336 17684 13388
rect 17736 13336 17742 13388
rect 17788 13385 17816 13416
rect 18782 13404 18788 13416
rect 18840 13404 18846 13456
rect 20898 13444 20904 13456
rect 20272 13416 20904 13444
rect 18230 13385 18236 13391
rect 17773 13379 17831 13385
rect 17773 13345 17785 13379
rect 17819 13345 17831 13379
rect 17773 13339 17831 13345
rect 17865 13379 17923 13385
rect 17865 13345 17877 13379
rect 17911 13345 17923 13379
rect 17865 13339 17923 13345
rect 18222 13379 18236 13385
rect 18222 13345 18234 13379
rect 18222 13339 18236 13345
rect 18288 13339 18294 13391
rect 18414 13385 18420 13388
rect 18381 13379 18420 13385
rect 18381 13345 18393 13379
rect 18381 13339 18420 13345
rect 17586 13268 17592 13320
rect 17644 13308 17650 13320
rect 17880 13308 17908 13339
rect 18414 13336 18420 13339
rect 18472 13336 18478 13388
rect 18509 13379 18567 13385
rect 18509 13345 18521 13379
rect 18555 13345 18567 13379
rect 18509 13339 18567 13345
rect 17644 13280 17908 13308
rect 17644 13268 17650 13280
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18524 13308 18552 13339
rect 18598 13336 18604 13388
rect 18656 13336 18662 13388
rect 18690 13336 18696 13388
rect 18748 13385 18754 13388
rect 18748 13376 18756 13385
rect 18969 13379 19027 13385
rect 18748 13348 18793 13376
rect 18748 13339 18756 13348
rect 18969 13345 18981 13379
rect 19015 13345 19027 13379
rect 19132 13379 19190 13385
rect 19132 13376 19144 13379
rect 18969 13339 19027 13345
rect 19076 13348 19144 13376
rect 18748 13336 18754 13339
rect 18012 13280 18552 13308
rect 18012 13268 18018 13280
rect 18984 13240 19012 13339
rect 19076 13308 19104 13348
rect 19132 13345 19144 13348
rect 19178 13345 19190 13379
rect 19132 13339 19190 13345
rect 19242 13336 19248 13388
rect 19300 13336 19306 13388
rect 19334 13336 19340 13388
rect 19392 13336 19398 13388
rect 19889 13379 19947 13385
rect 19889 13345 19901 13379
rect 19935 13345 19947 13379
rect 19889 13339 19947 13345
rect 19426 13308 19432 13320
rect 19076 13280 19432 13308
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 19904 13308 19932 13339
rect 20070 13336 20076 13388
rect 20128 13336 20134 13388
rect 20162 13336 20168 13388
rect 20220 13336 20226 13388
rect 20272 13385 20300 13416
rect 20898 13404 20904 13416
rect 20956 13404 20962 13456
rect 22186 13404 22192 13456
rect 22244 13444 22250 13456
rect 24854 13453 24860 13456
rect 22382 13447 22440 13453
rect 22382 13444 22394 13447
rect 22244 13416 22394 13444
rect 22244 13404 22250 13416
rect 22382 13413 22394 13416
rect 22428 13413 22440 13447
rect 24848 13444 24860 13453
rect 22382 13407 22440 13413
rect 22664 13416 24624 13444
rect 24815 13416 24860 13444
rect 20257 13379 20315 13385
rect 20257 13345 20269 13379
rect 20303 13345 20315 13379
rect 20257 13339 20315 13345
rect 20622 13336 20628 13388
rect 20680 13336 20686 13388
rect 22664 13385 22692 13416
rect 22649 13379 22707 13385
rect 22649 13345 22661 13379
rect 22695 13345 22707 13379
rect 22649 13339 22707 13345
rect 22922 13336 22928 13388
rect 22980 13336 22986 13388
rect 23032 13385 23060 13416
rect 23017 13379 23075 13385
rect 23017 13345 23029 13379
rect 23063 13345 23075 13379
rect 23017 13339 23075 13345
rect 23284 13379 23342 13385
rect 23284 13345 23296 13379
rect 23330 13376 23342 13379
rect 23842 13376 23848 13388
rect 23330 13348 23848 13376
rect 23330 13345 23342 13348
rect 23284 13339 23342 13345
rect 23842 13336 23848 13348
rect 23900 13336 23906 13388
rect 24596 13385 24624 13416
rect 24848 13407 24860 13416
rect 24854 13404 24860 13407
rect 24912 13404 24918 13456
rect 24581 13379 24639 13385
rect 24581 13345 24593 13379
rect 24627 13376 24639 13379
rect 24670 13376 24676 13388
rect 24627 13348 24676 13376
rect 24627 13345 24639 13348
rect 24581 13339 24639 13345
rect 24670 13336 24676 13348
rect 24728 13336 24734 13388
rect 27062 13336 27068 13388
rect 27120 13336 27126 13388
rect 21174 13308 21180 13320
rect 19904 13280 21180 13308
rect 19904 13240 19932 13280
rect 21174 13268 21180 13280
rect 21232 13268 21238 13320
rect 16816 13212 17540 13240
rect 16816 13200 16822 13212
rect 11716 13144 14688 13172
rect 9861 13135 9919 13141
rect 15102 13132 15108 13184
rect 15160 13172 15166 13184
rect 15381 13175 15439 13181
rect 15381 13172 15393 13175
rect 15160 13144 15393 13172
rect 15160 13132 15166 13144
rect 15381 13141 15393 13144
rect 15427 13141 15439 13175
rect 17512 13172 17540 13212
rect 17880 13212 19932 13240
rect 20809 13243 20867 13249
rect 17880 13172 17908 13212
rect 20809 13209 20821 13243
rect 20855 13240 20867 13243
rect 20990 13240 20996 13252
rect 20855 13212 20996 13240
rect 20855 13209 20867 13212
rect 20809 13203 20867 13209
rect 20990 13200 20996 13212
rect 21048 13200 21054 13252
rect 17512 13144 17908 13172
rect 15381 13135 15439 13141
rect 18138 13132 18144 13184
rect 18196 13172 18202 13184
rect 18690 13172 18696 13184
rect 18196 13144 18696 13172
rect 18196 13132 18202 13144
rect 18690 13132 18696 13144
rect 18748 13132 18754 13184
rect 18877 13175 18935 13181
rect 18877 13141 18889 13175
rect 18923 13172 18935 13175
rect 19978 13172 19984 13184
rect 18923 13144 19984 13172
rect 18923 13141 18935 13144
rect 18877 13135 18935 13141
rect 19978 13132 19984 13144
rect 20036 13132 20042 13184
rect 22462 13132 22468 13184
rect 22520 13172 22526 13184
rect 22833 13175 22891 13181
rect 22833 13172 22845 13175
rect 22520 13144 22845 13172
rect 22520 13132 22526 13144
rect 22833 13141 22845 13144
rect 22879 13141 22891 13175
rect 22833 13135 22891 13141
rect 24946 13132 24952 13184
rect 25004 13172 25010 13184
rect 26421 13175 26479 13181
rect 26421 13172 26433 13175
rect 25004 13144 26433 13172
rect 25004 13132 25010 13144
rect 26421 13141 26433 13144
rect 26467 13141 26479 13175
rect 26421 13135 26479 13141
rect 552 13082 27416 13104
rect 552 13030 3756 13082
rect 3808 13030 3820 13082
rect 3872 13030 3884 13082
rect 3936 13030 3948 13082
rect 4000 13030 4012 13082
rect 4064 13030 10472 13082
rect 10524 13030 10536 13082
rect 10588 13030 10600 13082
rect 10652 13030 10664 13082
rect 10716 13030 10728 13082
rect 10780 13030 17188 13082
rect 17240 13030 17252 13082
rect 17304 13030 17316 13082
rect 17368 13030 17380 13082
rect 17432 13030 17444 13082
rect 17496 13030 23904 13082
rect 23956 13030 23968 13082
rect 24020 13030 24032 13082
rect 24084 13030 24096 13082
rect 24148 13030 24160 13082
rect 24212 13030 27416 13082
rect 552 13008 27416 13030
rect 4065 12971 4123 12977
rect 4065 12937 4077 12971
rect 4111 12968 4123 12971
rect 4154 12968 4160 12980
rect 4111 12940 4160 12968
rect 4111 12937 4123 12940
rect 4065 12931 4123 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 7466 12928 7472 12980
rect 7524 12968 7530 12980
rect 9398 12968 9404 12980
rect 7524 12940 9404 12968
rect 7524 12928 7530 12940
rect 9398 12928 9404 12940
rect 9456 12968 9462 12980
rect 14182 12968 14188 12980
rect 9456 12940 14188 12968
rect 9456 12928 9462 12940
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 15286 12968 15292 12980
rect 14292 12940 15292 12968
rect 2777 12903 2835 12909
rect 2777 12869 2789 12903
rect 2823 12900 2835 12903
rect 6181 12903 6239 12909
rect 2823 12872 4660 12900
rect 2823 12869 2835 12872
rect 2777 12863 2835 12869
rect 4632 12844 4660 12872
rect 6181 12869 6193 12903
rect 6227 12869 6239 12903
rect 6181 12863 6239 12869
rect 2961 12835 3019 12841
rect 2961 12801 2973 12835
rect 3007 12832 3019 12835
rect 3786 12832 3792 12844
rect 3007 12804 3792 12832
rect 3007 12801 3019 12804
rect 2961 12795 3019 12801
rect 3786 12792 3792 12804
rect 3844 12832 3850 12844
rect 4246 12832 4252 12844
rect 3844 12804 4252 12832
rect 3844 12792 3850 12804
rect 4246 12792 4252 12804
rect 4304 12792 4310 12844
rect 4614 12792 4620 12844
rect 4672 12792 4678 12844
rect 6196 12832 6224 12863
rect 6730 12860 6736 12912
rect 6788 12900 6794 12912
rect 12434 12900 12440 12912
rect 6788 12872 7328 12900
rect 6788 12860 6794 12872
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 6196 12804 6377 12832
rect 6365 12801 6377 12804
rect 6411 12832 6423 12835
rect 7006 12832 7012 12844
rect 6411 12804 7012 12832
rect 6411 12801 6423 12804
rect 6365 12795 6423 12801
rect 7006 12792 7012 12804
rect 7064 12792 7070 12844
rect 7300 12832 7328 12872
rect 9968 12872 12440 12900
rect 9968 12832 9996 12872
rect 12434 12860 12440 12872
rect 12492 12860 12498 12912
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 14292 12900 14320 12940
rect 15286 12928 15292 12940
rect 15344 12968 15350 12980
rect 16298 12968 16304 12980
rect 15344 12940 16304 12968
rect 15344 12928 15350 12940
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 17497 12971 17555 12977
rect 17497 12937 17509 12971
rect 17543 12968 17555 12971
rect 18230 12968 18236 12980
rect 17543 12940 18236 12968
rect 17543 12937 17555 12940
rect 17497 12931 17555 12937
rect 18230 12928 18236 12940
rect 18288 12928 18294 12980
rect 18598 12928 18604 12980
rect 18656 12968 18662 12980
rect 20346 12968 20352 12980
rect 18656 12940 20352 12968
rect 18656 12928 18662 12940
rect 20346 12928 20352 12940
rect 20404 12928 20410 12980
rect 23014 12928 23020 12980
rect 23072 12968 23078 12980
rect 23477 12971 23535 12977
rect 23477 12968 23489 12971
rect 23072 12940 23489 12968
rect 23072 12928 23078 12940
rect 23477 12937 23489 12940
rect 23523 12937 23535 12971
rect 23477 12931 23535 12937
rect 25038 12928 25044 12980
rect 25096 12968 25102 12980
rect 26053 12971 26111 12977
rect 26053 12968 26065 12971
rect 25096 12940 26065 12968
rect 25096 12928 25102 12940
rect 26053 12937 26065 12940
rect 26099 12937 26111 12971
rect 26053 12931 26111 12937
rect 17862 12900 17868 12912
rect 12584 12872 14320 12900
rect 15212 12872 17868 12900
rect 12584 12860 12590 12872
rect 15212 12844 15240 12872
rect 17862 12860 17868 12872
rect 17920 12900 17926 12912
rect 19153 12903 19211 12909
rect 19153 12900 19165 12903
rect 17920 12872 19165 12900
rect 17920 12860 17926 12872
rect 19153 12869 19165 12872
rect 19199 12900 19211 12903
rect 19242 12900 19248 12912
rect 19199 12872 19248 12900
rect 19199 12869 19211 12872
rect 19153 12863 19211 12869
rect 19242 12860 19248 12872
rect 19300 12900 19306 12912
rect 22005 12903 22063 12909
rect 19300 12872 20668 12900
rect 19300 12860 19306 12872
rect 7300 12804 9996 12832
rect 1394 12724 1400 12776
rect 1452 12724 1458 12776
rect 3050 12724 3056 12776
rect 3108 12724 3114 12776
rect 3142 12724 3148 12776
rect 3200 12764 3206 12776
rect 3881 12767 3939 12773
rect 3881 12764 3893 12767
rect 3200 12736 3893 12764
rect 3200 12724 3206 12736
rect 3881 12733 3893 12736
rect 3927 12733 3939 12767
rect 3881 12727 3939 12733
rect 4798 12724 4804 12776
rect 4856 12724 4862 12776
rect 6546 12724 6552 12776
rect 6604 12724 6610 12776
rect 7101 12767 7159 12773
rect 7101 12733 7113 12767
rect 7147 12764 7159 12767
rect 7466 12764 7472 12776
rect 7147 12736 7472 12764
rect 7147 12733 7159 12736
rect 7101 12727 7159 12733
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 7558 12724 7564 12776
rect 7616 12724 7622 12776
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12764 7987 12767
rect 8202 12764 8208 12776
rect 7975 12736 8208 12764
rect 7975 12733 7987 12736
rect 7929 12727 7987 12733
rect 8202 12724 8208 12736
rect 8260 12764 8266 12776
rect 8496 12773 8524 12804
rect 8389 12767 8447 12773
rect 8389 12764 8401 12767
rect 8260 12736 8401 12764
rect 8260 12724 8266 12736
rect 8389 12733 8401 12736
rect 8435 12733 8447 12767
rect 8389 12727 8447 12733
rect 8481 12767 8539 12773
rect 8481 12733 8493 12767
rect 8527 12733 8539 12767
rect 8481 12727 8539 12733
rect 8662 12724 8668 12776
rect 8720 12724 8726 12776
rect 8754 12724 8760 12776
rect 8812 12724 8818 12776
rect 9490 12724 9496 12776
rect 9548 12724 9554 12776
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 9858 12764 9864 12776
rect 9723 12736 9864 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 9968 12773 9996 12804
rect 11164 12804 11744 12832
rect 10134 12773 10140 12776
rect 9953 12767 10011 12773
rect 9953 12733 9965 12767
rect 9999 12733 10011 12767
rect 9953 12727 10011 12733
rect 10101 12767 10140 12773
rect 10101 12733 10113 12767
rect 10101 12727 10140 12733
rect 10134 12724 10140 12727
rect 10192 12724 10198 12776
rect 10226 12724 10232 12776
rect 10284 12724 10290 12776
rect 10318 12724 10324 12776
rect 10376 12724 10382 12776
rect 10459 12767 10517 12773
rect 10459 12733 10471 12767
rect 10505 12764 10517 12767
rect 10505 12736 10640 12764
rect 10505 12733 10517 12736
rect 10459 12727 10517 12733
rect 1664 12699 1722 12705
rect 1664 12665 1676 12699
rect 1710 12696 1722 12699
rect 4062 12696 4068 12708
rect 1710 12668 4068 12696
rect 1710 12665 1722 12668
rect 1664 12659 1722 12665
rect 4062 12656 4068 12668
rect 4120 12656 4126 12708
rect 4890 12656 4896 12708
rect 4948 12696 4954 12708
rect 5046 12699 5104 12705
rect 5046 12696 5058 12699
rect 4948 12668 5058 12696
rect 4948 12656 4954 12668
rect 5046 12665 5058 12668
rect 5092 12665 5104 12699
rect 5046 12659 5104 12665
rect 6733 12699 6791 12705
rect 6733 12665 6745 12699
rect 6779 12696 6791 12699
rect 6917 12699 6975 12705
rect 6917 12696 6929 12699
rect 6779 12668 6929 12696
rect 6779 12665 6791 12668
rect 6733 12659 6791 12665
rect 6917 12665 6929 12668
rect 6963 12665 6975 12699
rect 9214 12696 9220 12708
rect 6917 12659 6975 12665
rect 7024 12668 9220 12696
rect 3326 12588 3332 12640
rect 3384 12588 3390 12640
rect 3418 12588 3424 12640
rect 3476 12628 3482 12640
rect 7024 12628 7052 12668
rect 3476 12600 7052 12628
rect 7285 12631 7343 12637
rect 3476 12588 3482 12600
rect 7285 12597 7297 12631
rect 7331 12628 7343 12631
rect 7466 12628 7472 12640
rect 7331 12600 7472 12628
rect 7331 12597 7343 12600
rect 7285 12591 7343 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 7760 12637 7788 12668
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 10612 12696 10640 12736
rect 10686 12724 10692 12776
rect 10744 12724 10750 12776
rect 10962 12696 10968 12708
rect 10612 12668 10968 12696
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 7745 12631 7803 12637
rect 7745 12597 7757 12631
rect 7791 12628 7803 12631
rect 7926 12628 7932 12640
rect 7791 12600 7932 12628
rect 7791 12597 7803 12600
rect 7745 12591 7803 12597
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 8113 12631 8171 12637
rect 8113 12597 8125 12631
rect 8159 12628 8171 12631
rect 8846 12628 8852 12640
rect 8159 12600 8852 12628
rect 8159 12597 8171 12600
rect 8113 12591 8171 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 8938 12588 8944 12640
rect 8996 12588 9002 12640
rect 9030 12588 9036 12640
rect 9088 12628 9094 12640
rect 9309 12631 9367 12637
rect 9309 12628 9321 12631
rect 9088 12600 9321 12628
rect 9088 12588 9094 12600
rect 9309 12597 9321 12600
rect 9355 12597 9367 12631
rect 9309 12591 9367 12597
rect 10597 12631 10655 12637
rect 10597 12597 10609 12631
rect 10643 12628 10655 12631
rect 11164 12628 11192 12804
rect 11425 12767 11483 12773
rect 11425 12733 11437 12767
rect 11471 12733 11483 12767
rect 11425 12727 11483 12733
rect 11440 12696 11468 12727
rect 11606 12724 11612 12776
rect 11664 12724 11670 12776
rect 11716 12773 11744 12804
rect 11808 12804 13400 12832
rect 11808 12776 11836 12804
rect 13372 12776 13400 12804
rect 15194 12792 15200 12844
rect 15252 12792 15258 12844
rect 16577 12835 16635 12841
rect 16577 12832 16589 12835
rect 15396 12804 16589 12832
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12733 11759 12767
rect 11701 12727 11759 12733
rect 11790 12724 11796 12776
rect 11848 12724 11854 12776
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12892 12767 12950 12773
rect 12892 12764 12904 12767
rect 12032 12736 12904 12764
rect 12032 12724 12038 12736
rect 12892 12733 12904 12736
rect 12938 12733 12950 12767
rect 13262 12764 13268 12776
rect 13223 12736 13268 12764
rect 12892 12727 12950 12733
rect 12526 12696 12532 12708
rect 11440 12668 12532 12696
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 10643 12600 11192 12628
rect 10643 12597 10655 12600
rect 10597 12591 10655 12597
rect 11330 12588 11336 12640
rect 11388 12588 11394 12640
rect 12066 12588 12072 12640
rect 12124 12588 12130 12640
rect 12250 12588 12256 12640
rect 12308 12628 12314 12640
rect 12713 12631 12771 12637
rect 12713 12628 12725 12631
rect 12308 12600 12725 12628
rect 12308 12588 12314 12600
rect 12713 12597 12725 12600
rect 12759 12597 12771 12631
rect 12912 12628 12940 12727
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 13354 12724 13360 12776
rect 13412 12724 13418 12776
rect 14941 12767 14999 12773
rect 14941 12733 14953 12767
rect 14987 12764 14999 12767
rect 15102 12764 15108 12776
rect 14987 12736 15108 12764
rect 14987 12733 14999 12736
rect 14941 12727 14999 12733
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 15286 12724 15292 12776
rect 15344 12724 15350 12776
rect 12986 12656 12992 12708
rect 13044 12656 13050 12708
rect 13081 12699 13139 12705
rect 13081 12665 13093 12699
rect 13127 12696 13139 12699
rect 13170 12696 13176 12708
rect 13127 12668 13176 12696
rect 13127 12665 13139 12668
rect 13081 12659 13139 12665
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 14274 12696 14280 12708
rect 13832 12668 14280 12696
rect 13446 12628 13452 12640
rect 12912 12600 13452 12628
rect 12713 12591 12771 12597
rect 13446 12588 13452 12600
rect 13504 12588 13510 12640
rect 13832 12637 13860 12668
rect 14274 12656 14280 12668
rect 14332 12696 14338 12708
rect 15396 12696 15424 12804
rect 16577 12801 16589 12804
rect 16623 12801 16635 12835
rect 16577 12795 16635 12801
rect 16666 12792 16672 12844
rect 16724 12832 16730 12844
rect 20640 12841 20668 12872
rect 22005 12869 22017 12903
rect 22051 12900 22063 12903
rect 24489 12903 24547 12909
rect 22051 12872 22876 12900
rect 22051 12869 22063 12872
rect 22005 12863 22063 12869
rect 22848 12841 22876 12872
rect 24489 12869 24501 12903
rect 24535 12869 24547 12903
rect 24489 12863 24547 12869
rect 20625 12835 20683 12841
rect 16724 12804 17356 12832
rect 16724 12792 16730 12804
rect 15470 12724 15476 12776
rect 15528 12724 15534 12776
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12733 15623 12767
rect 15565 12727 15623 12733
rect 15657 12767 15715 12773
rect 15657 12733 15669 12767
rect 15703 12764 15715 12767
rect 16482 12764 16488 12776
rect 15703 12736 16488 12764
rect 15703 12733 15715 12736
rect 15657 12727 15715 12733
rect 14332 12668 15424 12696
rect 15580 12696 15608 12727
rect 16482 12724 16488 12736
rect 16540 12724 16546 12776
rect 16942 12724 16948 12776
rect 17000 12724 17006 12776
rect 17328 12773 17356 12804
rect 20625 12801 20637 12835
rect 20671 12801 20683 12835
rect 22833 12835 22891 12841
rect 20625 12795 20683 12801
rect 21652 12804 22416 12832
rect 17313 12767 17371 12773
rect 17313 12733 17325 12767
rect 17359 12733 17371 12767
rect 17313 12727 17371 12733
rect 18322 12724 18328 12776
rect 18380 12724 18386 12776
rect 21652 12764 21680 12804
rect 20272 12736 21680 12764
rect 20272 12708 20300 12736
rect 22094 12724 22100 12776
rect 22152 12724 22158 12776
rect 22278 12724 22284 12776
rect 22336 12724 22342 12776
rect 22388 12773 22416 12804
rect 22833 12801 22845 12835
rect 22879 12801 22891 12835
rect 22833 12795 22891 12801
rect 23658 12792 23664 12844
rect 23716 12832 23722 12844
rect 24504 12832 24532 12863
rect 24854 12860 24860 12912
rect 24912 12900 24918 12912
rect 24912 12872 25636 12900
rect 24912 12860 24918 12872
rect 23716 12804 24164 12832
rect 24504 12804 25544 12832
rect 23716 12792 23722 12804
rect 22373 12767 22431 12773
rect 22373 12733 22385 12767
rect 22419 12733 22431 12767
rect 22373 12727 22431 12733
rect 22465 12767 22523 12773
rect 22465 12733 22477 12767
rect 22511 12764 22523 12767
rect 23014 12764 23020 12776
rect 22511 12736 23020 12764
rect 22511 12733 22523 12736
rect 22465 12727 22523 12733
rect 23014 12724 23020 12736
rect 23072 12724 23078 12776
rect 23382 12724 23388 12776
rect 23440 12764 23446 12776
rect 24136 12773 24164 12804
rect 23845 12767 23903 12773
rect 23845 12764 23857 12767
rect 23440 12736 23857 12764
rect 23440 12724 23446 12736
rect 23845 12733 23857 12736
rect 23891 12733 23903 12767
rect 23845 12727 23903 12733
rect 23938 12767 23996 12773
rect 23938 12733 23950 12767
rect 23984 12733 23996 12767
rect 23938 12727 23996 12733
rect 24121 12767 24179 12773
rect 24121 12733 24133 12767
rect 24167 12733 24179 12767
rect 24121 12727 24179 12733
rect 15746 12696 15752 12708
rect 15580 12668 15752 12696
rect 14332 12656 14338 12668
rect 15746 12656 15752 12668
rect 15804 12656 15810 12708
rect 15933 12699 15991 12705
rect 15933 12665 15945 12699
rect 15979 12696 15991 12699
rect 16666 12696 16672 12708
rect 15979 12668 16672 12696
rect 15979 12665 15991 12668
rect 15933 12659 15991 12665
rect 16666 12656 16672 12668
rect 16724 12656 16730 12708
rect 18230 12696 18236 12708
rect 17144 12668 18236 12696
rect 13817 12631 13875 12637
rect 13817 12597 13829 12631
rect 13863 12597 13875 12631
rect 13817 12591 13875 12597
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 17144 12637 17172 12668
rect 18230 12656 18236 12668
rect 18288 12696 18294 12708
rect 20254 12696 20260 12708
rect 18288 12668 20260 12696
rect 18288 12656 18294 12668
rect 20254 12656 20260 12668
rect 20312 12656 20318 12708
rect 20438 12656 20444 12708
rect 20496 12656 20502 12708
rect 20892 12699 20950 12705
rect 20892 12665 20904 12699
rect 20938 12696 20950 12699
rect 22741 12699 22799 12705
rect 22741 12696 22753 12699
rect 20938 12668 22753 12696
rect 20938 12665 20950 12668
rect 20892 12659 20950 12665
rect 22741 12665 22753 12668
rect 22787 12665 22799 12699
rect 23952 12696 23980 12727
rect 24302 12724 24308 12776
rect 24360 12773 24366 12776
rect 24360 12764 24368 12773
rect 24360 12736 24405 12764
rect 24360 12727 24368 12736
rect 24360 12724 24366 12727
rect 24486 12724 24492 12776
rect 24544 12764 24550 12776
rect 24581 12767 24639 12773
rect 24581 12764 24593 12767
rect 24544 12736 24593 12764
rect 24544 12724 24550 12736
rect 24581 12733 24593 12736
rect 24627 12733 24639 12767
rect 24581 12727 24639 12733
rect 24670 12724 24676 12776
rect 24728 12764 24734 12776
rect 24765 12767 24823 12773
rect 24765 12764 24777 12767
rect 24728 12736 24777 12764
rect 24728 12724 24734 12736
rect 24765 12733 24777 12736
rect 24811 12733 24823 12767
rect 24765 12727 24823 12733
rect 24854 12724 24860 12776
rect 24912 12724 24918 12776
rect 24946 12724 24952 12776
rect 25004 12724 25010 12776
rect 25314 12724 25320 12776
rect 25372 12724 25378 12776
rect 25516 12773 25544 12804
rect 25608 12773 25636 12872
rect 25866 12860 25872 12912
rect 25924 12900 25930 12912
rect 25961 12903 26019 12909
rect 25961 12900 25973 12903
rect 25924 12872 25973 12900
rect 25924 12860 25930 12872
rect 25961 12869 25973 12872
rect 26007 12869 26019 12903
rect 25961 12863 26019 12869
rect 25700 12804 26372 12832
rect 25700 12776 25728 12804
rect 25501 12767 25559 12773
rect 25501 12733 25513 12767
rect 25547 12733 25559 12767
rect 25501 12727 25559 12733
rect 25593 12767 25651 12773
rect 25593 12733 25605 12767
rect 25639 12733 25651 12767
rect 25593 12727 25651 12733
rect 25682 12724 25688 12776
rect 25740 12724 25746 12776
rect 25774 12724 25780 12776
rect 25832 12764 25838 12776
rect 26191 12767 26249 12773
rect 26191 12764 26203 12767
rect 25832 12736 26203 12764
rect 25832 12724 25838 12736
rect 26191 12733 26203 12736
rect 26237 12733 26249 12767
rect 26344 12764 26372 12804
rect 26418 12792 26424 12844
rect 26476 12832 26482 12844
rect 26476 12804 26740 12832
rect 26476 12792 26482 12804
rect 26712 12773 26740 12804
rect 26549 12767 26607 12773
rect 26549 12764 26561 12767
rect 26344 12736 26561 12764
rect 26191 12727 26249 12733
rect 26549 12733 26561 12736
rect 26595 12733 26607 12767
rect 26549 12727 26607 12733
rect 26697 12767 26755 12773
rect 26697 12733 26709 12767
rect 26743 12733 26755 12767
rect 26697 12727 26755 12733
rect 22741 12659 22799 12665
rect 23032 12668 23980 12696
rect 24213 12699 24271 12705
rect 16025 12631 16083 12637
rect 16025 12628 16037 12631
rect 14884 12600 16037 12628
rect 14884 12588 14890 12600
rect 16025 12597 16037 12600
rect 16071 12597 16083 12631
rect 16025 12591 16083 12597
rect 17129 12631 17187 12637
rect 17129 12597 17141 12631
rect 17175 12597 17187 12631
rect 17129 12591 17187 12597
rect 17678 12588 17684 12640
rect 17736 12588 17742 12640
rect 21174 12588 21180 12640
rect 21232 12628 21238 12640
rect 21818 12628 21824 12640
rect 21232 12600 21824 12628
rect 21232 12588 21238 12600
rect 21818 12588 21824 12600
rect 21876 12588 21882 12640
rect 21910 12588 21916 12640
rect 21968 12628 21974 12640
rect 23032 12628 23060 12668
rect 24213 12665 24225 12699
rect 24259 12696 24271 12699
rect 24259 12668 24440 12696
rect 24259 12665 24271 12668
rect 24213 12659 24271 12665
rect 24412 12640 24440 12668
rect 26326 12656 26332 12708
rect 26384 12656 26390 12708
rect 26418 12656 26424 12708
rect 26476 12656 26482 12708
rect 21968 12600 23060 12628
rect 21968 12588 21974 12600
rect 24394 12588 24400 12640
rect 24452 12588 24458 12640
rect 25222 12588 25228 12640
rect 25280 12588 25286 12640
rect 552 12538 27576 12560
rect 552 12486 7114 12538
rect 7166 12486 7178 12538
rect 7230 12486 7242 12538
rect 7294 12486 7306 12538
rect 7358 12486 7370 12538
rect 7422 12486 13830 12538
rect 13882 12486 13894 12538
rect 13946 12486 13958 12538
rect 14010 12486 14022 12538
rect 14074 12486 14086 12538
rect 14138 12486 20546 12538
rect 20598 12486 20610 12538
rect 20662 12486 20674 12538
rect 20726 12486 20738 12538
rect 20790 12486 20802 12538
rect 20854 12486 27262 12538
rect 27314 12486 27326 12538
rect 27378 12486 27390 12538
rect 27442 12486 27454 12538
rect 27506 12486 27518 12538
rect 27570 12486 27576 12538
rect 552 12464 27576 12486
rect 2682 12384 2688 12436
rect 2740 12424 2746 12436
rect 4798 12424 4804 12436
rect 2740 12396 4804 12424
rect 2740 12384 2746 12396
rect 4798 12384 4804 12396
rect 4856 12424 4862 12436
rect 6914 12424 6920 12436
rect 4856 12396 6920 12424
rect 4856 12384 4862 12396
rect 6914 12384 6920 12396
rect 6972 12424 6978 12436
rect 7742 12424 7748 12436
rect 6972 12396 7748 12424
rect 6972 12384 6978 12396
rect 7742 12384 7748 12396
rect 7800 12424 7806 12436
rect 7929 12427 7987 12433
rect 7929 12424 7941 12427
rect 7800 12396 7941 12424
rect 7800 12384 7806 12396
rect 7929 12393 7941 12396
rect 7975 12393 7987 12427
rect 7929 12387 7987 12393
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 10870 12424 10876 12436
rect 8076 12396 10876 12424
rect 8076 12384 8082 12396
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 14645 12427 14703 12433
rect 14645 12393 14657 12427
rect 14691 12424 14703 12427
rect 14734 12424 14740 12436
rect 14691 12396 14740 12424
rect 14691 12393 14703 12396
rect 14645 12387 14703 12393
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 14918 12384 14924 12436
rect 14976 12384 14982 12436
rect 16482 12384 16488 12436
rect 16540 12424 16546 12436
rect 16853 12427 16911 12433
rect 16853 12424 16865 12427
rect 16540 12396 16865 12424
rect 16540 12384 16546 12396
rect 16853 12393 16865 12396
rect 16899 12393 16911 12427
rect 16853 12387 16911 12393
rect 18322 12384 18328 12436
rect 18380 12424 18386 12436
rect 18969 12427 19027 12433
rect 18969 12424 18981 12427
rect 18380 12396 18981 12424
rect 18380 12384 18386 12396
rect 18969 12393 18981 12396
rect 19015 12393 19027 12427
rect 18969 12387 19027 12393
rect 26237 12427 26295 12433
rect 26237 12393 26249 12427
rect 26283 12424 26295 12427
rect 27062 12424 27068 12436
rect 26283 12396 27068 12424
rect 26283 12393 26295 12396
rect 26237 12387 26295 12393
rect 27062 12384 27068 12396
rect 27120 12384 27126 12436
rect 1394 12316 1400 12368
rect 1452 12356 1458 12368
rect 2700 12356 2728 12384
rect 1452 12328 2728 12356
rect 1452 12316 1458 12328
rect 1780 12297 1808 12328
rect 3602 12316 3608 12368
rect 3660 12316 3666 12368
rect 4154 12316 4160 12368
rect 4212 12356 4218 12368
rect 4249 12359 4307 12365
rect 4249 12356 4261 12359
rect 4212 12328 4261 12356
rect 4212 12316 4218 12328
rect 4249 12325 4261 12328
rect 4295 12325 4307 12359
rect 4249 12319 4307 12325
rect 4338 12316 4344 12368
rect 4396 12356 4402 12368
rect 4433 12359 4491 12365
rect 4433 12356 4445 12359
rect 4396 12328 4445 12356
rect 4396 12316 4402 12328
rect 4433 12325 4445 12328
rect 4479 12325 4491 12359
rect 4433 12319 4491 12325
rect 5166 12316 5172 12368
rect 5224 12356 5230 12368
rect 5997 12359 6055 12365
rect 5997 12356 6009 12359
rect 5224 12328 6009 12356
rect 5224 12316 5230 12328
rect 5997 12325 6009 12328
rect 6043 12325 6055 12359
rect 5997 12319 6055 12325
rect 8846 12316 8852 12368
rect 8904 12356 8910 12368
rect 10045 12359 10103 12365
rect 8904 12328 9996 12356
rect 8904 12316 8910 12328
rect 2038 12297 2044 12300
rect 1765 12291 1823 12297
rect 1765 12257 1777 12291
rect 1811 12257 1823 12291
rect 2032 12288 2044 12297
rect 1999 12260 2044 12288
rect 1765 12251 1823 12257
rect 2032 12251 2044 12260
rect 2038 12248 2044 12251
rect 2096 12248 2102 12300
rect 3326 12248 3332 12300
rect 3384 12288 3390 12300
rect 3513 12291 3571 12297
rect 3513 12288 3525 12291
rect 3384 12260 3525 12288
rect 3384 12248 3390 12260
rect 3513 12257 3525 12260
rect 3559 12257 3571 12291
rect 3620 12288 3648 12316
rect 3697 12291 3755 12297
rect 3697 12288 3709 12291
rect 3620 12260 3709 12288
rect 3513 12251 3571 12257
rect 3697 12257 3709 12260
rect 3743 12257 3755 12291
rect 3697 12251 3755 12257
rect 3881 12291 3939 12297
rect 3881 12257 3893 12291
rect 3927 12257 3939 12291
rect 3881 12251 3939 12257
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 3418 12180 3424 12232
rect 3476 12180 3482 12232
rect 3605 12223 3663 12229
rect 3605 12189 3617 12223
rect 3651 12220 3663 12223
rect 3786 12220 3792 12232
rect 3651 12192 3792 12220
rect 3651 12189 3663 12192
rect 3605 12183 3663 12189
rect 3786 12180 3792 12192
rect 3844 12180 3850 12232
rect 3142 12044 3148 12096
rect 3200 12044 3206 12096
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 3896 12084 3924 12251
rect 4522 12248 4528 12300
rect 4580 12248 4586 12300
rect 4798 12248 4804 12300
rect 4856 12288 4862 12300
rect 5077 12291 5135 12297
rect 5077 12288 5089 12291
rect 4856 12260 5089 12288
rect 4856 12248 4862 12260
rect 5077 12257 5089 12260
rect 5123 12288 5135 12291
rect 5353 12291 5411 12297
rect 5353 12288 5365 12291
rect 5123 12260 5365 12288
rect 5123 12257 5135 12260
rect 5077 12251 5135 12257
rect 5353 12257 5365 12260
rect 5399 12257 5411 12291
rect 5353 12251 5411 12257
rect 6638 12248 6644 12300
rect 6696 12248 6702 12300
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 8665 12291 8723 12297
rect 8665 12288 8677 12291
rect 8628 12260 8677 12288
rect 8628 12248 8634 12260
rect 8665 12257 8677 12260
rect 8711 12257 8723 12291
rect 8665 12251 8723 12257
rect 8938 12248 8944 12300
rect 8996 12248 9002 12300
rect 9030 12248 9036 12300
rect 9088 12248 9094 12300
rect 9214 12248 9220 12300
rect 9272 12248 9278 12300
rect 9490 12248 9496 12300
rect 9548 12288 9554 12300
rect 9585 12291 9643 12297
rect 9585 12288 9597 12291
rect 9548 12260 9597 12288
rect 9548 12248 9554 12260
rect 9585 12257 9597 12260
rect 9631 12257 9643 12291
rect 9585 12251 9643 12257
rect 9674 12248 9680 12300
rect 9732 12248 9738 12300
rect 9858 12248 9864 12300
rect 9916 12248 9922 12300
rect 9968 12288 9996 12328
rect 10045 12325 10057 12359
rect 10091 12356 10103 12359
rect 11606 12356 11612 12368
rect 10091 12328 11612 12356
rect 10091 12325 10103 12328
rect 10045 12319 10103 12325
rect 11606 12316 11612 12328
rect 11664 12316 11670 12368
rect 12713 12359 12771 12365
rect 12713 12325 12725 12359
rect 12759 12356 12771 12359
rect 12802 12356 12808 12368
rect 12759 12328 12808 12356
rect 12759 12325 12771 12328
rect 12713 12319 12771 12325
rect 12802 12316 12808 12328
rect 12860 12316 12866 12368
rect 14182 12316 14188 12368
rect 14240 12356 14246 12368
rect 14936 12356 14964 12384
rect 16758 12356 16764 12368
rect 14240 12328 14964 12356
rect 15304 12328 16764 12356
rect 14240 12316 14246 12328
rect 9968 12260 10916 12288
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 4203 12192 5396 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 5368 12164 5396 12192
rect 5442 12180 5448 12232
rect 5500 12220 5506 12232
rect 5905 12223 5963 12229
rect 5905 12220 5917 12223
rect 5500 12192 5917 12220
rect 5500 12180 5506 12192
rect 5905 12189 5917 12192
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 6089 12223 6147 12229
rect 6089 12189 6101 12223
rect 6135 12220 6147 12223
rect 8849 12223 8907 12229
rect 6135 12192 8800 12220
rect 6135 12189 6147 12192
rect 6089 12183 6147 12189
rect 4062 12112 4068 12164
rect 4120 12112 4126 12164
rect 4430 12112 4436 12164
rect 4488 12152 4494 12164
rect 4798 12152 4804 12164
rect 4488 12124 4804 12152
rect 4488 12112 4494 12124
rect 4798 12112 4804 12124
rect 4856 12112 4862 12164
rect 5350 12112 5356 12164
rect 5408 12112 5414 12164
rect 8772 12152 8800 12192
rect 8849 12189 8861 12223
rect 8895 12220 8907 12223
rect 9692 12220 9720 12248
rect 8895 12192 9720 12220
rect 8895 12189 8907 12192
rect 8849 12183 8907 12189
rect 9876 12152 9904 12248
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 10008 12192 10149 12220
rect 10008 12180 10014 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10686 12220 10692 12232
rect 10284 12192 10692 12220
rect 10284 12180 10290 12192
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 10888 12220 10916 12260
rect 10962 12248 10968 12300
rect 11020 12248 11026 12300
rect 11054 12248 11060 12300
rect 11112 12288 11118 12300
rect 11112 12260 14504 12288
rect 11112 12248 11118 12260
rect 11238 12220 11244 12232
rect 10888 12192 11244 12220
rect 11238 12180 11244 12192
rect 11296 12220 11302 12232
rect 11790 12220 11796 12232
rect 11296 12192 11796 12220
rect 11296 12180 11302 12192
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 13078 12180 13084 12232
rect 13136 12220 13142 12232
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 13136 12192 13185 12220
rect 13136 12180 13142 12192
rect 13173 12189 13185 12192
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 12710 12152 12716 12164
rect 8772 12124 9536 12152
rect 9876 12124 12716 12152
rect 3660 12056 3924 12084
rect 3973 12087 4031 12093
rect 3660 12044 3666 12056
rect 3973 12053 3985 12087
rect 4019 12084 4031 12087
rect 4249 12087 4307 12093
rect 4249 12084 4261 12087
rect 4019 12056 4261 12084
rect 4019 12053 4031 12056
rect 3973 12047 4031 12053
rect 4249 12053 4261 12056
rect 4295 12053 4307 12087
rect 4249 12047 4307 12053
rect 5537 12087 5595 12093
rect 5537 12053 5549 12087
rect 5583 12084 5595 12087
rect 5626 12084 5632 12096
rect 5583 12056 5632 12084
rect 5583 12053 5595 12056
rect 5537 12047 5595 12053
rect 5626 12044 5632 12056
rect 5684 12044 5690 12096
rect 6457 12087 6515 12093
rect 6457 12053 6469 12087
rect 6503 12084 6515 12087
rect 6638 12084 6644 12096
rect 6503 12056 6644 12084
rect 6503 12053 6515 12056
rect 6457 12047 6515 12053
rect 6638 12044 6644 12056
rect 6696 12044 6702 12096
rect 8478 12044 8484 12096
rect 8536 12044 8542 12096
rect 8570 12044 8576 12096
rect 8628 12084 8634 12096
rect 9030 12084 9036 12096
rect 8628 12056 9036 12084
rect 8628 12044 8634 12056
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 9398 12044 9404 12096
rect 9456 12044 9462 12096
rect 9508 12084 9536 12124
rect 12710 12112 12716 12124
rect 12768 12112 12774 12164
rect 12802 12112 12808 12164
rect 12860 12152 12866 12164
rect 13909 12155 13967 12161
rect 13909 12152 13921 12155
rect 12860 12124 13921 12152
rect 12860 12112 12866 12124
rect 13909 12121 13921 12124
rect 13955 12121 13967 12155
rect 13909 12115 13967 12121
rect 13722 12084 13728 12096
rect 9508 12056 13728 12084
rect 13722 12044 13728 12056
rect 13780 12044 13786 12096
rect 13814 12044 13820 12096
rect 13872 12044 13878 12096
rect 14476 12084 14504 12260
rect 14550 12180 14556 12232
rect 14608 12180 14614 12232
rect 14753 12220 14781 12328
rect 14826 12248 14832 12300
rect 14884 12297 14890 12300
rect 14884 12291 14933 12297
rect 14884 12257 14887 12291
rect 14921 12257 14933 12291
rect 14884 12251 14933 12257
rect 15013 12291 15071 12297
rect 15013 12257 15025 12291
rect 15059 12257 15071 12291
rect 15013 12251 15071 12257
rect 14884 12248 14890 12251
rect 15028 12220 15056 12251
rect 15102 12248 15108 12300
rect 15160 12248 15166 12300
rect 15304 12297 15332 12328
rect 16758 12316 16764 12328
rect 16816 12316 16822 12368
rect 16868 12328 18368 12356
rect 15289 12291 15347 12297
rect 15289 12257 15301 12291
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 16666 12248 16672 12300
rect 16724 12248 16730 12300
rect 14753 12192 15056 12220
rect 16298 12180 16304 12232
rect 16356 12220 16362 12232
rect 16868 12220 16896 12328
rect 17586 12248 17592 12300
rect 17644 12248 17650 12300
rect 17682 12291 17740 12297
rect 17682 12257 17694 12291
rect 17728 12257 17740 12291
rect 17682 12251 17740 12257
rect 16356 12192 16896 12220
rect 16356 12180 16362 12192
rect 16942 12180 16948 12232
rect 17000 12220 17006 12232
rect 17405 12223 17463 12229
rect 17405 12220 17417 12223
rect 17000 12192 17417 12220
rect 17000 12180 17006 12192
rect 17405 12189 17417 12192
rect 17451 12220 17463 12223
rect 17696 12220 17724 12251
rect 17862 12248 17868 12300
rect 17920 12248 17926 12300
rect 17954 12248 17960 12300
rect 18012 12248 18018 12300
rect 18138 12297 18144 12300
rect 18095 12291 18144 12297
rect 18095 12257 18107 12291
rect 18141 12257 18144 12291
rect 18095 12251 18144 12257
rect 18138 12248 18144 12251
rect 18196 12248 18202 12300
rect 18340 12297 18368 12328
rect 18414 12316 18420 12368
rect 18472 12356 18478 12368
rect 18472 12328 18736 12356
rect 18472 12316 18478 12328
rect 18325 12291 18383 12297
rect 18325 12257 18337 12291
rect 18371 12257 18383 12291
rect 18325 12251 18383 12257
rect 18509 12291 18567 12297
rect 18509 12257 18521 12291
rect 18555 12257 18567 12291
rect 18509 12251 18567 12257
rect 18524 12220 18552 12251
rect 18598 12248 18604 12300
rect 18656 12248 18662 12300
rect 18708 12297 18736 12328
rect 19794 12316 19800 12368
rect 19852 12356 19858 12368
rect 21269 12359 21327 12365
rect 21269 12356 21281 12359
rect 19852 12328 21281 12356
rect 19852 12316 19858 12328
rect 21269 12325 21281 12328
rect 21315 12325 21327 12359
rect 21269 12319 21327 12325
rect 25124 12359 25182 12365
rect 25124 12325 25136 12359
rect 25170 12356 25182 12359
rect 25222 12356 25228 12368
rect 25170 12328 25228 12356
rect 25170 12325 25182 12328
rect 25124 12319 25182 12325
rect 25222 12316 25228 12328
rect 25280 12316 25286 12368
rect 19518 12297 19524 12300
rect 18693 12291 18751 12297
rect 18693 12257 18705 12291
rect 18739 12257 18751 12291
rect 18693 12251 18751 12257
rect 19512 12251 19524 12297
rect 19518 12248 19524 12251
rect 19576 12248 19582 12300
rect 20438 12248 20444 12300
rect 20496 12288 20502 12300
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 20496 12260 22017 12288
rect 20496 12248 20502 12260
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 26234 12248 26240 12300
rect 26292 12288 26298 12300
rect 26878 12288 26884 12300
rect 26292 12260 26884 12288
rect 26292 12248 26298 12260
rect 26878 12248 26884 12260
rect 26936 12288 26942 12300
rect 27065 12291 27123 12297
rect 27065 12288 27077 12291
rect 26936 12260 27077 12288
rect 26936 12248 26942 12260
rect 27065 12257 27077 12260
rect 27111 12257 27123 12291
rect 27065 12251 27123 12257
rect 17451 12192 17724 12220
rect 18248 12192 18552 12220
rect 17451 12189 17463 12192
rect 17405 12183 17463 12189
rect 18248 12161 18276 12192
rect 19242 12180 19248 12232
rect 19300 12180 19306 12232
rect 21821 12223 21879 12229
rect 21821 12189 21833 12223
rect 21867 12220 21879 12223
rect 21910 12220 21916 12232
rect 21867 12192 21916 12220
rect 21867 12189 21879 12192
rect 21821 12183 21879 12189
rect 18233 12155 18291 12161
rect 15396 12124 16252 12152
rect 15396 12084 15424 12124
rect 14476 12056 15424 12084
rect 16114 12044 16120 12096
rect 16172 12044 16178 12096
rect 16224 12084 16252 12124
rect 18233 12121 18245 12155
rect 18279 12121 18291 12155
rect 18233 12115 18291 12121
rect 20625 12155 20683 12161
rect 20625 12121 20637 12155
rect 20671 12152 20683 12155
rect 21836 12152 21864 12183
rect 21910 12180 21916 12192
rect 21968 12180 21974 12232
rect 23750 12180 23756 12232
rect 23808 12180 23814 12232
rect 24394 12180 24400 12232
rect 24452 12180 24458 12232
rect 24762 12180 24768 12232
rect 24820 12220 24826 12232
rect 24857 12223 24915 12229
rect 24857 12220 24869 12223
rect 24820 12192 24869 12220
rect 24820 12180 24826 12192
rect 24857 12189 24869 12192
rect 24903 12189 24915 12223
rect 24857 12183 24915 12189
rect 26418 12180 26424 12232
rect 26476 12180 26482 12232
rect 20671 12124 21864 12152
rect 20671 12121 20683 12124
rect 20625 12115 20683 12121
rect 23014 12084 23020 12096
rect 16224 12056 23020 12084
rect 23014 12044 23020 12056
rect 23072 12044 23078 12096
rect 23474 12044 23480 12096
rect 23532 12084 23538 12096
rect 23845 12087 23903 12093
rect 23845 12084 23857 12087
rect 23532 12056 23857 12084
rect 23532 12044 23538 12056
rect 23845 12053 23857 12056
rect 23891 12053 23903 12087
rect 23845 12047 23903 12053
rect 552 11994 27416 12016
rect 552 11942 3756 11994
rect 3808 11942 3820 11994
rect 3872 11942 3884 11994
rect 3936 11942 3948 11994
rect 4000 11942 4012 11994
rect 4064 11942 10472 11994
rect 10524 11942 10536 11994
rect 10588 11942 10600 11994
rect 10652 11942 10664 11994
rect 10716 11942 10728 11994
rect 10780 11942 17188 11994
rect 17240 11942 17252 11994
rect 17304 11942 17316 11994
rect 17368 11942 17380 11994
rect 17432 11942 17444 11994
rect 17496 11942 23904 11994
rect 23956 11942 23968 11994
rect 24020 11942 24032 11994
rect 24084 11942 24096 11994
rect 24148 11942 24160 11994
rect 24212 11942 27416 11994
rect 552 11920 27416 11942
rect 3602 11840 3608 11892
rect 3660 11880 3666 11892
rect 3973 11883 4031 11889
rect 3973 11880 3985 11883
rect 3660 11852 3985 11880
rect 3660 11840 3666 11852
rect 3973 11849 3985 11852
rect 4019 11849 4031 11883
rect 3973 11843 4031 11849
rect 4801 11883 4859 11889
rect 4801 11849 4813 11883
rect 4847 11880 4859 11883
rect 4890 11880 4896 11892
rect 4847 11852 4896 11880
rect 4847 11849 4859 11852
rect 4801 11843 4859 11849
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 5629 11883 5687 11889
rect 5629 11849 5641 11883
rect 5675 11880 5687 11883
rect 5902 11880 5908 11892
rect 5675 11852 5908 11880
rect 5675 11849 5687 11852
rect 5629 11843 5687 11849
rect 5902 11840 5908 11852
rect 5960 11840 5966 11892
rect 9950 11880 9956 11892
rect 8588 11852 9956 11880
rect 8588 11812 8616 11852
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 10045 11883 10103 11889
rect 10045 11849 10057 11883
rect 10091 11880 10103 11883
rect 10226 11880 10232 11892
rect 10091 11852 10232 11880
rect 10091 11849 10103 11852
rect 10045 11843 10103 11849
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 13170 11880 13176 11892
rect 10520 11852 13176 11880
rect 4816 11784 8616 11812
rect 4816 11756 4844 11784
rect 9582 11772 9588 11824
rect 9640 11812 9646 11824
rect 10520 11812 10548 11852
rect 13170 11840 13176 11852
rect 13228 11880 13234 11892
rect 13446 11880 13452 11892
rect 13228 11852 13452 11880
rect 13228 11840 13234 11852
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 13722 11840 13728 11892
rect 13780 11880 13786 11892
rect 13780 11852 14504 11880
rect 13780 11840 13786 11852
rect 9640 11784 10548 11812
rect 9640 11772 9646 11784
rect 12710 11772 12716 11824
rect 12768 11812 12774 11824
rect 12897 11815 12955 11821
rect 12897 11812 12909 11815
rect 12768 11784 12909 11812
rect 12768 11772 12774 11784
rect 12897 11781 12909 11784
rect 12943 11781 12955 11815
rect 14476 11812 14504 11852
rect 14550 11840 14556 11892
rect 14608 11880 14614 11892
rect 14921 11883 14979 11889
rect 14921 11880 14933 11883
rect 14608 11852 14933 11880
rect 14608 11840 14614 11852
rect 14921 11849 14933 11852
rect 14967 11849 14979 11883
rect 16390 11880 16396 11892
rect 14921 11843 14979 11849
rect 15028 11852 16396 11880
rect 15028 11812 15056 11852
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 16577 11883 16635 11889
rect 16577 11849 16589 11883
rect 16623 11880 16635 11883
rect 16942 11880 16948 11892
rect 16623 11852 16948 11880
rect 16623 11849 16635 11852
rect 16577 11843 16635 11849
rect 16942 11840 16948 11852
rect 17000 11840 17006 11892
rect 18414 11840 18420 11892
rect 18472 11880 18478 11892
rect 18693 11883 18751 11889
rect 18693 11880 18705 11883
rect 18472 11852 18705 11880
rect 18472 11840 18478 11852
rect 18693 11849 18705 11852
rect 18739 11849 18751 11883
rect 18693 11843 18751 11849
rect 20346 11840 20352 11892
rect 20404 11880 20410 11892
rect 21082 11880 21088 11892
rect 20404 11852 21088 11880
rect 20404 11840 20410 11852
rect 21082 11840 21088 11852
rect 21140 11880 21146 11892
rect 21361 11883 21419 11889
rect 21361 11880 21373 11883
rect 21140 11852 21373 11880
rect 21140 11840 21146 11852
rect 21361 11849 21373 11852
rect 21407 11849 21419 11883
rect 21361 11843 21419 11849
rect 23569 11883 23627 11889
rect 23569 11849 23581 11883
rect 23615 11880 23627 11883
rect 24394 11880 24400 11892
rect 23615 11852 24400 11880
rect 23615 11849 23627 11852
rect 23569 11843 23627 11849
rect 24394 11840 24400 11852
rect 24452 11840 24458 11892
rect 26418 11840 26424 11892
rect 26476 11840 26482 11892
rect 14476 11784 15056 11812
rect 18325 11815 18383 11821
rect 12897 11775 12955 11781
rect 18325 11781 18337 11815
rect 18371 11812 18383 11815
rect 19889 11815 19947 11821
rect 18371 11784 19288 11812
rect 18371 11781 18383 11784
rect 18325 11775 18383 11781
rect 4798 11704 4804 11756
rect 4856 11704 4862 11756
rect 7006 11744 7012 11756
rect 6932 11716 7012 11744
rect 3050 11636 3056 11688
rect 3108 11676 3114 11688
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 3108 11648 3801 11676
rect 3108 11636 3114 11648
rect 3789 11645 3801 11648
rect 3835 11645 3847 11679
rect 3789 11639 3847 11645
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11645 4031 11679
rect 3973 11639 4031 11645
rect 3988 11540 4016 11639
rect 4706 11636 4712 11688
rect 4764 11636 4770 11688
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11676 4951 11679
rect 5350 11676 5356 11688
rect 4939 11648 5356 11676
rect 4939 11645 4951 11648
rect 4893 11639 4951 11645
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 5445 11679 5503 11685
rect 5445 11645 5457 11679
rect 5491 11676 5503 11679
rect 5994 11676 6000 11688
rect 5491 11648 6000 11676
rect 5491 11645 5503 11648
rect 5445 11639 5503 11645
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 6638 11636 6644 11688
rect 6696 11636 6702 11688
rect 6932 11685 6960 11716
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 19260 11753 19288 11784
rect 19889 11781 19901 11815
rect 19935 11781 19947 11815
rect 19889 11775 19947 11781
rect 19245 11747 19303 11753
rect 19245 11713 19257 11747
rect 19291 11713 19303 11747
rect 19245 11707 19303 11713
rect 6917 11679 6975 11685
rect 6917 11645 6929 11679
rect 6963 11645 6975 11679
rect 6917 11639 6975 11645
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11676 8631 11679
rect 9122 11676 9128 11688
rect 8619 11648 9128 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 9122 11636 9128 11648
rect 9180 11676 9186 11688
rect 9306 11676 9312 11688
rect 9180 11648 9312 11676
rect 9180 11636 9186 11648
rect 9306 11636 9312 11648
rect 9364 11676 9370 11688
rect 13814 11685 13820 11688
rect 11425 11679 11483 11685
rect 11425 11676 11437 11679
rect 9364 11648 11437 11676
rect 9364 11636 9370 11648
rect 11072 11620 11100 11648
rect 11425 11645 11437 11648
rect 11471 11676 11483 11679
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11471 11648 11529 11676
rect 11471 11645 11483 11648
rect 11425 11639 11483 11645
rect 11517 11645 11529 11648
rect 11563 11676 11575 11679
rect 13541 11679 13599 11685
rect 11563 11648 13124 11676
rect 11563 11645 11575 11648
rect 11517 11639 11575 11645
rect 7009 11611 7067 11617
rect 7009 11577 7021 11611
rect 7055 11608 7067 11611
rect 7653 11611 7711 11617
rect 7653 11608 7665 11611
rect 7055 11580 7665 11608
rect 7055 11577 7067 11580
rect 7009 11571 7067 11577
rect 7653 11577 7665 11580
rect 7699 11608 7711 11611
rect 8386 11608 8392 11620
rect 7699 11580 8392 11608
rect 7699 11577 7711 11580
rect 7653 11571 7711 11577
rect 8386 11568 8392 11580
rect 8444 11568 8450 11620
rect 8478 11568 8484 11620
rect 8536 11608 8542 11620
rect 8818 11611 8876 11617
rect 8818 11608 8830 11611
rect 8536 11580 8830 11608
rect 8536 11568 8542 11580
rect 8818 11577 8830 11580
rect 8864 11577 8876 11611
rect 9858 11608 9864 11620
rect 8818 11571 8876 11577
rect 8956 11580 9864 11608
rect 7561 11543 7619 11549
rect 7561 11540 7573 11543
rect 3988 11512 7573 11540
rect 7561 11509 7573 11512
rect 7607 11540 7619 11543
rect 8956 11540 8984 11580
rect 9858 11568 9864 11580
rect 9916 11568 9922 11620
rect 10134 11568 10140 11620
rect 10192 11608 10198 11620
rect 10962 11608 10968 11620
rect 10192 11580 10968 11608
rect 10192 11568 10198 11580
rect 10962 11568 10968 11580
rect 11020 11568 11026 11620
rect 11054 11568 11060 11620
rect 11112 11568 11118 11620
rect 11180 11611 11238 11617
rect 11180 11577 11192 11611
rect 11226 11608 11238 11611
rect 11606 11608 11612 11620
rect 11226 11580 11612 11608
rect 11226 11577 11238 11580
rect 11180 11571 11238 11577
rect 11606 11568 11612 11580
rect 11664 11568 11670 11620
rect 11784 11611 11842 11617
rect 11784 11577 11796 11611
rect 11830 11608 11842 11611
rect 12066 11608 12072 11620
rect 11830 11580 12072 11608
rect 11830 11577 11842 11580
rect 11784 11571 11842 11577
rect 12066 11568 12072 11580
rect 12124 11568 12130 11620
rect 13096 11608 13124 11648
rect 13541 11645 13553 11679
rect 13587 11645 13599 11679
rect 13808 11676 13820 11685
rect 13775 11648 13820 11676
rect 13541 11639 13599 11645
rect 13808 11639 13820 11648
rect 13170 11608 13176 11620
rect 13096 11580 13176 11608
rect 13170 11568 13176 11580
rect 13228 11608 13234 11620
rect 13556 11608 13584 11639
rect 13814 11636 13820 11639
rect 13872 11636 13878 11688
rect 15194 11636 15200 11688
rect 15252 11676 15258 11688
rect 16945 11679 17003 11685
rect 16945 11676 16957 11679
rect 15252 11648 16957 11676
rect 15252 11636 15258 11648
rect 16945 11645 16957 11648
rect 16991 11645 17003 11679
rect 16945 11639 17003 11645
rect 17212 11679 17270 11685
rect 17212 11645 17224 11679
rect 17258 11676 17270 11679
rect 17678 11676 17684 11688
rect 17258 11648 17684 11676
rect 17258 11645 17270 11648
rect 17212 11639 17270 11645
rect 17678 11636 17684 11648
rect 17736 11636 17742 11688
rect 19904 11676 19932 11775
rect 21266 11704 21272 11756
rect 21324 11744 21330 11756
rect 21324 11716 22094 11744
rect 21324 11704 21330 11716
rect 21913 11679 21971 11685
rect 21913 11676 21925 11679
rect 19904 11648 21925 11676
rect 21913 11645 21925 11648
rect 21959 11645 21971 11679
rect 22066 11676 22094 11716
rect 23750 11704 23756 11756
rect 23808 11744 23814 11756
rect 24762 11744 24768 11756
rect 23808 11716 24768 11744
rect 23808 11704 23814 11716
rect 24762 11704 24768 11716
rect 24820 11744 24826 11756
rect 25041 11747 25099 11753
rect 25041 11744 25053 11747
rect 24820 11716 25053 11744
rect 24820 11704 24826 11716
rect 25041 11713 25053 11716
rect 25087 11713 25099 11747
rect 25041 11707 25099 11713
rect 22189 11679 22247 11685
rect 22189 11676 22201 11679
rect 22066 11648 22201 11676
rect 21913 11639 21971 11645
rect 22189 11645 22201 11648
rect 22235 11676 22247 11679
rect 23768 11676 23796 11704
rect 22235 11648 23796 11676
rect 22235 11645 22247 11648
rect 22189 11639 22247 11645
rect 24394 11636 24400 11688
rect 24452 11636 24458 11688
rect 13228 11580 13584 11608
rect 15464 11611 15522 11617
rect 13228 11568 13234 11580
rect 15464 11577 15476 11611
rect 15510 11608 15522 11611
rect 16114 11608 16120 11620
rect 15510 11580 16120 11608
rect 15510 11577 15522 11580
rect 15464 11571 15522 11577
rect 16114 11568 16120 11580
rect 16172 11568 16178 11620
rect 16482 11568 16488 11620
rect 16540 11608 16546 11620
rect 18046 11608 18052 11620
rect 16540 11580 18052 11608
rect 16540 11568 16546 11580
rect 18046 11568 18052 11580
rect 18104 11568 18110 11620
rect 21024 11611 21082 11617
rect 21024 11577 21036 11611
rect 21070 11608 21082 11611
rect 21634 11608 21640 11620
rect 21070 11580 21640 11608
rect 21070 11577 21082 11580
rect 21024 11571 21082 11577
rect 21634 11568 21640 11580
rect 21692 11568 21698 11620
rect 22456 11611 22514 11617
rect 22456 11577 22468 11611
rect 22502 11608 22514 11611
rect 23845 11611 23903 11617
rect 23845 11608 23857 11611
rect 22502 11580 23857 11608
rect 22502 11577 22514 11580
rect 22456 11571 22514 11577
rect 23845 11577 23857 11580
rect 23891 11577 23903 11611
rect 23845 11571 23903 11577
rect 25308 11611 25366 11617
rect 25308 11577 25320 11611
rect 25354 11608 25366 11611
rect 25590 11608 25596 11620
rect 25354 11580 25596 11608
rect 25354 11577 25366 11580
rect 25308 11571 25366 11577
rect 25590 11568 25596 11580
rect 25648 11568 25654 11620
rect 7607 11512 8984 11540
rect 7607 11509 7619 11512
rect 7561 11503 7619 11509
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 9582 11540 9588 11552
rect 9088 11512 9588 11540
rect 9088 11500 9094 11512
rect 9582 11500 9588 11512
rect 9640 11540 9646 11552
rect 9953 11543 10011 11549
rect 9953 11540 9965 11543
rect 9640 11512 9965 11540
rect 9640 11500 9646 11512
rect 9953 11509 9965 11512
rect 9999 11509 10011 11543
rect 9953 11503 10011 11509
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 16022 11540 16028 11552
rect 10376 11512 16028 11540
rect 10376 11500 10382 11512
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 552 11450 27576 11472
rect 552 11398 7114 11450
rect 7166 11398 7178 11450
rect 7230 11398 7242 11450
rect 7294 11398 7306 11450
rect 7358 11398 7370 11450
rect 7422 11398 13830 11450
rect 13882 11398 13894 11450
rect 13946 11398 13958 11450
rect 14010 11398 14022 11450
rect 14074 11398 14086 11450
rect 14138 11398 20546 11450
rect 20598 11398 20610 11450
rect 20662 11398 20674 11450
rect 20726 11398 20738 11450
rect 20790 11398 20802 11450
rect 20854 11398 27262 11450
rect 27314 11398 27326 11450
rect 27378 11398 27390 11450
rect 27442 11398 27454 11450
rect 27506 11398 27518 11450
rect 27570 11398 27576 11450
rect 552 11376 27576 11398
rect 4430 11296 4436 11348
rect 4488 11336 4494 11348
rect 4982 11336 4988 11348
rect 4488 11308 4988 11336
rect 4488 11296 4494 11308
rect 4982 11296 4988 11308
rect 5040 11296 5046 11348
rect 8386 11296 8392 11348
rect 8444 11336 8450 11348
rect 10226 11336 10232 11348
rect 8444 11308 10232 11336
rect 8444 11296 8450 11308
rect 10226 11296 10232 11308
rect 10284 11336 10290 11348
rect 10284 11308 10364 11336
rect 10284 11296 10290 11308
rect 3228 11271 3286 11277
rect 3228 11237 3240 11271
rect 3274 11268 3286 11271
rect 4525 11271 4583 11277
rect 4525 11268 4537 11271
rect 3274 11240 4537 11268
rect 3274 11237 3286 11240
rect 3228 11231 3286 11237
rect 4525 11237 4537 11240
rect 4571 11237 4583 11271
rect 10042 11268 10048 11280
rect 4525 11231 4583 11237
rect 5276 11240 5580 11268
rect 2682 11160 2688 11212
rect 2740 11200 2746 11212
rect 2961 11203 3019 11209
rect 2961 11200 2973 11203
rect 2740 11172 2973 11200
rect 2740 11160 2746 11172
rect 2961 11169 2973 11172
rect 3007 11169 3019 11203
rect 2961 11163 3019 11169
rect 4430 11160 4436 11212
rect 4488 11160 4494 11212
rect 4617 11203 4675 11209
rect 4617 11169 4629 11203
rect 4663 11169 4675 11203
rect 4617 11163 4675 11169
rect 4632 11132 4660 11163
rect 4982 11160 4988 11212
rect 5040 11160 5046 11212
rect 5166 11160 5172 11212
rect 5224 11160 5230 11212
rect 5276 11209 5304 11240
rect 5552 11212 5580 11240
rect 6104 11240 10048 11268
rect 5261 11203 5319 11209
rect 5261 11169 5273 11203
rect 5307 11169 5319 11203
rect 5261 11163 5319 11169
rect 5350 11160 5356 11212
rect 5408 11200 5414 11212
rect 5445 11203 5503 11209
rect 5445 11200 5457 11203
rect 5408 11172 5457 11200
rect 5408 11160 5414 11172
rect 5445 11169 5457 11172
rect 5491 11169 5503 11203
rect 5445 11163 5503 11169
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 5629 11203 5687 11209
rect 5629 11200 5641 11203
rect 5592 11172 5641 11200
rect 5592 11160 5598 11172
rect 5629 11169 5641 11172
rect 5675 11169 5687 11203
rect 5629 11163 5687 11169
rect 5718 11160 5724 11212
rect 5776 11200 5782 11212
rect 5813 11203 5871 11209
rect 5813 11200 5825 11203
rect 5776 11172 5825 11200
rect 5776 11160 5782 11172
rect 5813 11169 5825 11172
rect 5859 11169 5871 11203
rect 5813 11163 5871 11169
rect 5994 11160 6000 11212
rect 6052 11160 6058 11212
rect 6104 11209 6132 11240
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 10336 11277 10364 11308
rect 11606 11296 11612 11348
rect 11664 11296 11670 11348
rect 12618 11336 12624 11348
rect 11707 11308 12624 11336
rect 10321 11271 10379 11277
rect 10321 11237 10333 11271
rect 10367 11237 10379 11271
rect 10321 11231 10379 11237
rect 10870 11228 10876 11280
rect 10928 11268 10934 11280
rect 11707 11268 11735 11308
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 13078 11296 13084 11348
rect 13136 11296 13142 11348
rect 13446 11296 13452 11348
rect 13504 11296 13510 11348
rect 14553 11339 14611 11345
rect 14553 11305 14565 11339
rect 14599 11336 14611 11339
rect 14826 11336 14832 11348
rect 14599 11308 14832 11336
rect 14599 11305 14611 11308
rect 14553 11299 14611 11305
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 15470 11336 15476 11348
rect 15335 11308 15476 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 17313 11339 17371 11345
rect 17313 11305 17325 11339
rect 17359 11336 17371 11339
rect 17954 11336 17960 11348
rect 17359 11308 17960 11336
rect 17359 11305 17371 11308
rect 17313 11299 17371 11305
rect 17954 11296 17960 11308
rect 18012 11336 18018 11348
rect 18012 11308 19380 11336
rect 18012 11296 18018 11308
rect 10928 11240 11735 11268
rect 10928 11228 10934 11240
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 6914 11160 6920 11212
rect 6972 11160 6978 11212
rect 7184 11203 7242 11209
rect 7184 11169 7196 11203
rect 7230 11200 7242 11203
rect 7558 11200 7564 11212
rect 7230 11172 7564 11200
rect 7230 11169 7242 11172
rect 7184 11163 7242 11169
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 8294 11160 8300 11212
rect 8352 11200 8358 11212
rect 8662 11200 8668 11212
rect 8352 11172 8668 11200
rect 8352 11160 8358 11172
rect 8662 11160 8668 11172
rect 8720 11200 8726 11212
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 8720 11172 9045 11200
rect 8720 11160 8726 11172
rect 9033 11169 9045 11172
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 10980 11209 11008 11240
rect 12250 11228 12256 11280
rect 12308 11268 12314 11280
rect 13464 11268 13492 11296
rect 14921 11271 14979 11277
rect 14921 11268 14933 11271
rect 12308 11240 12664 11268
rect 13464 11240 14933 11268
rect 12308 11228 12314 11240
rect 10137 11203 10195 11209
rect 10137 11200 10149 11203
rect 9824 11172 10149 11200
rect 9824 11160 9830 11172
rect 10137 11169 10149 11172
rect 10183 11169 10195 11203
rect 10137 11163 10195 11169
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11169 11207 11203
rect 11149 11163 11207 11169
rect 11241 11203 11299 11209
rect 11241 11169 11253 11203
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 8389 11135 8447 11141
rect 4632 11104 5856 11132
rect 5828 11073 5856 11104
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 10505 11135 10563 11141
rect 10505 11101 10517 11135
rect 10551 11132 10563 11135
rect 11164 11132 11192 11163
rect 10551 11104 11192 11132
rect 10551 11101 10563 11104
rect 10505 11095 10563 11101
rect 5813 11067 5871 11073
rect 5813 11033 5825 11067
rect 5859 11033 5871 11067
rect 5813 11027 5871 11033
rect 8297 11067 8355 11073
rect 8297 11033 8309 11067
rect 8343 11064 8355 11067
rect 8404 11064 8432 11095
rect 8343 11036 8432 11064
rect 8343 11033 8355 11036
rect 8297 11027 8355 11033
rect 4341 10999 4399 11005
rect 4341 10965 4353 10999
rect 4387 10996 4399 10999
rect 5166 10996 5172 11008
rect 4387 10968 5172 10996
rect 4387 10965 4399 10968
rect 4341 10959 4399 10965
rect 5166 10956 5172 10968
rect 5224 10956 5230 11008
rect 5534 10956 5540 11008
rect 5592 10956 5598 11008
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 11256 10996 11284 11163
rect 11330 11160 11336 11212
rect 11388 11160 11394 11212
rect 12434 11160 12440 11212
rect 12492 11160 12498 11212
rect 12636 11209 12664 11240
rect 14921 11237 14933 11240
rect 14967 11268 14979 11271
rect 17862 11268 17868 11280
rect 14967 11240 17868 11268
rect 14967 11237 14979 11240
rect 14921 11231 14979 11237
rect 17862 11228 17868 11240
rect 17920 11228 17926 11280
rect 12621 11203 12679 11209
rect 12621 11169 12633 11203
rect 12667 11169 12679 11203
rect 12621 11163 12679 11169
rect 12713 11203 12771 11209
rect 12713 11169 12725 11203
rect 12759 11169 12771 11203
rect 12713 11163 12771 11169
rect 12728 11132 12756 11163
rect 12802 11160 12808 11212
rect 12860 11160 12866 11212
rect 13170 11160 13176 11212
rect 13228 11160 13234 11212
rect 13446 11209 13452 11212
rect 13440 11163 13452 11209
rect 13446 11160 13452 11163
rect 13504 11160 13510 11212
rect 14645 11203 14703 11209
rect 14645 11200 14657 11203
rect 14476 11172 14657 11200
rect 12728 11104 13216 11132
rect 13188 11076 13216 11104
rect 12710 11024 12716 11076
rect 12768 11064 12774 11076
rect 13078 11064 13084 11076
rect 12768 11036 13084 11064
rect 12768 11024 12774 11036
rect 13078 11024 13084 11036
rect 13136 11024 13142 11076
rect 13170 11024 13176 11076
rect 13228 11024 13234 11076
rect 14476 11064 14504 11172
rect 14645 11169 14657 11172
rect 14691 11169 14703 11203
rect 14645 11163 14703 11169
rect 14738 11203 14796 11209
rect 14738 11169 14750 11203
rect 14784 11169 14796 11203
rect 14738 11163 14796 11169
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 14752 11132 14780 11163
rect 14826 11160 14832 11212
rect 14884 11200 14890 11212
rect 15013 11203 15071 11209
rect 15013 11200 15025 11203
rect 14884 11172 15025 11200
rect 14884 11160 14890 11172
rect 15013 11169 15025 11172
rect 15059 11169 15071 11203
rect 15013 11163 15071 11169
rect 15102 11160 15108 11212
rect 15160 11209 15166 11212
rect 15160 11163 15168 11209
rect 15160 11160 15166 11163
rect 15470 11160 15476 11212
rect 15528 11200 15534 11212
rect 15746 11200 15752 11212
rect 15528 11172 15752 11200
rect 15528 11160 15534 11172
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 18437 11203 18495 11209
rect 18437 11169 18449 11203
rect 18483 11200 18495 11203
rect 18598 11200 18604 11212
rect 18483 11172 18604 11200
rect 18483 11169 18495 11172
rect 18437 11163 18495 11169
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 18693 11203 18751 11209
rect 18693 11169 18705 11203
rect 18739 11200 18751 11203
rect 19242 11200 19248 11212
rect 18739 11172 19248 11200
rect 18739 11169 18751 11172
rect 18693 11163 18751 11169
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 19352 11209 19380 11308
rect 19518 11296 19524 11348
rect 19576 11296 19582 11348
rect 20990 11336 20996 11348
rect 20180 11308 20996 11336
rect 19337 11203 19395 11209
rect 19337 11169 19349 11203
rect 19383 11169 19395 11203
rect 19337 11163 19395 11169
rect 19794 11160 19800 11212
rect 19852 11160 19858 11212
rect 19889 11203 19947 11209
rect 19889 11169 19901 11203
rect 19935 11169 19947 11203
rect 19889 11163 19947 11169
rect 14608 11104 14780 11132
rect 14608 11092 14614 11104
rect 18782 11092 18788 11144
rect 18840 11132 18846 11144
rect 19904 11132 19932 11163
rect 19978 11160 19984 11212
rect 20036 11160 20042 11212
rect 20180 11209 20208 11308
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 22646 11296 22652 11348
rect 22704 11296 22710 11348
rect 25501 11339 25559 11345
rect 25501 11305 25513 11339
rect 25547 11336 25559 11339
rect 26234 11336 26240 11348
rect 25547 11308 26240 11336
rect 25547 11305 25559 11308
rect 25501 11299 25559 11305
rect 26234 11296 26240 11308
rect 26292 11296 26298 11348
rect 20901 11271 20959 11277
rect 20901 11237 20913 11271
rect 20947 11268 20959 11271
rect 22186 11268 22192 11280
rect 20947 11240 22192 11268
rect 20947 11237 20959 11240
rect 20901 11231 20959 11237
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 20165 11203 20223 11209
rect 20165 11169 20177 11203
rect 20211 11169 20223 11203
rect 20165 11163 20223 11169
rect 20257 11203 20315 11209
rect 20257 11169 20269 11203
rect 20303 11169 20315 11203
rect 20257 11163 20315 11169
rect 20441 11203 20499 11209
rect 20441 11169 20453 11203
rect 20487 11169 20499 11203
rect 20441 11163 20499 11169
rect 20272 11132 20300 11163
rect 18840 11104 19932 11132
rect 20180 11104 20300 11132
rect 20456 11132 20484 11163
rect 20530 11160 20536 11212
rect 20588 11160 20594 11212
rect 20625 11203 20683 11209
rect 20625 11169 20637 11203
rect 20671 11200 20683 11203
rect 21082 11200 21088 11212
rect 20671 11172 21088 11200
rect 20671 11169 20683 11172
rect 20625 11163 20683 11169
rect 21082 11160 21088 11172
rect 21140 11160 21146 11212
rect 21266 11160 21272 11212
rect 21324 11160 21330 11212
rect 21542 11209 21548 11212
rect 21536 11163 21548 11209
rect 21542 11160 21548 11163
rect 21600 11160 21606 11212
rect 22664 11200 22692 11296
rect 26344 11240 26648 11268
rect 23293 11203 23351 11209
rect 23293 11200 23305 11203
rect 22664 11172 23305 11200
rect 23293 11169 23305 11172
rect 23339 11169 23351 11203
rect 23293 11163 23351 11169
rect 24388 11203 24446 11209
rect 24388 11169 24400 11203
rect 24434 11200 24446 11203
rect 24946 11200 24952 11212
rect 24434 11172 24952 11200
rect 24434 11169 24446 11172
rect 24388 11163 24446 11169
rect 24946 11160 24952 11172
rect 25004 11160 25010 11212
rect 26234 11160 26240 11212
rect 26292 11160 26298 11212
rect 20806 11132 20812 11144
rect 20456 11104 20812 11132
rect 18840 11092 18846 11104
rect 17586 11064 17592 11076
rect 14108 11036 17592 11064
rect 12158 10996 12164 11008
rect 7708 10968 12164 10996
rect 7708 10956 7714 10968
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 14108 10996 14136 11036
rect 17586 11024 17592 11036
rect 17644 11024 17650 11076
rect 20180 11008 20208 11104
rect 20806 11092 20812 11104
rect 20864 11092 20870 11144
rect 23750 11092 23756 11144
rect 23808 11132 23814 11144
rect 24121 11135 24179 11141
rect 24121 11132 24133 11135
rect 23808 11104 24133 11132
rect 23808 11092 23814 11104
rect 24121 11101 24133 11104
rect 24167 11101 24179 11135
rect 24121 11095 24179 11101
rect 25314 11092 25320 11144
rect 25372 11132 25378 11144
rect 26344 11132 26372 11240
rect 26620 11209 26648 11240
rect 26421 11203 26479 11209
rect 26421 11169 26433 11203
rect 26467 11169 26479 11203
rect 26421 11163 26479 11169
rect 26605 11203 26663 11209
rect 26605 11169 26617 11203
rect 26651 11169 26663 11203
rect 26605 11163 26663 11169
rect 26697 11203 26755 11209
rect 26697 11169 26709 11203
rect 26743 11169 26755 11203
rect 26697 11163 26755 11169
rect 26789 11203 26847 11209
rect 26789 11169 26801 11203
rect 26835 11200 26847 11203
rect 26878 11200 26884 11212
rect 26835 11172 26884 11200
rect 26835 11169 26847 11172
rect 26789 11163 26847 11169
rect 25372 11104 26372 11132
rect 25372 11092 25378 11104
rect 20346 11024 20352 11076
rect 20404 11064 20410 11076
rect 20530 11064 20536 11076
rect 20404 11036 20536 11064
rect 20404 11024 20410 11036
rect 20530 11024 20536 11036
rect 20588 11024 20594 11076
rect 25130 11024 25136 11076
rect 25188 11064 25194 11076
rect 25593 11067 25651 11073
rect 25593 11064 25605 11067
rect 25188 11036 25605 11064
rect 25188 11024 25194 11036
rect 25593 11033 25605 11036
rect 25639 11033 25651 11067
rect 26436 11064 26464 11163
rect 26712 11132 26740 11163
rect 26878 11160 26884 11172
rect 26936 11160 26942 11212
rect 25593 11027 25651 11033
rect 25700 11036 26464 11064
rect 26528 11104 26740 11132
rect 13412 10968 14136 10996
rect 13412 10956 13418 10968
rect 18046 10956 18052 11008
rect 18104 10996 18110 11008
rect 18785 10999 18843 11005
rect 18785 10996 18797 10999
rect 18104 10968 18797 10996
rect 18104 10956 18110 10968
rect 18785 10965 18797 10968
rect 18831 10965 18843 10999
rect 18785 10959 18843 10965
rect 20162 10956 20168 11008
rect 20220 10956 20226 11008
rect 22370 10956 22376 11008
rect 22428 10996 22434 11008
rect 22741 10999 22799 11005
rect 22741 10996 22753 10999
rect 22428 10968 22753 10996
rect 22428 10956 22434 10968
rect 22741 10965 22753 10968
rect 22787 10965 22799 10999
rect 22741 10959 22799 10965
rect 24486 10956 24492 11008
rect 24544 10996 24550 11008
rect 24762 10996 24768 11008
rect 24544 10968 24768 10996
rect 24544 10956 24550 10968
rect 24762 10956 24768 10968
rect 24820 10996 24826 11008
rect 25700 10996 25728 11036
rect 24820 10968 25728 10996
rect 24820 10956 24826 10968
rect 25774 10956 25780 11008
rect 25832 10996 25838 11008
rect 26528 10996 26556 11104
rect 25832 10968 26556 10996
rect 25832 10956 25838 10968
rect 27062 10956 27068 11008
rect 27120 10956 27126 11008
rect 552 10906 27416 10928
rect 552 10854 3756 10906
rect 3808 10854 3820 10906
rect 3872 10854 3884 10906
rect 3936 10854 3948 10906
rect 4000 10854 4012 10906
rect 4064 10854 10472 10906
rect 10524 10854 10536 10906
rect 10588 10854 10600 10906
rect 10652 10854 10664 10906
rect 10716 10854 10728 10906
rect 10780 10854 17188 10906
rect 17240 10854 17252 10906
rect 17304 10854 17316 10906
rect 17368 10854 17380 10906
rect 17432 10854 17444 10906
rect 17496 10854 23904 10906
rect 23956 10854 23968 10906
rect 24020 10854 24032 10906
rect 24084 10854 24096 10906
rect 24148 10854 24160 10906
rect 24212 10854 27416 10906
rect 552 10832 27416 10854
rect 7834 10792 7840 10804
rect 6380 10764 7840 10792
rect 6380 10733 6408 10764
rect 7834 10752 7840 10764
rect 7892 10752 7898 10804
rect 8404 10764 16528 10792
rect 6365 10727 6423 10733
rect 6365 10693 6377 10727
rect 6411 10693 6423 10727
rect 8018 10724 8024 10736
rect 6365 10687 6423 10693
rect 6840 10696 8024 10724
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 4632 10628 4813 10656
rect 4632 10600 4660 10628
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5040 10628 6316 10656
rect 5040 10616 5046 10628
rect 3142 10548 3148 10600
rect 3200 10588 3206 10600
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 3200 10560 3801 10588
rect 3200 10548 3206 10560
rect 3789 10557 3801 10560
rect 3835 10588 3847 10591
rect 3835 10560 4476 10588
rect 3835 10557 3847 10560
rect 3789 10551 3847 10557
rect 3881 10523 3939 10529
rect 3881 10489 3893 10523
rect 3927 10520 3939 10523
rect 4154 10520 4160 10532
rect 3927 10492 4160 10520
rect 3927 10489 3939 10492
rect 3881 10483 3939 10489
rect 4154 10480 4160 10492
rect 4212 10480 4218 10532
rect 4065 10455 4123 10461
rect 4065 10421 4077 10455
rect 4111 10452 4123 10455
rect 4338 10452 4344 10464
rect 4111 10424 4344 10452
rect 4111 10421 4123 10424
rect 4065 10415 4123 10421
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 4448 10452 4476 10560
rect 4614 10548 4620 10600
rect 4672 10548 4678 10600
rect 5445 10591 5503 10597
rect 5445 10588 5457 10591
rect 4816 10560 5457 10588
rect 4816 10532 4844 10560
rect 5445 10557 5457 10560
rect 5491 10557 5503 10591
rect 5445 10551 5503 10557
rect 5994 10548 6000 10600
rect 6052 10548 6058 10600
rect 6288 10597 6316 10628
rect 6840 10600 6868 10696
rect 8018 10684 8024 10696
rect 8076 10684 8082 10736
rect 7466 10656 7472 10668
rect 7208 10628 7472 10656
rect 6273 10591 6331 10597
rect 6273 10557 6285 10591
rect 6319 10557 6331 10591
rect 6273 10551 6331 10557
rect 6822 10548 6828 10600
rect 6880 10588 6886 10600
rect 6917 10591 6975 10597
rect 6917 10588 6929 10591
rect 6880 10560 6929 10588
rect 6880 10548 6886 10560
rect 6917 10557 6929 10560
rect 6963 10557 6975 10591
rect 6917 10551 6975 10557
rect 7006 10548 7012 10600
rect 7064 10588 7070 10600
rect 7208 10597 7236 10628
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 7101 10591 7159 10597
rect 7101 10588 7113 10591
rect 7064 10560 7113 10588
rect 7064 10548 7070 10560
rect 7101 10557 7113 10560
rect 7147 10557 7159 10591
rect 7101 10551 7159 10557
rect 7193 10591 7251 10597
rect 7193 10557 7205 10591
rect 7239 10557 7251 10591
rect 7193 10551 7251 10557
rect 7285 10591 7343 10597
rect 7285 10557 7297 10591
rect 7331 10588 7343 10591
rect 8294 10588 8300 10600
rect 7331 10560 8300 10588
rect 7331 10557 7343 10560
rect 7285 10551 7343 10557
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 4798 10480 4804 10532
rect 4856 10480 4862 10532
rect 5074 10480 5080 10532
rect 5132 10480 5138 10532
rect 5169 10523 5227 10529
rect 5169 10489 5181 10523
rect 5215 10520 5227 10523
rect 6012 10520 6040 10548
rect 8404 10520 8432 10764
rect 10042 10684 10048 10736
rect 10100 10684 10106 10736
rect 12529 10727 12587 10733
rect 12529 10693 12541 10727
rect 12575 10693 12587 10727
rect 16500 10724 16528 10764
rect 16574 10752 16580 10804
rect 16632 10752 16638 10804
rect 18138 10792 18144 10804
rect 17604 10764 18144 10792
rect 17604 10724 17632 10764
rect 18138 10752 18144 10764
rect 18196 10752 18202 10804
rect 18598 10752 18604 10804
rect 18656 10792 18662 10804
rect 18693 10795 18751 10801
rect 18693 10792 18705 10795
rect 18656 10764 18705 10792
rect 18656 10752 18662 10764
rect 18693 10761 18705 10764
rect 18739 10761 18751 10795
rect 18693 10755 18751 10761
rect 20806 10752 20812 10804
rect 20864 10752 20870 10804
rect 21542 10752 21548 10804
rect 21600 10752 21606 10804
rect 21634 10752 21640 10804
rect 21692 10752 21698 10804
rect 23385 10795 23443 10801
rect 23385 10761 23397 10795
rect 23431 10792 23443 10795
rect 24394 10792 24400 10804
rect 23431 10764 24400 10792
rect 23431 10761 23443 10764
rect 23385 10755 23443 10761
rect 24394 10752 24400 10764
rect 24452 10752 24458 10804
rect 24946 10752 24952 10804
rect 25004 10792 25010 10804
rect 25041 10795 25099 10801
rect 25041 10792 25053 10795
rect 25004 10764 25053 10792
rect 25004 10752 25010 10764
rect 25041 10761 25053 10764
rect 25087 10761 25099 10795
rect 25041 10755 25099 10761
rect 20073 10727 20131 10733
rect 20073 10724 20085 10727
rect 16500 10696 17632 10724
rect 17696 10696 20085 10724
rect 12529 10687 12587 10693
rect 8570 10616 8576 10668
rect 8628 10656 8634 10668
rect 9398 10656 9404 10668
rect 8628 10628 9404 10656
rect 8628 10616 8634 10628
rect 9398 10616 9404 10628
rect 9456 10656 9462 10668
rect 9456 10628 9536 10656
rect 9456 10616 9462 10628
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 8662 10588 8668 10600
rect 8527 10560 8668 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 9508 10597 9536 10628
rect 10318 10616 10324 10668
rect 10376 10616 10382 10668
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11149 10659 11207 10665
rect 11149 10656 11161 10659
rect 11112 10628 11161 10656
rect 11112 10616 11118 10628
rect 11149 10625 11161 10628
rect 11195 10625 11207 10659
rect 12544 10656 12572 10687
rect 12986 10656 12992 10668
rect 12544 10628 12992 10656
rect 11149 10619 11207 10625
rect 12986 10616 12992 10628
rect 13044 10656 13050 10668
rect 13173 10659 13231 10665
rect 13173 10656 13185 10659
rect 13044 10628 13185 10656
rect 13044 10616 13050 10628
rect 13173 10625 13185 10628
rect 13219 10625 13231 10659
rect 13173 10619 13231 10625
rect 14734 10616 14740 10668
rect 14792 10616 14798 10668
rect 14826 10616 14832 10668
rect 14884 10656 14890 10668
rect 17696 10656 17724 10696
rect 20073 10693 20085 10696
rect 20119 10724 20131 10727
rect 20162 10724 20168 10736
rect 20119 10696 20168 10724
rect 20119 10693 20131 10696
rect 20073 10687 20131 10693
rect 20162 10684 20168 10696
rect 20220 10724 20226 10736
rect 20220 10696 22784 10724
rect 20220 10684 20226 10696
rect 18230 10656 18236 10668
rect 14884 10628 17724 10656
rect 14884 10616 14890 10628
rect 9263 10591 9321 10597
rect 9263 10588 9275 10591
rect 8812 10560 9275 10588
rect 8812 10548 8818 10560
rect 9263 10557 9275 10560
rect 9309 10557 9321 10591
rect 9263 10551 9321 10557
rect 9493 10591 9551 10597
rect 9493 10557 9505 10591
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 9582 10548 9588 10600
rect 9640 10588 9646 10600
rect 9676 10591 9734 10597
rect 9676 10588 9688 10591
rect 9640 10560 9688 10588
rect 9640 10548 9646 10560
rect 9676 10557 9688 10560
rect 9722 10557 9734 10591
rect 9676 10551 9734 10557
rect 9769 10591 9827 10597
rect 9769 10557 9781 10591
rect 9815 10588 9827 10591
rect 11238 10588 11244 10600
rect 9815 10560 11244 10588
rect 9815 10557 9827 10560
rect 9769 10551 9827 10557
rect 11238 10548 11244 10560
rect 11296 10548 11302 10600
rect 15654 10548 15660 10600
rect 15712 10588 15718 10600
rect 17696 10597 17724 10628
rect 17972 10628 18236 10656
rect 16117 10591 16175 10597
rect 16117 10588 16129 10591
rect 15712 10560 16129 10588
rect 15712 10548 15718 10560
rect 16117 10557 16129 10560
rect 16163 10557 16175 10591
rect 16117 10551 16175 10557
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10557 16451 10591
rect 16393 10551 16451 10557
rect 17681 10591 17739 10597
rect 17681 10557 17693 10591
rect 17727 10557 17739 10591
rect 17681 10551 17739 10557
rect 9401 10523 9459 10529
rect 9401 10520 9413 10523
rect 5215 10492 5488 10520
rect 6012 10492 8432 10520
rect 9048 10492 9413 10520
rect 5215 10489 5227 10492
rect 5169 10483 5227 10489
rect 5460 10464 5488 10492
rect 4985 10455 5043 10461
rect 4985 10452 4997 10455
rect 4448 10424 4997 10452
rect 4985 10421 4997 10424
rect 5031 10421 5043 10455
rect 4985 10415 5043 10421
rect 5350 10412 5356 10464
rect 5408 10412 5414 10464
rect 5442 10412 5448 10464
rect 5500 10412 5506 10464
rect 7558 10412 7564 10464
rect 7616 10412 7622 10464
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 9048 10461 9076 10492
rect 9401 10489 9413 10492
rect 9447 10489 9459 10523
rect 9401 10483 9459 10489
rect 11416 10523 11474 10529
rect 11416 10489 11428 10523
rect 11462 10520 11474 10523
rect 11974 10520 11980 10532
rect 11462 10492 11980 10520
rect 11462 10489 11474 10492
rect 11416 10483 11474 10489
rect 11974 10480 11980 10492
rect 12032 10480 12038 10532
rect 12250 10480 12256 10532
rect 12308 10520 12314 10532
rect 12621 10523 12679 10529
rect 12621 10520 12633 10523
rect 12308 10492 12633 10520
rect 12308 10480 12314 10492
rect 12621 10489 12633 10492
rect 12667 10489 12679 10523
rect 16408 10520 16436 10551
rect 17862 10548 17868 10600
rect 17920 10548 17926 10600
rect 17972 10597 18000 10628
rect 18230 10616 18236 10628
rect 18288 10616 18294 10668
rect 18325 10659 18383 10665
rect 18325 10625 18337 10659
rect 18371 10656 18383 10659
rect 19245 10659 19303 10665
rect 19245 10656 19257 10659
rect 18371 10628 19257 10656
rect 18371 10625 18383 10628
rect 18325 10619 18383 10625
rect 19245 10625 19257 10628
rect 19291 10625 19303 10659
rect 19978 10656 19984 10668
rect 19245 10619 19303 10625
rect 19812 10628 19984 10656
rect 17957 10591 18015 10597
rect 17957 10557 17969 10591
rect 18003 10557 18015 10591
rect 17957 10551 18015 10557
rect 18046 10548 18052 10600
rect 18104 10548 18110 10600
rect 18138 10548 18144 10600
rect 18196 10588 18202 10600
rect 19812 10588 19840 10628
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 20530 10616 20536 10668
rect 20588 10656 20594 10668
rect 22094 10656 22100 10668
rect 20588 10628 22100 10656
rect 20588 10616 20594 10628
rect 18196 10560 19840 10588
rect 19889 10591 19947 10597
rect 18196 10548 18202 10560
rect 19889 10557 19901 10591
rect 19935 10588 19947 10591
rect 20162 10588 20168 10600
rect 19935 10560 20168 10588
rect 19935 10557 19947 10560
rect 19889 10551 19947 10557
rect 20162 10548 20168 10560
rect 20220 10548 20226 10600
rect 20346 10548 20352 10600
rect 20404 10548 20410 10600
rect 20625 10591 20683 10597
rect 20625 10557 20637 10591
rect 20671 10557 20683 10591
rect 20625 10551 20683 10557
rect 20901 10591 20959 10597
rect 20901 10557 20913 10591
rect 20947 10588 20959 10591
rect 20990 10588 20996 10600
rect 20947 10560 20996 10588
rect 20947 10557 20959 10560
rect 20901 10551 20959 10557
rect 17586 10520 17592 10532
rect 12621 10483 12679 10489
rect 16132 10492 17592 10520
rect 9033 10455 9091 10461
rect 9033 10452 9045 10455
rect 8352 10424 9045 10452
rect 8352 10412 8358 10424
rect 9033 10421 9045 10424
rect 9079 10421 9091 10455
rect 9033 10415 9091 10421
rect 9125 10455 9183 10461
rect 9125 10421 9137 10455
rect 9171 10452 9183 10455
rect 9214 10452 9220 10464
rect 9171 10424 9220 10452
rect 9171 10421 9183 10424
rect 9125 10415 9183 10421
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 9861 10455 9919 10461
rect 9861 10452 9873 10455
rect 9824 10424 9873 10452
rect 9824 10412 9830 10424
rect 9861 10421 9873 10424
rect 9907 10421 9919 10455
rect 9861 10415 9919 10421
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 14185 10455 14243 10461
rect 14185 10452 14197 10455
rect 13780 10424 14197 10452
rect 13780 10412 13786 10424
rect 14185 10421 14197 10424
rect 14231 10421 14243 10455
rect 14185 10415 14243 10421
rect 15378 10412 15384 10464
rect 15436 10452 15442 10464
rect 16132 10452 16160 10492
rect 17586 10480 17592 10492
rect 17644 10480 17650 10532
rect 19058 10480 19064 10532
rect 19116 10520 19122 10532
rect 20640 10520 20668 10551
rect 20990 10548 20996 10560
rect 21048 10548 21054 10600
rect 21082 10548 21088 10600
rect 21140 10548 21146 10600
rect 21192 10597 21220 10628
rect 22094 10616 22100 10628
rect 22152 10616 22158 10668
rect 22186 10616 22192 10668
rect 22244 10616 22250 10668
rect 22756 10656 22784 10696
rect 24762 10656 24768 10668
rect 22756 10628 24768 10656
rect 21177 10591 21235 10597
rect 21177 10557 21189 10591
rect 21223 10557 21235 10591
rect 21177 10551 21235 10557
rect 21269 10591 21327 10597
rect 21269 10557 21281 10591
rect 21315 10588 21327 10591
rect 22370 10588 22376 10600
rect 21315 10560 22376 10588
rect 21315 10557 21327 10560
rect 21269 10551 21327 10557
rect 22370 10548 22376 10560
rect 22428 10548 22434 10600
rect 22756 10597 22784 10628
rect 22741 10591 22799 10597
rect 22741 10557 22753 10591
rect 22787 10557 22799 10591
rect 22741 10551 22799 10557
rect 22922 10548 22928 10600
rect 22980 10548 22986 10600
rect 23017 10591 23075 10597
rect 23017 10557 23029 10591
rect 23063 10557 23075 10591
rect 23017 10551 23075 10557
rect 23109 10591 23167 10597
rect 23109 10557 23121 10591
rect 23155 10588 23167 10591
rect 23474 10588 23480 10600
rect 23155 10560 23480 10588
rect 23155 10557 23167 10560
rect 23109 10551 23167 10557
rect 22830 10520 22836 10532
rect 19116 10492 22836 10520
rect 19116 10480 19122 10492
rect 22830 10480 22836 10492
rect 22888 10480 22894 10532
rect 23032 10520 23060 10551
rect 23474 10548 23480 10560
rect 23532 10548 23538 10600
rect 24320 10597 24348 10628
rect 24762 10616 24768 10628
rect 24820 10616 24826 10668
rect 24949 10659 25007 10665
rect 24949 10625 24961 10659
rect 24995 10656 25007 10659
rect 25593 10659 25651 10665
rect 25593 10656 25605 10659
rect 24995 10628 25605 10656
rect 24995 10625 25007 10628
rect 24949 10619 25007 10625
rect 25593 10625 25605 10628
rect 25639 10625 25651 10659
rect 25593 10619 25651 10625
rect 26786 10616 26792 10668
rect 26844 10616 26850 10668
rect 24305 10591 24363 10597
rect 24305 10557 24317 10591
rect 24351 10557 24363 10591
rect 24305 10551 24363 10557
rect 24486 10548 24492 10600
rect 24544 10548 24550 10600
rect 24581 10591 24639 10597
rect 24581 10557 24593 10591
rect 24627 10557 24639 10591
rect 24581 10551 24639 10557
rect 24673 10591 24731 10597
rect 24673 10557 24685 10591
rect 24719 10588 24731 10591
rect 25130 10588 25136 10600
rect 24719 10560 25136 10588
rect 24719 10557 24731 10560
rect 24673 10551 24731 10557
rect 24596 10520 24624 10551
rect 25130 10548 25136 10560
rect 25188 10548 25194 10600
rect 24854 10520 24860 10532
rect 23032 10492 24860 10520
rect 15436 10424 16160 10452
rect 16209 10455 16267 10461
rect 15436 10412 15442 10424
rect 16209 10421 16221 10455
rect 16255 10452 16267 10455
rect 17678 10452 17684 10464
rect 16255 10424 17684 10452
rect 16255 10421 16267 10424
rect 16209 10415 16267 10421
rect 17678 10412 17684 10424
rect 17736 10412 17742 10464
rect 18874 10412 18880 10464
rect 18932 10452 18938 10464
rect 19794 10452 19800 10464
rect 18932 10424 19800 10452
rect 18932 10412 18938 10424
rect 19794 10412 19800 10424
rect 19852 10412 19858 10464
rect 20254 10412 20260 10464
rect 20312 10452 20318 10464
rect 20441 10455 20499 10461
rect 20441 10452 20453 10455
rect 20312 10424 20453 10452
rect 20312 10412 20318 10424
rect 20441 10421 20453 10424
rect 20487 10421 20499 10455
rect 20441 10415 20499 10421
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 23032 10452 23060 10492
rect 24854 10480 24860 10492
rect 24912 10520 24918 10532
rect 25774 10520 25780 10532
rect 24912 10492 25780 10520
rect 24912 10480 24918 10492
rect 25148 10464 25176 10492
rect 25774 10480 25780 10492
rect 25832 10480 25838 10532
rect 22152 10424 23060 10452
rect 22152 10412 22158 10424
rect 25130 10412 25136 10464
rect 25188 10412 25194 10464
rect 25222 10412 25228 10464
rect 25280 10452 25286 10464
rect 26145 10455 26203 10461
rect 26145 10452 26157 10455
rect 25280 10424 26157 10452
rect 25280 10412 25286 10424
rect 26145 10421 26157 10424
rect 26191 10421 26203 10455
rect 26145 10415 26203 10421
rect 552 10362 27576 10384
rect 552 10310 7114 10362
rect 7166 10310 7178 10362
rect 7230 10310 7242 10362
rect 7294 10310 7306 10362
rect 7358 10310 7370 10362
rect 7422 10310 13830 10362
rect 13882 10310 13894 10362
rect 13946 10310 13958 10362
rect 14010 10310 14022 10362
rect 14074 10310 14086 10362
rect 14138 10310 20546 10362
rect 20598 10310 20610 10362
rect 20662 10310 20674 10362
rect 20726 10310 20738 10362
rect 20790 10310 20802 10362
rect 20854 10310 27262 10362
rect 27314 10310 27326 10362
rect 27378 10310 27390 10362
rect 27442 10310 27454 10362
rect 27506 10310 27518 10362
rect 27570 10310 27576 10362
rect 552 10288 27576 10310
rect 3973 10251 4031 10257
rect 3973 10217 3985 10251
rect 4019 10248 4031 10251
rect 4614 10248 4620 10260
rect 4019 10220 4620 10248
rect 4019 10217 4031 10220
rect 3973 10211 4031 10217
rect 4614 10208 4620 10220
rect 4672 10248 4678 10260
rect 5258 10248 5264 10260
rect 4672 10220 5264 10248
rect 4672 10208 4678 10220
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 5500 10220 7236 10248
rect 5500 10208 5506 10220
rect 7208 10180 7236 10220
rect 8662 10208 8668 10260
rect 8720 10208 8726 10260
rect 11974 10208 11980 10260
rect 12032 10208 12038 10260
rect 12526 10208 12532 10260
rect 12584 10248 12590 10260
rect 12584 10220 13400 10248
rect 12584 10208 12590 10220
rect 10318 10180 10324 10192
rect 5000 10152 6224 10180
rect 5000 10124 5028 10152
rect 2593 10115 2651 10121
rect 2593 10081 2605 10115
rect 2639 10112 2651 10115
rect 2682 10112 2688 10124
rect 2639 10084 2688 10112
rect 2639 10081 2651 10084
rect 2593 10075 2651 10081
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 2866 10121 2872 10124
rect 2860 10112 2872 10121
rect 2827 10084 2872 10112
rect 2860 10075 2872 10084
rect 2866 10072 2872 10075
rect 2924 10072 2930 10124
rect 4062 10072 4068 10124
rect 4120 10072 4126 10124
rect 4157 10115 4215 10121
rect 4157 10081 4169 10115
rect 4203 10112 4215 10115
rect 4709 10115 4767 10121
rect 4709 10112 4721 10115
rect 4203 10084 4721 10112
rect 4203 10081 4215 10084
rect 4157 10075 4215 10081
rect 4709 10081 4721 10084
rect 4755 10112 4767 10115
rect 4982 10112 4988 10124
rect 4755 10084 4988 10112
rect 4755 10081 4767 10084
rect 4709 10075 4767 10081
rect 4982 10072 4988 10084
rect 5040 10072 5046 10124
rect 5258 10072 5264 10124
rect 5316 10112 5322 10124
rect 6196 10121 6224 10152
rect 7208 10152 10324 10180
rect 7208 10121 7236 10152
rect 10318 10140 10324 10152
rect 10376 10140 10382 10192
rect 11514 10140 11520 10192
rect 11572 10180 11578 10192
rect 12158 10180 12164 10192
rect 11572 10152 12164 10180
rect 11572 10140 11578 10152
rect 12158 10140 12164 10152
rect 12216 10180 12222 10192
rect 13372 10180 13400 10220
rect 13446 10208 13452 10260
rect 13504 10248 13510 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 13504 10220 13553 10248
rect 13504 10208 13510 10220
rect 13541 10217 13553 10220
rect 13587 10217 13599 10251
rect 13541 10211 13599 10217
rect 13648 10220 14412 10248
rect 13648 10180 13676 10220
rect 14384 10180 14412 10220
rect 15194 10208 15200 10260
rect 15252 10208 15258 10260
rect 15396 10220 16436 10248
rect 15396 10180 15424 10220
rect 12216 10152 13308 10180
rect 13372 10152 13676 10180
rect 13740 10152 13952 10180
rect 14384 10152 15424 10180
rect 15565 10183 15623 10189
rect 12216 10140 12222 10152
rect 7558 10121 7564 10124
rect 5997 10115 6055 10121
rect 5997 10112 6009 10115
rect 5316 10084 6009 10112
rect 5316 10072 5322 10084
rect 5997 10081 6009 10084
rect 6043 10081 6055 10115
rect 5997 10075 6055 10081
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10081 7251 10115
rect 7193 10075 7251 10081
rect 7552 10075 7564 10121
rect 7558 10072 7564 10075
rect 7616 10072 7622 10124
rect 9122 10072 9128 10124
rect 9180 10072 9186 10124
rect 9398 10121 9404 10124
rect 9392 10075 9404 10121
rect 9398 10072 9404 10075
rect 9456 10072 9462 10124
rect 12250 10072 12256 10124
rect 12308 10072 12314 10124
rect 12360 10121 12388 10152
rect 12345 10115 12403 10121
rect 12345 10081 12357 10115
rect 12391 10081 12403 10115
rect 12345 10075 12403 10081
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10112 12495 10115
rect 12526 10112 12532 10124
rect 12483 10084 12532 10112
rect 12483 10081 12495 10084
rect 12437 10075 12495 10081
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 12621 10115 12679 10121
rect 12621 10081 12633 10115
rect 12667 10112 12679 10115
rect 12802 10112 12808 10124
rect 12667 10084 12808 10112
rect 12667 10081 12679 10084
rect 12621 10075 12679 10081
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 13096 10121 13124 10152
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10081 13047 10115
rect 12989 10075 13047 10081
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10081 13139 10115
rect 13081 10075 13139 10081
rect 13173 10115 13231 10121
rect 13173 10081 13185 10115
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 4080 9976 4108 10072
rect 4338 10004 4344 10056
rect 4396 10004 4402 10056
rect 4617 10047 4675 10053
rect 4617 10044 4629 10047
rect 4448 10016 4629 10044
rect 4448 9976 4476 10016
rect 4617 10013 4629 10016
rect 4663 10044 4675 10047
rect 4798 10044 4804 10056
rect 4663 10016 4804 10044
rect 4663 10013 4675 10016
rect 4617 10007 4675 10013
rect 4798 10004 4804 10016
rect 4856 10044 4862 10056
rect 4856 10016 6040 10044
rect 4856 10004 4862 10016
rect 4080 9948 4476 9976
rect 4246 9868 4252 9920
rect 4304 9868 4310 9920
rect 4338 9868 4344 9920
rect 4396 9908 4402 9920
rect 4433 9911 4491 9917
rect 4433 9908 4445 9911
rect 4396 9880 4445 9908
rect 4396 9868 4402 9880
rect 4433 9877 4445 9880
rect 4479 9877 4491 9911
rect 4433 9871 4491 9877
rect 5810 9868 5816 9920
rect 5868 9868 5874 9920
rect 6012 9917 6040 10016
rect 6914 10004 6920 10056
rect 6972 10044 6978 10056
rect 7285 10047 7343 10053
rect 7285 10044 7297 10047
rect 6972 10016 7297 10044
rect 6972 10004 6978 10016
rect 7285 10013 7297 10016
rect 7331 10013 7343 10047
rect 7285 10007 7343 10013
rect 11238 10004 11244 10056
rect 11296 10004 11302 10056
rect 13004 10044 13032 10075
rect 11992 10016 13032 10044
rect 11992 9920 12020 10016
rect 12158 9936 12164 9988
rect 12216 9976 12222 9988
rect 13188 9976 13216 10075
rect 13280 10044 13308 10152
rect 13354 10072 13360 10124
rect 13412 10072 13418 10124
rect 13446 10044 13452 10056
rect 13280 10016 13452 10044
rect 13446 10004 13452 10016
rect 13504 10044 13510 10056
rect 13740 10044 13768 10152
rect 13814 10121 13820 10124
rect 13797 10115 13820 10121
rect 13797 10081 13809 10115
rect 13797 10075 13820 10081
rect 13814 10072 13820 10075
rect 13872 10072 13878 10124
rect 13924 10121 13952 10152
rect 15565 10149 15577 10183
rect 15611 10180 15623 10183
rect 16298 10180 16304 10192
rect 15611 10152 16304 10180
rect 15611 10149 15623 10152
rect 15565 10143 15623 10149
rect 16298 10140 16304 10152
rect 16356 10140 16362 10192
rect 16408 10180 16436 10220
rect 16666 10208 16672 10260
rect 16724 10248 16730 10260
rect 17034 10248 17040 10260
rect 16724 10220 17040 10248
rect 16724 10208 16730 10220
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 17678 10208 17684 10260
rect 17736 10208 17742 10260
rect 17862 10208 17868 10260
rect 17920 10248 17926 10260
rect 18969 10251 19027 10257
rect 18969 10248 18981 10251
rect 17920 10220 18981 10248
rect 17920 10208 17926 10220
rect 18969 10217 18981 10220
rect 19015 10217 19027 10251
rect 18969 10211 19027 10217
rect 19058 10208 19064 10260
rect 19116 10248 19122 10260
rect 19889 10251 19947 10257
rect 19116 10220 19748 10248
rect 19116 10208 19122 10220
rect 19521 10183 19579 10189
rect 19521 10180 19533 10183
rect 16408 10152 19533 10180
rect 19521 10149 19533 10152
rect 19567 10149 19579 10183
rect 19521 10143 19579 10149
rect 13909 10115 13967 10121
rect 13909 10081 13921 10115
rect 13955 10081 13967 10115
rect 13909 10075 13967 10081
rect 14022 10115 14080 10121
rect 14022 10081 14034 10115
rect 14068 10112 14080 10115
rect 14068 10084 14136 10112
rect 14068 10081 14080 10084
rect 14022 10075 14080 10081
rect 13504 10016 13768 10044
rect 14108 10044 14136 10084
rect 14182 10072 14188 10124
rect 14240 10112 14246 10124
rect 14826 10112 14832 10124
rect 14240 10084 14832 10112
rect 14240 10072 14246 10084
rect 14826 10072 14832 10084
rect 14884 10072 14890 10124
rect 15378 10072 15384 10124
rect 15436 10072 15442 10124
rect 15654 10072 15660 10124
rect 15712 10072 15718 10124
rect 15746 10072 15752 10124
rect 15804 10072 15810 10124
rect 15933 10115 15991 10121
rect 15933 10081 15945 10115
rect 15979 10112 15991 10115
rect 17034 10112 17040 10124
rect 15979 10084 17040 10112
rect 15979 10081 15991 10084
rect 15933 10075 15991 10081
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 18598 10072 18604 10124
rect 18656 10072 18662 10124
rect 18785 10115 18843 10121
rect 18785 10081 18797 10115
rect 18831 10081 18843 10115
rect 18785 10075 18843 10081
rect 14108 10016 14964 10044
rect 13504 10004 13510 10016
rect 12216 9948 13216 9976
rect 12216 9936 12222 9948
rect 13354 9936 13360 9988
rect 13412 9976 13418 9988
rect 14182 9976 14188 9988
rect 13412 9948 14188 9976
rect 13412 9936 13418 9948
rect 14182 9936 14188 9948
rect 14240 9936 14246 9988
rect 14936 9976 14964 10016
rect 15010 10004 15016 10056
rect 15068 10044 15074 10056
rect 15672 10044 15700 10072
rect 15068 10016 15700 10044
rect 15841 10047 15899 10053
rect 15068 10004 15074 10016
rect 15841 10013 15853 10047
rect 15887 10044 15899 10047
rect 16209 10047 16267 10053
rect 16209 10044 16221 10047
rect 15887 10016 16221 10044
rect 15887 10013 15899 10016
rect 15841 10007 15899 10013
rect 16209 10013 16221 10016
rect 16255 10013 16267 10047
rect 16209 10007 16267 10013
rect 16298 10004 16304 10056
rect 16356 10044 16362 10056
rect 16945 10047 17003 10053
rect 16945 10044 16957 10047
rect 16356 10016 16957 10044
rect 16356 10004 16362 10016
rect 16945 10013 16957 10016
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 18230 10004 18236 10056
rect 18288 10004 18294 10056
rect 18417 9979 18475 9985
rect 18417 9976 18429 9979
rect 14936 9948 18429 9976
rect 18417 9945 18429 9948
rect 18463 9945 18475 9979
rect 18800 9976 18828 10075
rect 18874 10072 18880 10124
rect 18932 10072 18938 10124
rect 19058 10072 19064 10124
rect 19116 10112 19122 10124
rect 19153 10115 19211 10121
rect 19153 10112 19165 10115
rect 19116 10084 19165 10112
rect 19116 10072 19122 10084
rect 19153 10081 19165 10084
rect 19199 10081 19211 10115
rect 19153 10075 19211 10081
rect 19334 10072 19340 10124
rect 19392 10072 19398 10124
rect 19720 10121 19748 10220
rect 19889 10217 19901 10251
rect 19935 10248 19947 10251
rect 20990 10248 20996 10260
rect 19935 10220 20996 10248
rect 19935 10217 19947 10220
rect 19889 10211 19947 10217
rect 20990 10208 20996 10220
rect 21048 10208 21054 10260
rect 21082 10208 21088 10260
rect 21140 10248 21146 10260
rect 21269 10251 21327 10257
rect 21269 10248 21281 10251
rect 21140 10220 21281 10248
rect 21140 10208 21146 10220
rect 21269 10217 21281 10220
rect 21315 10217 21327 10251
rect 22278 10248 22284 10260
rect 21269 10211 21327 10217
rect 21652 10220 22284 10248
rect 20717 10183 20775 10189
rect 20717 10149 20729 10183
rect 20763 10180 20775 10183
rect 21358 10180 21364 10192
rect 20763 10152 21364 10180
rect 20763 10149 20775 10152
rect 20717 10143 20775 10149
rect 21358 10140 21364 10152
rect 21416 10140 21422 10192
rect 21652 10180 21680 10220
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 22922 10208 22928 10260
rect 22980 10248 22986 10260
rect 23109 10251 23167 10257
rect 23109 10248 23121 10251
rect 22980 10220 23121 10248
rect 22980 10208 22986 10220
rect 23109 10217 23121 10220
rect 23155 10217 23167 10251
rect 23109 10211 23167 10217
rect 23477 10251 23535 10257
rect 23477 10217 23489 10251
rect 23523 10248 23535 10251
rect 24394 10248 24400 10260
rect 23523 10220 24400 10248
rect 23523 10217 23535 10220
rect 23477 10211 23535 10217
rect 24394 10208 24400 10220
rect 24452 10208 24458 10260
rect 24486 10208 24492 10260
rect 24544 10248 24550 10260
rect 24765 10251 24823 10257
rect 24765 10248 24777 10251
rect 24544 10220 24777 10248
rect 24544 10208 24550 10220
rect 24765 10217 24777 10220
rect 24811 10217 24823 10251
rect 24765 10211 24823 10217
rect 25590 10208 25596 10260
rect 25648 10208 25654 10260
rect 21560 10152 21680 10180
rect 21744 10152 23612 10180
rect 19429 10115 19487 10121
rect 19429 10081 19441 10115
rect 19475 10081 19487 10115
rect 19429 10075 19487 10081
rect 19705 10115 19763 10121
rect 19705 10081 19717 10115
rect 19751 10081 19763 10115
rect 19705 10075 19763 10081
rect 18892 10044 18920 10072
rect 19444 10044 19472 10075
rect 19978 10072 19984 10124
rect 20036 10072 20042 10124
rect 20162 10072 20168 10124
rect 20220 10072 20226 10124
rect 20346 10072 20352 10124
rect 20404 10112 20410 10124
rect 20625 10115 20683 10121
rect 20625 10112 20637 10115
rect 20404 10084 20637 10112
rect 20404 10072 20410 10084
rect 20625 10081 20637 10084
rect 20671 10081 20683 10115
rect 20625 10075 20683 10081
rect 20364 10044 20392 10072
rect 18892 10016 20392 10044
rect 20640 9976 20668 10075
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20864 10084 20913 10112
rect 20864 10072 20870 10084
rect 20901 10081 20913 10084
rect 20947 10112 20959 10115
rect 21453 10115 21511 10121
rect 21453 10112 21465 10115
rect 20947 10084 21465 10112
rect 20947 10081 20959 10084
rect 20901 10075 20959 10081
rect 21453 10081 21465 10084
rect 21499 10081 21511 10115
rect 21453 10075 21511 10081
rect 21085 10047 21143 10053
rect 21085 10013 21097 10047
rect 21131 10044 21143 10047
rect 21560 10044 21588 10152
rect 21744 10124 21772 10152
rect 21634 10072 21640 10124
rect 21692 10072 21698 10124
rect 21726 10072 21732 10124
rect 21784 10072 21790 10124
rect 22830 10072 22836 10124
rect 22888 10112 22894 10124
rect 23584 10121 23612 10152
rect 23658 10140 23664 10192
rect 23716 10180 23722 10192
rect 23845 10183 23903 10189
rect 23845 10180 23857 10183
rect 23716 10152 23857 10180
rect 23716 10140 23722 10152
rect 23845 10149 23857 10152
rect 23891 10149 23903 10183
rect 24213 10183 24271 10189
rect 23845 10143 23903 10149
rect 23952 10152 24164 10180
rect 23293 10115 23351 10121
rect 23293 10112 23305 10115
rect 22888 10084 23305 10112
rect 22888 10072 22894 10084
rect 23293 10081 23305 10084
rect 23339 10081 23351 10115
rect 23293 10075 23351 10081
rect 23569 10115 23627 10121
rect 23569 10081 23581 10115
rect 23615 10112 23627 10115
rect 23753 10115 23811 10121
rect 23753 10112 23765 10115
rect 23615 10084 23765 10112
rect 23615 10081 23627 10084
rect 23569 10075 23627 10081
rect 23753 10081 23765 10084
rect 23799 10112 23811 10115
rect 23952 10112 23980 10152
rect 23799 10084 23980 10112
rect 24029 10115 24087 10121
rect 23799 10081 23811 10084
rect 23753 10075 23811 10081
rect 24029 10081 24041 10115
rect 24075 10081 24087 10115
rect 24136 10112 24164 10152
rect 24213 10149 24225 10183
rect 24259 10180 24271 10183
rect 25314 10180 25320 10192
rect 24259 10152 25320 10180
rect 24259 10149 24271 10152
rect 24213 10143 24271 10149
rect 25314 10140 25320 10152
rect 25372 10140 25378 10192
rect 24302 10112 24308 10124
rect 24136 10084 24308 10112
rect 24029 10075 24087 10081
rect 21131 10016 21588 10044
rect 23308 10044 23336 10075
rect 24044 10044 24072 10075
rect 24302 10072 24308 10084
rect 24360 10072 24366 10124
rect 24397 10115 24455 10121
rect 24397 10081 24409 10115
rect 24443 10112 24455 10115
rect 24486 10112 24492 10124
rect 24443 10084 24492 10112
rect 24443 10081 24455 10084
rect 24397 10075 24455 10081
rect 24486 10072 24492 10084
rect 24544 10072 24550 10124
rect 24581 10115 24639 10121
rect 24581 10081 24593 10115
rect 24627 10081 24639 10115
rect 24581 10075 24639 10081
rect 24596 10044 24624 10075
rect 24762 10072 24768 10124
rect 24820 10112 24826 10124
rect 24857 10115 24915 10121
rect 24857 10112 24869 10115
rect 24820 10084 24869 10112
rect 24820 10072 24826 10084
rect 24857 10081 24869 10084
rect 24903 10081 24915 10115
rect 24857 10075 24915 10081
rect 25041 10115 25099 10121
rect 25041 10081 25053 10115
rect 25087 10081 25099 10115
rect 25041 10075 25099 10081
rect 25056 10044 25084 10075
rect 25130 10072 25136 10124
rect 25188 10072 25194 10124
rect 25222 10072 25228 10124
rect 25280 10072 25286 10124
rect 26237 10115 26295 10121
rect 26237 10081 26249 10115
rect 26283 10112 26295 10115
rect 27062 10112 27068 10124
rect 26283 10084 27068 10112
rect 26283 10081 26295 10084
rect 26237 10075 26295 10081
rect 27062 10072 27068 10084
rect 27120 10072 27126 10124
rect 26878 10044 26884 10056
rect 23308 10016 24164 10044
rect 21131 10013 21143 10016
rect 21085 10007 21143 10013
rect 21726 9976 21732 9988
rect 18800 9948 19334 9976
rect 20640 9948 21732 9976
rect 18417 9939 18475 9945
rect 5997 9911 6055 9917
rect 5997 9877 6009 9911
rect 6043 9877 6055 9911
rect 5997 9871 6055 9877
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7009 9911 7067 9917
rect 7009 9908 7021 9911
rect 6972 9880 7021 9908
rect 6972 9868 6978 9880
rect 7009 9877 7021 9880
rect 7055 9877 7067 9911
rect 7009 9871 7067 9877
rect 10318 9868 10324 9920
rect 10376 9908 10382 9920
rect 10505 9911 10563 9917
rect 10505 9908 10517 9911
rect 10376 9880 10517 9908
rect 10376 9868 10382 9880
rect 10505 9877 10517 9880
rect 10551 9877 10563 9911
rect 10505 9871 10563 9877
rect 11885 9911 11943 9917
rect 11885 9877 11897 9911
rect 11931 9908 11943 9911
rect 11974 9908 11980 9920
rect 11931 9880 11980 9908
rect 11931 9877 11943 9880
rect 11885 9871 11943 9877
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 12710 9868 12716 9920
rect 12768 9868 12774 9920
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 13372 9908 13400 9936
rect 12860 9880 13400 9908
rect 12860 9868 12866 9880
rect 16850 9868 16856 9920
rect 16908 9868 16914 9920
rect 17589 9911 17647 9917
rect 17589 9877 17601 9911
rect 17635 9908 17647 9911
rect 17678 9908 17684 9920
rect 17635 9880 17684 9908
rect 17635 9877 17647 9880
rect 17589 9871 17647 9877
rect 17678 9868 17684 9880
rect 17736 9868 17742 9920
rect 17862 9868 17868 9920
rect 17920 9908 17926 9920
rect 18874 9908 18880 9920
rect 17920 9880 18880 9908
rect 17920 9868 17926 9880
rect 18874 9868 18880 9880
rect 18932 9868 18938 9920
rect 19306 9908 19334 9948
rect 21726 9936 21732 9948
rect 21784 9936 21790 9988
rect 24136 9976 24164 10016
rect 24596 10016 24900 10044
rect 25056 10016 26884 10044
rect 24596 9976 24624 10016
rect 24872 9988 24900 10016
rect 26878 10004 26884 10016
rect 26936 10004 26942 10056
rect 26973 10047 27031 10053
rect 26973 10013 26985 10047
rect 27019 10013 27031 10047
rect 26973 10007 27031 10013
rect 24136 9948 24624 9976
rect 24854 9936 24860 9988
rect 24912 9936 24918 9988
rect 25501 9979 25559 9985
rect 25501 9945 25513 9979
rect 25547 9976 25559 9979
rect 26988 9976 27016 10007
rect 25547 9948 27016 9976
rect 25547 9945 25559 9948
rect 25501 9939 25559 9945
rect 19610 9908 19616 9920
rect 19306 9880 19616 9908
rect 19610 9868 19616 9880
rect 19668 9868 19674 9920
rect 19794 9868 19800 9920
rect 19852 9908 19858 9920
rect 20441 9911 20499 9917
rect 20441 9908 20453 9911
rect 19852 9880 20453 9908
rect 19852 9868 19858 9880
rect 20441 9877 20453 9880
rect 20487 9908 20499 9911
rect 23474 9908 23480 9920
rect 20487 9880 23480 9908
rect 20487 9877 20499 9880
rect 20441 9871 20499 9877
rect 23474 9868 23480 9880
rect 23532 9868 23538 9920
rect 24486 9868 24492 9920
rect 24544 9908 24550 9920
rect 25130 9908 25136 9920
rect 24544 9880 25136 9908
rect 24544 9868 24550 9880
rect 25130 9868 25136 9880
rect 25188 9868 25194 9920
rect 25774 9868 25780 9920
rect 25832 9908 25838 9920
rect 26421 9911 26479 9917
rect 26421 9908 26433 9911
rect 25832 9880 26433 9908
rect 25832 9868 25838 9880
rect 26421 9877 26433 9880
rect 26467 9877 26479 9911
rect 26421 9871 26479 9877
rect 552 9818 27416 9840
rect 552 9766 3756 9818
rect 3808 9766 3820 9818
rect 3872 9766 3884 9818
rect 3936 9766 3948 9818
rect 4000 9766 4012 9818
rect 4064 9766 10472 9818
rect 10524 9766 10536 9818
rect 10588 9766 10600 9818
rect 10652 9766 10664 9818
rect 10716 9766 10728 9818
rect 10780 9766 17188 9818
rect 17240 9766 17252 9818
rect 17304 9766 17316 9818
rect 17368 9766 17380 9818
rect 17432 9766 17444 9818
rect 17496 9766 23904 9818
rect 23956 9766 23968 9818
rect 24020 9766 24032 9818
rect 24084 9766 24096 9818
rect 24148 9766 24160 9818
rect 24212 9766 27416 9818
rect 552 9744 27416 9766
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 3881 9707 3939 9713
rect 3881 9704 3893 9707
rect 2924 9676 3893 9704
rect 2924 9664 2930 9676
rect 3881 9673 3893 9676
rect 3927 9673 3939 9707
rect 3881 9667 3939 9673
rect 6181 9707 6239 9713
rect 6181 9673 6193 9707
rect 6227 9704 6239 9707
rect 7006 9704 7012 9716
rect 6227 9676 7012 9704
rect 6227 9673 6239 9676
rect 6181 9667 6239 9673
rect 7006 9664 7012 9676
rect 7064 9664 7070 9716
rect 7558 9664 7564 9716
rect 7616 9664 7622 9716
rect 9398 9664 9404 9716
rect 9456 9704 9462 9716
rect 9585 9707 9643 9713
rect 9585 9704 9597 9707
rect 9456 9676 9597 9704
rect 9456 9664 9462 9676
rect 9585 9673 9597 9676
rect 9631 9673 9643 9707
rect 11238 9704 11244 9716
rect 9585 9667 9643 9673
rect 10980 9676 11244 9704
rect 3605 9639 3663 9645
rect 3605 9605 3617 9639
rect 3651 9636 3663 9639
rect 4154 9636 4160 9648
rect 3651 9608 4160 9636
rect 3651 9605 3663 9608
rect 3605 9599 3663 9605
rect 4154 9596 4160 9608
rect 4212 9596 4218 9648
rect 4893 9639 4951 9645
rect 4893 9605 4905 9639
rect 4939 9636 4951 9639
rect 5534 9636 5540 9648
rect 4939 9608 5540 9636
rect 4939 9605 4951 9608
rect 4893 9599 4951 9605
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 5629 9639 5687 9645
rect 5629 9605 5641 9639
rect 5675 9636 5687 9639
rect 5718 9636 5724 9648
rect 5675 9608 5724 9636
rect 5675 9605 5687 9608
rect 5629 9599 5687 9605
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 10505 9639 10563 9645
rect 10505 9605 10517 9639
rect 10551 9636 10563 9639
rect 10980 9636 11008 9676
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 13170 9664 13176 9716
rect 13228 9704 13234 9716
rect 15470 9704 15476 9716
rect 13228 9676 15476 9704
rect 13228 9664 13234 9676
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 16117 9707 16175 9713
rect 16117 9673 16129 9707
rect 16163 9704 16175 9707
rect 16298 9704 16304 9716
rect 16163 9676 16304 9704
rect 16163 9673 16175 9676
rect 16117 9667 16175 9673
rect 16298 9664 16304 9676
rect 16356 9664 16362 9716
rect 20438 9704 20444 9716
rect 16592 9676 20444 9704
rect 10551 9608 11008 9636
rect 10551 9605 10563 9608
rect 10505 9599 10563 9605
rect 13262 9596 13268 9648
rect 13320 9636 13326 9648
rect 13357 9639 13415 9645
rect 13357 9636 13369 9639
rect 13320 9608 13369 9636
rect 13320 9596 13326 9608
rect 13357 9605 13369 9608
rect 13403 9605 13415 9639
rect 16592 9636 16620 9676
rect 20438 9664 20444 9676
rect 20496 9664 20502 9716
rect 23658 9664 23664 9716
rect 23716 9704 23722 9716
rect 25222 9704 25228 9716
rect 23716 9676 25228 9704
rect 23716 9664 23722 9676
rect 25222 9664 25228 9676
rect 25280 9664 25286 9716
rect 26786 9664 26792 9716
rect 26844 9704 26850 9716
rect 26881 9707 26939 9713
rect 26881 9704 26893 9707
rect 26844 9676 26893 9704
rect 26844 9664 26850 9676
rect 26881 9673 26893 9676
rect 26927 9673 26939 9707
rect 26881 9667 26939 9673
rect 13357 9599 13415 9605
rect 14292 9608 16620 9636
rect 14292 9580 14320 9608
rect 17586 9596 17592 9648
rect 17644 9596 17650 9648
rect 17770 9596 17776 9648
rect 17828 9636 17834 9648
rect 18693 9639 18751 9645
rect 18693 9636 18705 9639
rect 17828 9608 18705 9636
rect 17828 9596 17834 9608
rect 18693 9605 18705 9608
rect 18739 9605 18751 9639
rect 18693 9599 18751 9605
rect 19426 9596 19432 9648
rect 19484 9596 19490 9648
rect 20070 9596 20076 9648
rect 20128 9636 20134 9648
rect 20349 9639 20407 9645
rect 20349 9636 20361 9639
rect 20128 9608 20361 9636
rect 20128 9596 20134 9608
rect 20349 9605 20361 9608
rect 20395 9605 20407 9639
rect 20349 9599 20407 9605
rect 24670 9596 24676 9648
rect 24728 9596 24734 9648
rect 5810 9568 5816 9580
rect 4724 9540 5816 9568
rect 3326 9460 3332 9512
rect 3384 9460 3390 9512
rect 4157 9503 4215 9509
rect 4157 9469 4169 9503
rect 4203 9500 4215 9503
rect 4246 9500 4252 9512
rect 4203 9472 4252 9500
rect 4203 9469 4215 9472
rect 4157 9463 4215 9469
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 4724 9509 4752 9540
rect 5810 9528 5816 9540
rect 5868 9528 5874 9580
rect 7374 9568 7380 9580
rect 6656 9540 6960 9568
rect 6656 9512 6684 9540
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9469 4767 9503
rect 4709 9463 4767 9469
rect 4798 9460 4804 9512
rect 4856 9460 4862 9512
rect 5074 9460 5080 9512
rect 5132 9460 5138 9512
rect 5261 9503 5319 9509
rect 5261 9469 5273 9503
rect 5307 9500 5319 9503
rect 5350 9500 5356 9512
rect 5307 9472 5356 9500
rect 5307 9469 5319 9472
rect 5261 9463 5319 9469
rect 5350 9460 5356 9472
rect 5408 9500 5414 9512
rect 5445 9503 5503 9509
rect 5445 9500 5457 9503
rect 5408 9472 5457 9500
rect 5408 9460 5414 9472
rect 5445 9469 5457 9472
rect 5491 9469 5503 9503
rect 5445 9463 5503 9469
rect 6362 9460 6368 9512
rect 6420 9460 6426 9512
rect 6457 9503 6515 9509
rect 6457 9469 6469 9503
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 3234 9392 3240 9444
rect 3292 9432 3298 9444
rect 3605 9435 3663 9441
rect 3605 9432 3617 9435
rect 3292 9404 3617 9432
rect 3292 9392 3298 9404
rect 3605 9401 3617 9404
rect 3651 9432 3663 9435
rect 3881 9435 3939 9441
rect 3881 9432 3893 9435
rect 3651 9404 3893 9432
rect 3651 9401 3663 9404
rect 3605 9395 3663 9401
rect 3881 9401 3893 9404
rect 3927 9432 3939 9435
rect 4430 9432 4436 9444
rect 3927 9404 4436 9432
rect 3927 9401 3939 9404
rect 3881 9395 3939 9401
rect 4430 9392 4436 9404
rect 4488 9392 4494 9444
rect 4982 9392 4988 9444
rect 5040 9432 5046 9444
rect 6472 9432 6500 9463
rect 6638 9460 6644 9512
rect 6696 9460 6702 9512
rect 6733 9503 6791 9509
rect 6733 9469 6745 9503
rect 6779 9469 6791 9503
rect 6733 9463 6791 9469
rect 5040 9404 6500 9432
rect 5040 9392 5046 9404
rect 6546 9392 6552 9444
rect 6604 9432 6610 9444
rect 6748 9432 6776 9463
rect 6822 9460 6828 9512
rect 6880 9460 6886 9512
rect 6604 9404 6776 9432
rect 6604 9392 6610 9404
rect 2958 9324 2964 9376
rect 3016 9364 3022 9376
rect 3421 9367 3479 9373
rect 3421 9364 3433 9367
rect 3016 9336 3433 9364
rect 3016 9324 3022 9336
rect 3421 9333 3433 9336
rect 3467 9333 3479 9367
rect 3421 9327 3479 9333
rect 4065 9367 4123 9373
rect 4065 9333 4077 9367
rect 4111 9364 4123 9367
rect 4525 9367 4583 9373
rect 4525 9364 4537 9367
rect 4111 9336 4537 9364
rect 4111 9333 4123 9336
rect 4065 9327 4123 9333
rect 4525 9333 4537 9336
rect 4571 9364 4583 9367
rect 6270 9364 6276 9376
rect 4571 9336 6276 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6840 9364 6868 9460
rect 6932 9432 6960 9540
rect 7116 9540 7380 9568
rect 7006 9460 7012 9512
rect 7064 9460 7070 9512
rect 7116 9509 7144 9540
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 8113 9571 8171 9577
rect 8113 9568 8125 9571
rect 7515 9540 8125 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 8113 9537 8125 9540
rect 8159 9537 8171 9571
rect 9674 9568 9680 9580
rect 8113 9531 8171 9537
rect 9232 9540 9680 9568
rect 7101 9503 7159 9509
rect 7101 9469 7113 9503
rect 7147 9469 7159 9503
rect 7101 9463 7159 9469
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9500 7251 9503
rect 8294 9500 8300 9512
rect 7239 9472 8300 9500
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 8386 9460 8392 9512
rect 8444 9460 8450 9512
rect 8754 9460 8760 9512
rect 8812 9500 8818 9512
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 8812 9472 8953 9500
rect 8812 9460 8818 9472
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 9122 9460 9128 9512
rect 9180 9460 9186 9512
rect 9232 9509 9260 9540
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 14274 9528 14280 9580
rect 14332 9528 14338 9580
rect 17604 9568 17632 9596
rect 17604 9540 18184 9568
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9469 9275 9503
rect 9217 9463 9275 9469
rect 9306 9460 9312 9512
rect 9364 9500 9370 9512
rect 10318 9500 10324 9512
rect 9364 9472 10324 9500
rect 9364 9460 9370 9472
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 11054 9460 11060 9512
rect 11112 9500 11118 9512
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 11112 9472 11897 9500
rect 11112 9460 11118 9472
rect 11885 9469 11897 9472
rect 11931 9500 11943 9503
rect 11977 9503 12035 9509
rect 11977 9500 11989 9503
rect 11931 9472 11989 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 11977 9469 11989 9472
rect 12023 9469 12035 9503
rect 11977 9463 12035 9469
rect 13446 9460 13452 9512
rect 13504 9500 13510 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13504 9472 13921 9500
rect 13504 9460 13510 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 16850 9460 16856 9512
rect 16908 9500 16914 9512
rect 17230 9503 17288 9509
rect 17230 9500 17242 9503
rect 16908 9472 17242 9500
rect 16908 9460 16914 9472
rect 17230 9469 17242 9472
rect 17276 9469 17288 9503
rect 17230 9463 17288 9469
rect 17497 9503 17555 9509
rect 17497 9469 17509 9503
rect 17543 9500 17555 9503
rect 17586 9500 17592 9512
rect 17543 9472 17592 9500
rect 17543 9469 17555 9472
rect 17497 9463 17555 9469
rect 17586 9460 17592 9472
rect 17644 9460 17650 9512
rect 18156 9500 18184 9540
rect 18230 9528 18236 9580
rect 18288 9528 18294 9580
rect 23661 9571 23719 9577
rect 19168 9540 20852 9568
rect 18877 9503 18935 9509
rect 18877 9500 18889 9503
rect 18156 9472 18889 9500
rect 18877 9469 18889 9472
rect 18923 9469 18935 9503
rect 18877 9463 18935 9469
rect 6932 9404 8616 9432
rect 7558 9364 7564 9376
rect 6840 9336 7564 9364
rect 7558 9324 7564 9336
rect 7616 9324 7622 9376
rect 8588 9373 8616 9404
rect 11146 9392 11152 9444
rect 11204 9432 11210 9444
rect 11618 9435 11676 9441
rect 11618 9432 11630 9435
rect 11204 9404 11630 9432
rect 11204 9392 11210 9404
rect 11618 9401 11630 9404
rect 11664 9401 11676 9435
rect 11618 9395 11676 9401
rect 12066 9392 12072 9444
rect 12124 9432 12130 9444
rect 12222 9435 12280 9441
rect 12222 9432 12234 9435
rect 12124 9404 12234 9432
rect 12124 9392 12130 9404
rect 12222 9401 12234 9404
rect 12268 9401 12280 9435
rect 15378 9432 15384 9444
rect 12222 9395 12280 9401
rect 12406 9404 15384 9432
rect 8573 9367 8631 9373
rect 8573 9333 8585 9367
rect 8619 9364 8631 9367
rect 9398 9364 9404 9376
rect 8619 9336 9404 9364
rect 8619 9333 8631 9336
rect 8573 9327 8631 9333
rect 9398 9324 9404 9336
rect 9456 9364 9462 9376
rect 12406 9364 12434 9404
rect 15378 9392 15384 9404
rect 15436 9392 15442 9444
rect 16022 9392 16028 9444
rect 16080 9392 16086 9444
rect 17862 9432 17868 9444
rect 16684 9404 17868 9432
rect 9456 9336 12434 9364
rect 9456 9324 9462 9336
rect 12526 9324 12532 9376
rect 12584 9364 12590 9376
rect 12802 9364 12808 9376
rect 12584 9336 12808 9364
rect 12584 9324 12590 9336
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 14093 9367 14151 9373
rect 14093 9333 14105 9367
rect 14139 9364 14151 9367
rect 16684 9364 16712 9404
rect 17862 9392 17868 9404
rect 17920 9392 17926 9444
rect 18892 9432 18920 9463
rect 18966 9460 18972 9512
rect 19024 9500 19030 9512
rect 19168 9509 19196 9540
rect 19904 9509 19932 9540
rect 20824 9509 20852 9540
rect 21284 9540 21680 9568
rect 19153 9503 19211 9509
rect 19153 9500 19165 9503
rect 19024 9472 19165 9500
rect 19024 9460 19030 9472
rect 19153 9469 19165 9472
rect 19199 9469 19211 9503
rect 19153 9463 19211 9469
rect 19613 9503 19671 9509
rect 19613 9469 19625 9503
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9469 19947 9503
rect 19889 9463 19947 9469
rect 20533 9503 20591 9509
rect 20533 9469 20545 9503
rect 20579 9469 20591 9503
rect 20533 9463 20591 9469
rect 20809 9503 20867 9509
rect 20809 9469 20821 9503
rect 20855 9469 20867 9503
rect 20809 9463 20867 9469
rect 19628 9432 19656 9463
rect 20548 9432 20576 9463
rect 18892 9404 20576 9432
rect 14139 9336 16712 9364
rect 14139 9333 14151 9336
rect 14093 9327 14151 9333
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 17589 9367 17647 9373
rect 17589 9364 17601 9367
rect 16816 9336 17601 9364
rect 16816 9324 16822 9336
rect 17589 9333 17601 9336
rect 17635 9333 17647 9367
rect 17589 9327 17647 9333
rect 19058 9324 19064 9376
rect 19116 9324 19122 9376
rect 19797 9367 19855 9373
rect 19797 9333 19809 9367
rect 19843 9364 19855 9367
rect 20346 9364 20352 9376
rect 19843 9336 20352 9364
rect 19843 9333 19855 9336
rect 19797 9327 19855 9333
rect 20346 9324 20352 9336
rect 20404 9324 20410 9376
rect 20548 9364 20576 9404
rect 20717 9435 20775 9441
rect 20717 9401 20729 9435
rect 20763 9432 20775 9435
rect 21284 9432 21312 9540
rect 21358 9460 21364 9512
rect 21416 9500 21422 9512
rect 21545 9503 21603 9509
rect 21545 9500 21557 9503
rect 21416 9472 21557 9500
rect 21416 9460 21422 9472
rect 21545 9469 21557 9472
rect 21591 9469 21603 9503
rect 21545 9463 21603 9469
rect 21652 9500 21680 9540
rect 23661 9537 23673 9571
rect 23707 9568 23719 9571
rect 23750 9568 23756 9580
rect 23707 9540 23756 9568
rect 23707 9537 23719 9540
rect 23661 9531 23719 9537
rect 23750 9528 23756 9540
rect 23808 9568 23814 9580
rect 25501 9571 25559 9577
rect 25501 9568 25513 9571
rect 23808 9540 25513 9568
rect 23808 9528 23814 9540
rect 25501 9537 25513 9540
rect 25547 9537 25559 9571
rect 25501 9531 25559 9537
rect 23842 9500 23848 9512
rect 21652 9472 23848 9500
rect 20763 9404 21312 9432
rect 20763 9401 20775 9404
rect 20717 9395 20775 9401
rect 20806 9364 20812 9376
rect 20548 9336 20812 9364
rect 20806 9324 20812 9336
rect 20864 9324 20870 9376
rect 20898 9324 20904 9376
rect 20956 9364 20962 9376
rect 21269 9367 21327 9373
rect 21269 9364 21281 9367
rect 20956 9336 21281 9364
rect 20956 9324 20962 9336
rect 21269 9333 21281 9336
rect 21315 9333 21327 9367
rect 21269 9327 21327 9333
rect 21450 9324 21456 9376
rect 21508 9324 21514 9376
rect 21560 9364 21588 9463
rect 21652 9441 21680 9472
rect 23842 9460 23848 9472
rect 23900 9460 23906 9512
rect 24854 9460 24860 9512
rect 24912 9460 24918 9512
rect 25133 9503 25191 9509
rect 25133 9469 25145 9503
rect 25179 9500 25191 9503
rect 25406 9500 25412 9512
rect 25179 9472 25412 9500
rect 25179 9469 25191 9472
rect 25133 9463 25191 9469
rect 21637 9435 21695 9441
rect 21637 9401 21649 9435
rect 21683 9401 21695 9435
rect 21637 9395 21695 9401
rect 21726 9392 21732 9444
rect 21784 9432 21790 9444
rect 21821 9435 21879 9441
rect 21821 9432 21833 9435
rect 21784 9404 21833 9432
rect 21784 9392 21790 9404
rect 21821 9401 21833 9404
rect 21867 9401 21879 9435
rect 21821 9395 21879 9401
rect 23198 9392 23204 9444
rect 23256 9432 23262 9444
rect 23394 9435 23452 9441
rect 23394 9432 23406 9435
rect 23256 9404 23406 9432
rect 23256 9392 23262 9404
rect 23394 9401 23406 9404
rect 23440 9401 23452 9435
rect 24118 9432 24124 9444
rect 23394 9395 23452 9401
rect 23492 9404 24124 9432
rect 22281 9367 22339 9373
rect 22281 9364 22293 9367
rect 21560 9336 22293 9364
rect 22281 9333 22293 9336
rect 22327 9364 22339 9367
rect 22922 9364 22928 9376
rect 22327 9336 22928 9364
rect 22327 9333 22339 9336
rect 22281 9327 22339 9333
rect 22922 9324 22928 9336
rect 22980 9364 22986 9376
rect 23492 9364 23520 9404
rect 24118 9392 24124 9404
rect 24176 9392 24182 9444
rect 24302 9392 24308 9444
rect 24360 9432 24366 9444
rect 25148 9432 25176 9463
rect 25406 9460 25412 9472
rect 25464 9460 25470 9512
rect 25774 9509 25780 9512
rect 25768 9500 25780 9509
rect 25735 9472 25780 9500
rect 25768 9463 25780 9472
rect 25774 9460 25780 9463
rect 25832 9460 25838 9512
rect 24360 9404 25176 9432
rect 24360 9392 24366 9404
rect 22980 9336 23520 9364
rect 22980 9324 22986 9336
rect 23750 9324 23756 9376
rect 23808 9364 23814 9376
rect 23937 9367 23995 9373
rect 23937 9364 23949 9367
rect 23808 9336 23949 9364
rect 23808 9324 23814 9336
rect 23937 9333 23949 9336
rect 23983 9333 23995 9367
rect 23937 9327 23995 9333
rect 24578 9324 24584 9376
rect 24636 9364 24642 9376
rect 25041 9367 25099 9373
rect 25041 9364 25053 9367
rect 24636 9336 25053 9364
rect 24636 9324 24642 9336
rect 25041 9333 25053 9336
rect 25087 9333 25099 9367
rect 25041 9327 25099 9333
rect 552 9274 27576 9296
rect 552 9222 7114 9274
rect 7166 9222 7178 9274
rect 7230 9222 7242 9274
rect 7294 9222 7306 9274
rect 7358 9222 7370 9274
rect 7422 9222 13830 9274
rect 13882 9222 13894 9274
rect 13946 9222 13958 9274
rect 14010 9222 14022 9274
rect 14074 9222 14086 9274
rect 14138 9222 20546 9274
rect 20598 9222 20610 9274
rect 20662 9222 20674 9274
rect 20726 9222 20738 9274
rect 20790 9222 20802 9274
rect 20854 9222 27262 9274
rect 27314 9222 27326 9274
rect 27378 9222 27390 9274
rect 27442 9222 27454 9274
rect 27506 9222 27518 9274
rect 27570 9222 27576 9274
rect 552 9200 27576 9222
rect 6273 9163 6331 9169
rect 6273 9129 6285 9163
rect 6319 9160 6331 9163
rect 7006 9160 7012 9172
rect 6319 9132 7012 9160
rect 6319 9129 6331 9132
rect 6273 9123 6331 9129
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 11057 9163 11115 9169
rect 7116 9132 9168 9160
rect 6362 9052 6368 9104
rect 6420 9092 6426 9104
rect 6914 9092 6920 9104
rect 6420 9064 6920 9092
rect 6420 9052 6426 9064
rect 2124 9027 2182 9033
rect 2124 8993 2136 9027
rect 2170 9024 2182 9027
rect 3602 9024 3608 9036
rect 2170 8996 3608 9024
rect 2170 8993 2182 8996
rect 2124 8987 2182 8993
rect 3602 8984 3608 8996
rect 3660 8984 3666 9036
rect 6472 9033 6500 9064
rect 6914 9052 6920 9064
rect 6972 9092 6978 9104
rect 7116 9092 7144 9132
rect 8941 9095 8999 9101
rect 8941 9092 8953 9095
rect 6972 9064 7144 9092
rect 7392 9064 8953 9092
rect 6972 9052 6978 9064
rect 6457 9027 6515 9033
rect 6457 8993 6469 9027
rect 6503 8993 6515 9027
rect 6457 8987 6515 8993
rect 6549 9027 6607 9033
rect 6549 8993 6561 9027
rect 6595 8993 6607 9027
rect 6549 8987 6607 8993
rect 1578 8916 1584 8968
rect 1636 8956 1642 8968
rect 1857 8959 1915 8965
rect 1857 8956 1869 8959
rect 1636 8928 1869 8956
rect 1636 8916 1642 8928
rect 1857 8925 1869 8928
rect 1903 8925 1915 8959
rect 3513 8959 3571 8965
rect 3513 8956 3525 8959
rect 1857 8919 1915 8925
rect 3252 8928 3525 8956
rect 3252 8897 3280 8928
rect 3513 8925 3525 8928
rect 3559 8956 3571 8959
rect 4890 8956 4896 8968
rect 3559 8928 4896 8956
rect 3559 8925 3571 8928
rect 3513 8919 3571 8925
rect 4890 8916 4896 8928
rect 4948 8956 4954 8968
rect 6564 8956 6592 8987
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 6733 9027 6791 9033
rect 6733 9024 6745 9027
rect 6696 8996 6745 9024
rect 6696 8984 6702 8996
rect 6733 8993 6745 8996
rect 6779 8993 6791 9027
rect 6733 8987 6791 8993
rect 6822 8984 6828 9036
rect 6880 8984 6886 9036
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 8993 7251 9027
rect 7193 8987 7251 8993
rect 4948 8928 6592 8956
rect 7208 8956 7236 8987
rect 7282 8984 7288 9036
rect 7340 8984 7346 9036
rect 7392 9033 7420 9064
rect 8941 9061 8953 9064
rect 8987 9061 8999 9095
rect 8941 9055 8999 9061
rect 9140 9036 9168 9132
rect 11057 9129 11069 9163
rect 11103 9160 11115 9163
rect 11146 9160 11152 9172
rect 11103 9132 11152 9160
rect 11103 9129 11115 9132
rect 11057 9123 11115 9129
rect 11146 9120 11152 9132
rect 11204 9120 11210 9172
rect 12066 9120 12072 9172
rect 12124 9120 12130 9172
rect 12710 9160 12716 9172
rect 12176 9132 12716 9160
rect 7377 9027 7435 9033
rect 7377 8993 7389 9027
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 7558 8984 7564 9036
rect 7616 8984 7622 9036
rect 8202 8984 8208 9036
rect 8260 8984 8266 9036
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 8352 8996 8397 9024
rect 8352 8984 8358 8996
rect 8478 8984 8484 9036
rect 8536 8984 8542 9036
rect 8573 9027 8631 9033
rect 8573 8993 8585 9027
rect 8619 8993 8631 9027
rect 8573 8987 8631 8993
rect 7650 8956 7656 8968
rect 7208 8928 7656 8956
rect 4948 8916 4954 8928
rect 7650 8916 7656 8928
rect 7708 8956 7714 8968
rect 8588 8956 8616 8987
rect 8662 8984 8668 9036
rect 8720 9033 8726 9036
rect 8720 9024 8728 9033
rect 8720 8996 8765 9024
rect 8720 8987 8728 8996
rect 8720 8984 8726 8987
rect 9122 8984 9128 9036
rect 9180 8984 9186 9036
rect 9217 9027 9275 9033
rect 9217 8993 9229 9027
rect 9263 8993 9275 9027
rect 9217 8987 9275 8993
rect 9232 8956 9260 8987
rect 9398 8984 9404 9036
rect 9456 8984 9462 9036
rect 9490 8984 9496 9036
rect 9548 8984 9554 9036
rect 11701 9027 11759 9033
rect 11701 8993 11713 9027
rect 11747 9024 11759 9027
rect 12176 9024 12204 9132
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 15013 9163 15071 9169
rect 15013 9129 15025 9163
rect 15059 9160 15071 9163
rect 15749 9163 15807 9169
rect 15749 9160 15761 9163
rect 15059 9132 15761 9160
rect 15059 9129 15071 9132
rect 15013 9123 15071 9129
rect 15749 9129 15761 9132
rect 15795 9160 15807 9163
rect 16758 9160 16764 9172
rect 15795 9132 16764 9160
rect 15795 9129 15807 9132
rect 15749 9123 15807 9129
rect 16758 9120 16764 9132
rect 16816 9120 16822 9172
rect 17497 9163 17555 9169
rect 17497 9129 17509 9163
rect 17543 9160 17555 9163
rect 18230 9160 18236 9172
rect 17543 9132 18236 9160
rect 17543 9129 17555 9132
rect 17497 9123 17555 9129
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 19058 9120 19064 9172
rect 19116 9160 19122 9172
rect 19521 9163 19579 9169
rect 19116 9132 19472 9160
rect 19116 9120 19122 9132
rect 13262 9092 13268 9104
rect 12360 9064 13268 9092
rect 11747 8996 12204 9024
rect 11747 8993 11759 8996
rect 11701 8987 11759 8993
rect 12250 8984 12256 9036
rect 12308 9024 12314 9036
rect 12360 9033 12388 9064
rect 13262 9052 13268 9064
rect 13320 9052 13326 9104
rect 16574 9092 16580 9104
rect 14936 9064 15700 9092
rect 12345 9027 12403 9033
rect 12345 9024 12357 9027
rect 12308 8996 12357 9024
rect 12308 8984 12314 8996
rect 12345 8993 12357 8996
rect 12391 8993 12403 9027
rect 12345 8987 12403 8993
rect 12434 8984 12440 9036
rect 12492 8984 12498 9036
rect 12550 9027 12608 9033
rect 12550 8993 12562 9027
rect 12596 9024 12608 9027
rect 12713 9027 12771 9033
rect 12596 8996 12664 9024
rect 12596 8993 12608 8996
rect 12550 8987 12608 8993
rect 7708 8928 8616 8956
rect 8680 8928 9260 8956
rect 7708 8916 7714 8928
rect 3237 8891 3295 8897
rect 3237 8857 3249 8891
rect 3283 8857 3295 8891
rect 3237 8851 3295 8857
rect 7558 8848 7564 8900
rect 7616 8888 7622 8900
rect 8680 8888 8708 8928
rect 7616 8860 8708 8888
rect 7616 8848 7622 8860
rect 8846 8848 8852 8900
rect 8904 8848 8910 8900
rect 11330 8888 11336 8900
rect 9324 8860 11336 8888
rect 4157 8823 4215 8829
rect 4157 8789 4169 8823
rect 4203 8820 4215 8823
rect 4430 8820 4436 8832
rect 4203 8792 4436 8820
rect 4203 8789 4215 8792
rect 4157 8783 4215 8789
rect 4430 8780 4436 8792
rect 4488 8780 4494 8832
rect 6914 8780 6920 8832
rect 6972 8780 6978 8832
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 8938 8820 8944 8832
rect 8260 8792 8944 8820
rect 8260 8780 8266 8792
rect 8938 8780 8944 8792
rect 8996 8820 9002 8832
rect 9324 8820 9352 8860
rect 11330 8848 11336 8860
rect 11388 8848 11394 8900
rect 12526 8848 12532 8900
rect 12584 8888 12590 8900
rect 12636 8888 12664 8996
rect 12713 8993 12725 9027
rect 12759 9024 12771 9027
rect 12802 9024 12808 9036
rect 12759 8996 12808 9024
rect 12759 8993 12771 8996
rect 12713 8987 12771 8993
rect 12802 8984 12808 8996
rect 12860 9024 12866 9036
rect 14550 9024 14556 9036
rect 12860 8996 14556 9024
rect 12860 8984 12866 8996
rect 14550 8984 14556 8996
rect 14608 8984 14614 9036
rect 14936 9033 14964 9064
rect 15672 9036 15700 9064
rect 16132 9064 16580 9092
rect 14921 9027 14979 9033
rect 14921 8993 14933 9027
rect 14967 8993 14979 9027
rect 14921 8987 14979 8993
rect 15197 9027 15255 9033
rect 15197 8993 15209 9027
rect 15243 8993 15255 9027
rect 15197 8987 15255 8993
rect 15212 8956 15240 8987
rect 15654 8984 15660 9036
rect 15712 8984 15718 9036
rect 15930 8984 15936 9036
rect 15988 8984 15994 9036
rect 16132 9033 16160 9064
rect 16574 9052 16580 9064
rect 16632 9052 16638 9104
rect 17954 9092 17960 9104
rect 17788 9064 17960 9092
rect 17788 9033 17816 9064
rect 17954 9052 17960 9064
rect 18012 9092 18018 9104
rect 19337 9095 19395 9101
rect 19337 9092 19349 9095
rect 18012 9064 19349 9092
rect 18012 9052 18018 9064
rect 19337 9061 19349 9064
rect 19383 9061 19395 9095
rect 19444 9092 19472 9132
rect 19521 9129 19533 9163
rect 19567 9160 19579 9163
rect 20898 9160 20904 9172
rect 19567 9132 20904 9160
rect 19567 9129 19579 9132
rect 19521 9123 19579 9129
rect 20898 9120 20904 9132
rect 20956 9120 20962 9172
rect 21634 9120 21640 9172
rect 21692 9160 21698 9172
rect 21821 9163 21879 9169
rect 21821 9160 21833 9163
rect 21692 9132 21833 9160
rect 21692 9120 21698 9132
rect 21821 9129 21833 9132
rect 21867 9129 21879 9163
rect 21821 9123 21879 9129
rect 23198 9120 23204 9172
rect 23256 9120 23262 9172
rect 23842 9120 23848 9172
rect 23900 9160 23906 9172
rect 26237 9163 26295 9169
rect 26237 9160 26249 9163
rect 23900 9132 26249 9160
rect 23900 9120 23906 9132
rect 26237 9129 26249 9132
rect 26283 9129 26295 9163
rect 26237 9123 26295 9129
rect 26878 9120 26884 9172
rect 26936 9120 26942 9172
rect 19889 9095 19947 9101
rect 19889 9092 19901 9095
rect 19444 9064 19901 9092
rect 19337 9055 19395 9061
rect 19889 9061 19901 9064
rect 19935 9092 19947 9095
rect 20070 9092 20076 9104
rect 19935 9064 20076 9092
rect 19935 9061 19947 9064
rect 19889 9055 19947 9061
rect 20070 9052 20076 9064
rect 20128 9052 20134 9104
rect 23474 9052 23480 9104
rect 23532 9092 23538 9104
rect 25314 9092 25320 9104
rect 23532 9064 23980 9092
rect 23532 9052 23538 9064
rect 16117 9027 16175 9033
rect 16117 8993 16129 9027
rect 16163 8993 16175 9027
rect 16373 9027 16431 9033
rect 16373 9024 16385 9027
rect 16117 8987 16175 8993
rect 16224 8996 16385 9024
rect 16224 8956 16252 8996
rect 16373 8993 16385 8996
rect 16419 8993 16431 9027
rect 16373 8987 16431 8993
rect 17773 9027 17831 9033
rect 17773 8993 17785 9027
rect 17819 8993 17831 9027
rect 17773 8987 17831 8993
rect 17865 9027 17923 9033
rect 17865 8993 17877 9027
rect 17911 9024 17923 9027
rect 18230 9024 18236 9036
rect 17911 8996 18236 9024
rect 17911 8993 17923 8996
rect 17865 8987 17923 8993
rect 18230 8984 18236 8996
rect 18288 8984 18294 9036
rect 19518 8984 19524 9036
rect 19576 9024 19582 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 19576 8996 19625 9024
rect 19576 8984 19582 8996
rect 19613 8993 19625 8996
rect 19659 8993 19671 9027
rect 19613 8987 19671 8993
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 8993 19763 9027
rect 19705 8987 19763 8993
rect 15212 8928 15884 8956
rect 12584 8860 12664 8888
rect 15197 8891 15255 8897
rect 12584 8848 12590 8860
rect 15197 8857 15209 8891
rect 15243 8888 15255 8891
rect 15746 8888 15752 8900
rect 15243 8860 15752 8888
rect 15243 8857 15255 8860
rect 15197 8851 15255 8857
rect 15746 8848 15752 8860
rect 15804 8848 15810 8900
rect 8996 8792 9352 8820
rect 15856 8820 15884 8928
rect 15948 8928 16252 8956
rect 15948 8897 15976 8928
rect 17126 8916 17132 8968
rect 17184 8956 17190 8968
rect 17589 8959 17647 8965
rect 17589 8956 17601 8959
rect 17184 8928 17601 8956
rect 17184 8916 17190 8928
rect 17589 8925 17601 8928
rect 17635 8925 17647 8959
rect 17589 8919 17647 8925
rect 17678 8916 17684 8968
rect 17736 8956 17742 8968
rect 17957 8959 18015 8965
rect 17957 8956 17969 8959
rect 17736 8928 17969 8956
rect 17736 8916 17742 8928
rect 17957 8925 17969 8928
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 18046 8916 18052 8968
rect 18104 8956 18110 8968
rect 18690 8956 18696 8968
rect 18104 8928 18696 8956
rect 18104 8916 18110 8928
rect 18690 8916 18696 8928
rect 18748 8916 18754 8968
rect 19720 8956 19748 8987
rect 21450 8984 21456 9036
rect 21508 9024 21514 9036
rect 21508 8996 22094 9024
rect 21508 8984 21514 8996
rect 19794 8956 19800 8968
rect 19720 8928 19800 8956
rect 19794 8916 19800 8928
rect 19852 8956 19858 8968
rect 21634 8956 21640 8968
rect 19852 8928 21640 8956
rect 19852 8916 19858 8928
rect 21634 8916 21640 8928
rect 21692 8916 21698 8968
rect 22066 8956 22094 8996
rect 23382 8984 23388 9036
rect 23440 9024 23446 9036
rect 23569 9027 23627 9033
rect 23569 9024 23581 9027
rect 23440 8996 23581 9024
rect 23440 8984 23446 8996
rect 23569 8993 23581 8996
rect 23615 8993 23627 9027
rect 23569 8987 23627 8993
rect 23658 8984 23664 9036
rect 23716 8984 23722 9036
rect 23952 9033 23980 9064
rect 24872 9064 25320 9092
rect 23753 9027 23811 9033
rect 23753 8993 23765 9027
rect 23799 8993 23811 9027
rect 23753 8987 23811 8993
rect 23937 9027 23995 9033
rect 23937 8993 23949 9027
rect 23983 8993 23995 9027
rect 23937 8987 23995 8993
rect 22465 8959 22523 8965
rect 22465 8956 22477 8959
rect 22066 8928 22477 8956
rect 22465 8925 22477 8928
rect 22511 8925 22523 8959
rect 22465 8919 22523 8925
rect 22649 8959 22707 8965
rect 22649 8925 22661 8959
rect 22695 8956 22707 8959
rect 23293 8959 23351 8965
rect 23293 8956 23305 8959
rect 22695 8928 23305 8956
rect 22695 8925 22707 8928
rect 22649 8919 22707 8925
rect 23293 8925 23305 8928
rect 23339 8925 23351 8959
rect 23768 8956 23796 8987
rect 24118 8984 24124 9036
rect 24176 9024 24182 9036
rect 24872 9033 24900 9064
rect 25314 9052 25320 9064
rect 25372 9052 25378 9104
rect 25866 9052 25872 9104
rect 25924 9092 25930 9104
rect 26513 9095 26571 9101
rect 26513 9092 26525 9095
rect 25924 9064 26525 9092
rect 25924 9052 25930 9064
rect 26513 9061 26525 9064
rect 26559 9061 26571 9095
rect 26513 9055 26571 9061
rect 24489 9027 24547 9033
rect 24489 9024 24501 9027
rect 24176 8996 24501 9024
rect 24176 8984 24182 8996
rect 24489 8993 24501 8996
rect 24535 8993 24547 9027
rect 24489 8987 24547 8993
rect 24857 9027 24915 9033
rect 24857 8993 24869 9027
rect 24903 8993 24915 9027
rect 24857 8987 24915 8993
rect 24946 8984 24952 9036
rect 25004 9024 25010 9036
rect 25113 9027 25171 9033
rect 25113 9024 25125 9027
rect 25004 8996 25125 9024
rect 25004 8984 25010 8996
rect 25113 8993 25125 8996
rect 25159 8993 25171 9027
rect 25113 8987 25171 8993
rect 25406 8984 25412 9036
rect 25464 9024 25470 9036
rect 26421 9027 26479 9033
rect 26421 9024 26433 9027
rect 25464 8996 26433 9024
rect 25464 8984 25470 8996
rect 26421 8993 26433 8996
rect 26467 8993 26479 9027
rect 26421 8987 26479 8993
rect 26697 9027 26755 9033
rect 26697 8993 26709 9027
rect 26743 8993 26755 9027
rect 26697 8987 26755 8993
rect 24029 8959 24087 8965
rect 24029 8956 24041 8959
rect 23768 8928 24041 8956
rect 23293 8919 23351 8925
rect 24029 8925 24041 8928
rect 24075 8925 24087 8959
rect 24213 8959 24271 8965
rect 24213 8956 24225 8959
rect 24029 8919 24087 8925
rect 24136 8928 24225 8956
rect 15933 8891 15991 8897
rect 15933 8857 15945 8891
rect 15979 8857 15991 8891
rect 15933 8851 15991 8857
rect 17696 8820 17724 8916
rect 22480 8888 22508 8919
rect 24136 8900 24164 8928
rect 24213 8925 24225 8928
rect 24259 8925 24271 8959
rect 24213 8919 24271 8925
rect 24302 8916 24308 8968
rect 24360 8916 24366 8968
rect 24394 8916 24400 8968
rect 24452 8916 24458 8968
rect 23474 8888 23480 8900
rect 22480 8860 23480 8888
rect 23474 8848 23480 8860
rect 23532 8848 23538 8900
rect 24118 8848 24124 8900
rect 24176 8888 24182 8900
rect 24762 8888 24768 8900
rect 24176 8860 24768 8888
rect 24176 8848 24182 8860
rect 24762 8848 24768 8860
rect 24820 8848 24826 8900
rect 15856 8792 17724 8820
rect 8996 8780 9002 8792
rect 17770 8780 17776 8832
rect 17828 8820 17834 8832
rect 21266 8820 21272 8832
rect 17828 8792 21272 8820
rect 17828 8780 17834 8792
rect 21266 8780 21272 8792
rect 21324 8820 21330 8832
rect 22462 8820 22468 8832
rect 21324 8792 22468 8820
rect 21324 8780 21330 8792
rect 22462 8780 22468 8792
rect 22520 8780 22526 8832
rect 24854 8780 24860 8832
rect 24912 8820 24918 8832
rect 26712 8820 26740 8987
rect 24912 8792 26740 8820
rect 24912 8780 24918 8792
rect 552 8730 27416 8752
rect 552 8678 3756 8730
rect 3808 8678 3820 8730
rect 3872 8678 3884 8730
rect 3936 8678 3948 8730
rect 4000 8678 4012 8730
rect 4064 8678 10472 8730
rect 10524 8678 10536 8730
rect 10588 8678 10600 8730
rect 10652 8678 10664 8730
rect 10716 8678 10728 8730
rect 10780 8678 17188 8730
rect 17240 8678 17252 8730
rect 17304 8678 17316 8730
rect 17368 8678 17380 8730
rect 17432 8678 17444 8730
rect 17496 8678 23904 8730
rect 23956 8678 23968 8730
rect 24020 8678 24032 8730
rect 24084 8678 24096 8730
rect 24148 8678 24160 8730
rect 24212 8678 27416 8730
rect 552 8656 27416 8678
rect 3602 8576 3608 8628
rect 3660 8616 3666 8628
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3660 8588 3985 8616
rect 3660 8576 3666 8588
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 3973 8579 4031 8585
rect 7650 8576 7656 8628
rect 7708 8576 7714 8628
rect 8386 8576 8392 8628
rect 8444 8616 8450 8628
rect 8662 8616 8668 8628
rect 8444 8588 8668 8616
rect 8444 8576 8450 8588
rect 8662 8576 8668 8588
rect 8720 8616 8726 8628
rect 11790 8616 11796 8628
rect 8720 8588 11796 8616
rect 8720 8576 8726 8588
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 11977 8619 12035 8625
rect 11977 8585 11989 8619
rect 12023 8616 12035 8619
rect 12526 8616 12532 8628
rect 12023 8588 12532 8616
rect 12023 8585 12035 8588
rect 11977 8579 12035 8585
rect 12526 8576 12532 8588
rect 12584 8576 12590 8628
rect 15930 8576 15936 8628
rect 15988 8616 15994 8628
rect 16577 8619 16635 8625
rect 16577 8616 16589 8619
rect 15988 8588 16589 8616
rect 15988 8576 15994 8588
rect 16577 8585 16589 8588
rect 16623 8585 16635 8619
rect 16577 8579 16635 8585
rect 18325 8619 18383 8625
rect 18325 8585 18337 8619
rect 18371 8616 18383 8619
rect 18371 8588 19932 8616
rect 18371 8585 18383 8588
rect 18325 8579 18383 8585
rect 3326 8508 3332 8560
rect 3384 8548 3390 8560
rect 3878 8548 3884 8560
rect 3384 8520 3884 8548
rect 3384 8508 3390 8520
rect 3878 8508 3884 8520
rect 3936 8548 3942 8560
rect 4525 8551 4583 8557
rect 4525 8548 4537 8551
rect 3936 8520 4537 8548
rect 3936 8508 3942 8520
rect 4525 8517 4537 8520
rect 4571 8517 4583 8551
rect 4525 8511 4583 8517
rect 6825 8551 6883 8557
rect 6825 8517 6837 8551
rect 6871 8548 6883 8551
rect 6871 8520 7052 8548
rect 6871 8517 6883 8520
rect 6825 8511 6883 8517
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 2832 8452 4353 8480
rect 2832 8440 2838 8452
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4430 8440 4436 8492
rect 4488 8440 4494 8492
rect 4890 8440 4896 8492
rect 4948 8440 4954 8492
rect 7024 8489 7052 8520
rect 8570 8508 8576 8560
rect 8628 8548 8634 8560
rect 10689 8551 10747 8557
rect 8628 8520 10180 8548
rect 8628 8508 8634 8520
rect 7009 8483 7067 8489
rect 7009 8449 7021 8483
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 9674 8480 9680 8492
rect 8536 8452 9680 8480
rect 8536 8440 8542 8452
rect 1578 8372 1584 8424
rect 1636 8372 1642 8424
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8381 3939 8415
rect 3881 8375 3939 8381
rect 1848 8347 1906 8353
rect 1848 8313 1860 8347
rect 1894 8344 1906 8347
rect 2590 8344 2596 8356
rect 1894 8316 2596 8344
rect 1894 8313 1906 8316
rect 1848 8307 1906 8313
rect 2590 8304 2596 8316
rect 2648 8304 2654 8356
rect 3142 8344 3148 8356
rect 2976 8316 3148 8344
rect 2976 8285 3004 8316
rect 3142 8304 3148 8316
rect 3200 8344 3206 8356
rect 3896 8344 3924 8375
rect 4154 8372 4160 8424
rect 4212 8372 4218 8424
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8412 4767 8415
rect 4982 8412 4988 8424
rect 4755 8384 4988 8412
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 4724 8344 4752 8375
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 5442 8372 5448 8424
rect 5500 8372 5506 8424
rect 5712 8415 5770 8421
rect 5712 8381 5724 8415
rect 5758 8412 5770 8415
rect 6914 8412 6920 8424
rect 5758 8384 6920 8412
rect 5758 8381 5770 8384
rect 5712 8375 5770 8381
rect 6914 8372 6920 8384
rect 6972 8372 6978 8424
rect 8754 8372 8760 8424
rect 8812 8372 8818 8424
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 9048 8421 9076 8452
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8904 8384 8953 8412
rect 8904 8372 8910 8384
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8381 9183 8415
rect 9125 8375 9183 8381
rect 3200 8316 4752 8344
rect 3200 8304 3206 8316
rect 8662 8304 8668 8356
rect 8720 8344 8726 8356
rect 9140 8344 9168 8375
rect 8720 8316 9168 8344
rect 8720 8304 8726 8316
rect 2961 8279 3019 8285
rect 2961 8245 2973 8279
rect 3007 8245 3019 8279
rect 2961 8239 3019 8245
rect 3237 8279 3295 8285
rect 3237 8245 3249 8279
rect 3283 8276 3295 8279
rect 3510 8276 3516 8288
rect 3283 8248 3516 8276
rect 3283 8245 3295 8248
rect 3237 8239 3295 8245
rect 3510 8236 3516 8248
rect 3568 8236 3574 8288
rect 6086 8236 6092 8288
rect 6144 8276 6150 8288
rect 7282 8276 7288 8288
rect 6144 8248 7288 8276
rect 6144 8236 6150 8248
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 9398 8236 9404 8288
rect 9456 8236 9462 8288
rect 10152 8276 10180 8520
rect 10689 8517 10701 8551
rect 10735 8548 10747 8551
rect 12158 8548 12164 8560
rect 10735 8520 12164 8548
rect 10735 8517 10747 8520
rect 10689 8511 10747 8517
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 15654 8508 15660 8560
rect 15712 8548 15718 8560
rect 16669 8551 16727 8557
rect 16669 8548 16681 8551
rect 15712 8520 16681 8548
rect 15712 8508 15718 8520
rect 16669 8517 16681 8520
rect 16715 8548 16727 8551
rect 17954 8548 17960 8560
rect 16715 8520 17960 8548
rect 16715 8517 16727 8520
rect 16669 8511 16727 8517
rect 17954 8508 17960 8520
rect 18012 8508 18018 8560
rect 19904 8548 19932 8588
rect 20070 8576 20076 8628
rect 20128 8576 20134 8628
rect 20165 8619 20223 8625
rect 20165 8585 20177 8619
rect 20211 8616 20223 8619
rect 20346 8616 20352 8628
rect 20211 8588 20352 8616
rect 20211 8585 20223 8588
rect 20165 8579 20223 8585
rect 20346 8576 20352 8588
rect 20404 8616 20410 8628
rect 21726 8616 21732 8628
rect 20404 8588 21732 8616
rect 20404 8576 20410 8588
rect 21726 8576 21732 8588
rect 21784 8576 21790 8628
rect 22281 8619 22339 8625
rect 22281 8585 22293 8619
rect 22327 8616 22339 8619
rect 22554 8616 22560 8628
rect 22327 8588 22560 8616
rect 22327 8585 22339 8588
rect 22281 8579 22339 8585
rect 22554 8576 22560 8588
rect 22612 8576 22618 8628
rect 23569 8619 23627 8625
rect 23569 8585 23581 8619
rect 23615 8616 23627 8619
rect 23658 8616 23664 8628
rect 23615 8588 23664 8616
rect 23615 8585 23627 8588
rect 23569 8579 23627 8585
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 23937 8619 23995 8625
rect 23937 8585 23949 8619
rect 23983 8585 23995 8619
rect 23937 8579 23995 8585
rect 19904 8520 20208 8548
rect 20180 8492 20208 8520
rect 23382 8508 23388 8560
rect 23440 8548 23446 8560
rect 23842 8548 23848 8560
rect 23440 8520 23848 8548
rect 23440 8508 23446 8520
rect 23842 8508 23848 8520
rect 23900 8548 23906 8560
rect 23952 8548 23980 8579
rect 24486 8576 24492 8628
rect 24544 8576 24550 8628
rect 25133 8619 25191 8625
rect 25133 8585 25145 8619
rect 25179 8616 25191 8619
rect 25409 8619 25467 8625
rect 25409 8616 25421 8619
rect 25179 8588 25421 8616
rect 25179 8585 25191 8588
rect 25133 8579 25191 8585
rect 25409 8585 25421 8588
rect 25455 8585 25467 8619
rect 25409 8579 25467 8585
rect 23900 8520 24624 8548
rect 23900 8508 23906 8520
rect 10226 8440 10232 8492
rect 10284 8480 10290 8492
rect 10778 8480 10784 8492
rect 10284 8452 10784 8480
rect 10284 8440 10290 8452
rect 10778 8440 10784 8452
rect 10836 8480 10842 8492
rect 12710 8480 12716 8492
rect 10836 8452 11192 8480
rect 10836 8440 10842 8452
rect 10873 8415 10931 8421
rect 10873 8381 10885 8415
rect 10919 8381 10931 8415
rect 10873 8375 10931 8381
rect 10888 8344 10916 8375
rect 10962 8372 10968 8424
rect 11020 8372 11026 8424
rect 11164 8421 11192 8452
rect 11716 8452 12716 8480
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 11238 8372 11244 8424
rect 11296 8372 11302 8424
rect 11330 8372 11336 8424
rect 11388 8372 11394 8424
rect 11481 8415 11539 8421
rect 11481 8381 11493 8415
rect 11527 8412 11539 8415
rect 11716 8412 11744 8452
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 13354 8440 13360 8492
rect 13412 8480 13418 8492
rect 13412 8452 13860 8480
rect 13412 8440 13418 8452
rect 11527 8384 11744 8412
rect 11527 8381 11539 8384
rect 11481 8375 11539 8381
rect 11790 8372 11796 8424
rect 11848 8421 11854 8424
rect 11848 8412 11856 8421
rect 11848 8384 11893 8412
rect 11848 8375 11856 8384
rect 11848 8372 11854 8375
rect 12158 8372 12164 8424
rect 12216 8412 12222 8424
rect 12342 8412 12348 8424
rect 12216 8384 12348 8412
rect 12216 8372 12222 8384
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 12894 8372 12900 8424
rect 12952 8372 12958 8424
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8381 13599 8415
rect 13541 8375 13599 8381
rect 11054 8344 11060 8356
rect 10888 8316 11060 8344
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 11606 8344 11612 8356
rect 11256 8316 11612 8344
rect 11256 8276 11284 8316
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 11701 8347 11759 8353
rect 11701 8313 11713 8347
rect 11747 8344 11759 8347
rect 11974 8344 11980 8356
rect 11747 8316 11980 8344
rect 11747 8313 11759 8316
rect 11701 8307 11759 8313
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 12618 8304 12624 8356
rect 12676 8344 12682 8356
rect 13556 8344 13584 8375
rect 13630 8372 13636 8424
rect 13688 8412 13694 8424
rect 13832 8421 13860 8452
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 16482 8480 16488 8492
rect 16356 8452 16488 8480
rect 16356 8440 16362 8452
rect 16482 8440 16488 8452
rect 16540 8480 16546 8492
rect 16540 8452 17540 8480
rect 16540 8440 16546 8452
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 13688 8384 13737 8412
rect 13688 8372 13694 8384
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 13817 8415 13875 8421
rect 13817 8381 13829 8415
rect 13863 8381 13875 8415
rect 13817 8375 13875 8381
rect 13909 8415 13967 8421
rect 13909 8381 13921 8415
rect 13955 8412 13967 8415
rect 14366 8412 14372 8424
rect 13955 8384 14372 8412
rect 13955 8381 13967 8384
rect 13909 8375 13967 8381
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 16393 8415 16451 8421
rect 16393 8381 16405 8415
rect 16439 8381 16451 8415
rect 16393 8375 16451 8381
rect 12676 8316 13584 8344
rect 16408 8344 16436 8375
rect 16758 8372 16764 8424
rect 16816 8372 16822 8424
rect 17512 8412 17540 8452
rect 17586 8440 17592 8492
rect 17644 8480 17650 8492
rect 18693 8483 18751 8489
rect 18693 8480 18705 8483
rect 17644 8452 18705 8480
rect 17644 8440 17650 8452
rect 18693 8449 18705 8452
rect 18739 8449 18751 8483
rect 18693 8443 18751 8449
rect 20162 8440 20168 8492
rect 20220 8440 20226 8492
rect 21726 8440 21732 8492
rect 21784 8440 21790 8492
rect 22373 8491 22431 8497
rect 22373 8457 22385 8491
rect 22419 8480 22431 8491
rect 22462 8480 22468 8492
rect 22419 8457 22468 8480
rect 22373 8452 22468 8457
rect 22373 8451 22431 8452
rect 22462 8440 22468 8452
rect 22520 8440 22526 8492
rect 23750 8440 23756 8492
rect 23808 8480 23814 8492
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 23808 8452 23949 8480
rect 23808 8440 23814 8452
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 24596 8480 24624 8520
rect 24670 8508 24676 8560
rect 24728 8508 24734 8560
rect 25593 8551 25651 8557
rect 25593 8517 25605 8551
rect 25639 8517 25651 8551
rect 25593 8511 25651 8517
rect 25406 8480 25412 8492
rect 24596 8452 25412 8480
rect 23937 8443 23995 8449
rect 25406 8440 25412 8452
rect 25464 8440 25470 8492
rect 17770 8412 17776 8424
rect 17512 8384 17776 8412
rect 17770 8372 17776 8384
rect 17828 8372 17834 8424
rect 21545 8415 21603 8421
rect 21545 8381 21557 8415
rect 21591 8412 21603 8415
rect 21818 8412 21824 8424
rect 21591 8384 21824 8412
rect 21591 8381 21603 8384
rect 21545 8375 21603 8381
rect 21818 8372 21824 8384
rect 21876 8372 21882 8424
rect 22557 8415 22615 8421
rect 22557 8381 22569 8415
rect 22603 8381 22615 8415
rect 22557 8375 22615 8381
rect 16482 8344 16488 8356
rect 16408 8316 16488 8344
rect 12676 8304 12682 8316
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 18782 8304 18788 8356
rect 18840 8344 18846 8356
rect 18938 8347 18996 8353
rect 18938 8344 18950 8347
rect 18840 8316 18950 8344
rect 18840 8304 18846 8316
rect 18938 8313 18950 8316
rect 18984 8313 18996 8347
rect 18938 8307 18996 8313
rect 21082 8304 21088 8356
rect 21140 8344 21146 8356
rect 21278 8347 21336 8353
rect 21278 8344 21290 8347
rect 21140 8316 21290 8344
rect 21140 8304 21146 8316
rect 21278 8313 21290 8316
rect 21324 8313 21336 8347
rect 21278 8307 21336 8313
rect 22002 8304 22008 8356
rect 22060 8344 22066 8356
rect 22060 8316 22324 8344
rect 22060 8304 22066 8316
rect 10152 8248 11284 8276
rect 11330 8236 11336 8288
rect 11388 8276 11394 8288
rect 12066 8276 12072 8288
rect 11388 8248 12072 8276
rect 11388 8236 11394 8248
rect 12066 8236 12072 8248
rect 12124 8236 12130 8288
rect 12342 8236 12348 8288
rect 12400 8236 12406 8288
rect 14182 8236 14188 8288
rect 14240 8236 14246 8288
rect 14826 8236 14832 8288
rect 14884 8276 14890 8288
rect 15749 8279 15807 8285
rect 15749 8276 15761 8279
rect 14884 8248 15761 8276
rect 14884 8236 14890 8248
rect 15749 8245 15761 8248
rect 15795 8245 15807 8279
rect 15749 8239 15807 8245
rect 18322 8236 18328 8288
rect 18380 8236 18386 8288
rect 18509 8279 18567 8285
rect 18509 8245 18521 8279
rect 18555 8276 18567 8279
rect 18598 8276 18604 8288
rect 18555 8248 18604 8276
rect 18555 8245 18567 8248
rect 18509 8239 18567 8245
rect 18598 8236 18604 8248
rect 18656 8236 18662 8288
rect 19518 8236 19524 8288
rect 19576 8276 19582 8288
rect 21358 8276 21364 8288
rect 19576 8248 21364 8276
rect 19576 8236 19582 8248
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 22296 8276 22324 8316
rect 22462 8304 22468 8356
rect 22520 8344 22526 8356
rect 22572 8344 22600 8375
rect 22646 8372 22652 8424
rect 22704 8372 22710 8424
rect 23017 8415 23075 8421
rect 23017 8381 23029 8415
rect 23063 8412 23075 8415
rect 23474 8412 23480 8424
rect 23063 8384 23480 8412
rect 23063 8381 23075 8384
rect 23017 8375 23075 8381
rect 23474 8372 23480 8384
rect 23532 8412 23538 8424
rect 23845 8415 23903 8421
rect 23845 8412 23857 8415
rect 23532 8384 23857 8412
rect 23532 8372 23538 8384
rect 23845 8381 23857 8384
rect 23891 8381 23903 8415
rect 24949 8415 25007 8421
rect 23845 8375 23903 8381
rect 24228 8384 24424 8412
rect 22520 8316 22600 8344
rect 22520 8304 22526 8316
rect 22373 8279 22431 8285
rect 22373 8276 22385 8279
rect 22296 8248 22385 8276
rect 22373 8245 22385 8248
rect 22419 8245 22431 8279
rect 22373 8239 22431 8245
rect 23382 8236 23388 8288
rect 23440 8276 23446 8288
rect 24228 8285 24256 8384
rect 24305 8347 24363 8353
rect 24305 8313 24317 8347
rect 24351 8313 24363 8347
rect 24396 8344 24424 8384
rect 24949 8381 24961 8415
rect 24995 8412 25007 8415
rect 25608 8412 25636 8511
rect 25685 8415 25743 8421
rect 25685 8412 25697 8415
rect 24995 8384 25544 8412
rect 25608 8384 25697 8412
rect 24995 8381 25007 8384
rect 24949 8375 25007 8381
rect 24505 8347 24563 8353
rect 24505 8344 24517 8347
rect 24396 8316 24517 8344
rect 24305 8307 24363 8313
rect 24505 8313 24517 8316
rect 24551 8313 24563 8347
rect 24505 8307 24563 8313
rect 24596 8316 24716 8344
rect 24213 8279 24271 8285
rect 24213 8276 24225 8279
rect 23440 8248 24225 8276
rect 23440 8236 23446 8248
rect 24213 8245 24225 8248
rect 24259 8245 24271 8279
rect 24325 8276 24353 8307
rect 24596 8276 24624 8316
rect 24325 8248 24624 8276
rect 24688 8276 24716 8316
rect 24762 8304 24768 8356
rect 24820 8304 24826 8356
rect 24854 8304 24860 8356
rect 24912 8344 24918 8356
rect 25225 8347 25283 8353
rect 25225 8344 25237 8347
rect 24912 8316 25237 8344
rect 24912 8304 24918 8316
rect 25225 8313 25237 8316
rect 25271 8313 25283 8347
rect 25225 8307 25283 8313
rect 25406 8304 25412 8356
rect 25464 8353 25470 8356
rect 25464 8347 25483 8353
rect 25471 8313 25483 8347
rect 25516 8344 25544 8384
rect 25685 8381 25697 8384
rect 25731 8381 25743 8415
rect 25685 8375 25743 8381
rect 25590 8344 25596 8356
rect 25516 8316 25596 8344
rect 25464 8307 25483 8313
rect 25464 8304 25470 8307
rect 25590 8304 25596 8316
rect 25648 8344 25654 8356
rect 26878 8344 26884 8356
rect 25648 8316 26884 8344
rect 25648 8304 25654 8316
rect 26878 8304 26884 8316
rect 26936 8304 26942 8356
rect 24872 8276 24900 8304
rect 24688 8248 24900 8276
rect 24213 8239 24271 8245
rect 25774 8236 25780 8288
rect 25832 8276 25838 8288
rect 25869 8279 25927 8285
rect 25869 8276 25881 8279
rect 25832 8248 25881 8276
rect 25832 8236 25838 8248
rect 25869 8245 25881 8248
rect 25915 8245 25927 8279
rect 25869 8239 25927 8245
rect 552 8186 27576 8208
rect 552 8134 7114 8186
rect 7166 8134 7178 8186
rect 7230 8134 7242 8186
rect 7294 8134 7306 8186
rect 7358 8134 7370 8186
rect 7422 8134 13830 8186
rect 13882 8134 13894 8186
rect 13946 8134 13958 8186
rect 14010 8134 14022 8186
rect 14074 8134 14086 8186
rect 14138 8134 20546 8186
rect 20598 8134 20610 8186
rect 20662 8134 20674 8186
rect 20726 8134 20738 8186
rect 20790 8134 20802 8186
rect 20854 8134 27262 8186
rect 27314 8134 27326 8186
rect 27378 8134 27390 8186
rect 27442 8134 27454 8186
rect 27506 8134 27518 8186
rect 27570 8134 27576 8186
rect 552 8112 27576 8134
rect 2590 8032 2596 8084
rect 2648 8032 2654 8084
rect 2774 8032 2780 8084
rect 2832 8032 2838 8084
rect 8754 8032 8760 8084
rect 8812 8072 8818 8084
rect 12802 8072 12808 8084
rect 8812 8044 12808 8072
rect 8812 8032 8818 8044
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 12894 8032 12900 8084
rect 12952 8032 12958 8084
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 13679 8044 15424 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 3237 8007 3295 8013
rect 3237 8004 3249 8007
rect 2516 7976 3249 8004
rect 2516 7945 2544 7976
rect 3237 7973 3249 7976
rect 3283 7973 3295 8007
rect 3237 7967 3295 7973
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7905 2559 7939
rect 2501 7899 2559 7905
rect 2685 7939 2743 7945
rect 2685 7905 2697 7939
rect 2731 7936 2743 7939
rect 2774 7936 2780 7948
rect 2731 7908 2780 7936
rect 2731 7905 2743 7908
rect 2685 7899 2743 7905
rect 2774 7896 2780 7908
rect 2832 7896 2838 7948
rect 2958 7896 2964 7948
rect 3016 7896 3022 7948
rect 3142 7896 3148 7948
rect 3200 7896 3206 7948
rect 3510 7896 3516 7948
rect 3568 7896 3574 7948
rect 3602 7896 3608 7948
rect 3660 7936 3666 7948
rect 3878 7936 3884 7948
rect 3660 7908 3884 7936
rect 3660 7896 3666 7908
rect 3878 7896 3884 7908
rect 3936 7936 3942 7948
rect 3973 7939 4031 7945
rect 3973 7936 3985 7939
rect 3936 7908 3985 7936
rect 3936 7896 3942 7908
rect 3973 7905 3985 7908
rect 4019 7905 4031 7939
rect 3973 7899 4031 7905
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7905 4123 7939
rect 4065 7899 4123 7905
rect 2976 7800 3004 7896
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7868 3295 7871
rect 3326 7868 3332 7880
rect 3283 7840 3332 7868
rect 3283 7837 3295 7840
rect 3237 7831 3295 7837
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 4080 7868 4108 7899
rect 4246 7896 4252 7948
rect 4304 7896 4310 7948
rect 6454 7945 6460 7948
rect 6448 7899 6460 7945
rect 6454 7896 6460 7899
rect 6512 7896 6518 7948
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 8389 7939 8447 7945
rect 8389 7936 8401 7939
rect 8352 7908 8401 7936
rect 8352 7896 8358 7908
rect 8389 7905 8401 7908
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 8478 7896 8484 7948
rect 8536 7896 8542 7948
rect 8772 7945 8800 8032
rect 9674 8004 9680 8016
rect 8864 7976 9680 8004
rect 8864 7948 8892 7976
rect 9674 7964 9680 7976
rect 9732 8004 9738 8016
rect 9732 7976 11560 8004
rect 9732 7964 9738 7976
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7905 8631 7939
rect 8573 7899 8631 7905
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7905 8815 7939
rect 8757 7899 8815 7905
rect 3436 7840 4108 7868
rect 3436 7800 3464 7840
rect 5442 7828 5448 7880
rect 5500 7868 5506 7880
rect 6178 7868 6184 7880
rect 5500 7840 6184 7868
rect 5500 7828 5506 7840
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 8588 7868 8616 7899
rect 8846 7896 8852 7948
rect 8904 7896 8910 7948
rect 9116 7939 9174 7945
rect 9116 7905 9128 7939
rect 9162 7936 9174 7939
rect 9398 7936 9404 7948
rect 9162 7908 9404 7936
rect 9162 7905 9174 7908
rect 9116 7899 9174 7905
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 11532 7945 11560 7976
rect 13262 7964 13268 8016
rect 13320 7964 13326 8016
rect 13357 8007 13415 8013
rect 13357 7973 13369 8007
rect 13403 8004 13415 8007
rect 14366 8004 14372 8016
rect 13403 7976 14372 8004
rect 13403 7973 13415 7976
rect 13357 7967 13415 7973
rect 14366 7964 14372 7976
rect 14424 7964 14430 8016
rect 14550 7964 14556 8016
rect 14608 8004 14614 8016
rect 14608 7976 15240 8004
rect 14608 7964 14614 7976
rect 11790 7945 11796 7948
rect 11517 7939 11575 7945
rect 11517 7905 11529 7939
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 11784 7899 11796 7945
rect 11790 7896 11796 7899
rect 11848 7896 11854 7948
rect 12066 7896 12072 7948
rect 12124 7936 12130 7948
rect 12978 7939 13036 7945
rect 12978 7936 12990 7939
rect 12124 7908 12990 7936
rect 12124 7896 12130 7908
rect 12978 7905 12990 7908
rect 13024 7905 13036 7939
rect 12978 7899 13036 7905
rect 13082 7939 13140 7945
rect 13082 7905 13094 7939
rect 13128 7905 13140 7939
rect 13454 7939 13512 7945
rect 13454 7936 13466 7939
rect 13082 7899 13140 7905
rect 13188 7908 13466 7936
rect 8260 7840 8616 7868
rect 8260 7828 8266 7840
rect 12802 7828 12808 7880
rect 12860 7868 12866 7880
rect 13096 7868 13124 7899
rect 12860 7840 13124 7868
rect 12860 7828 12866 7840
rect 2976 7772 3464 7800
rect 3436 7744 3464 7772
rect 13188 7744 13216 7908
rect 13454 7905 13466 7908
rect 13500 7905 13512 7939
rect 13454 7899 13512 7905
rect 14467 7939 14525 7945
rect 14467 7905 14479 7939
rect 14513 7936 14525 7939
rect 14568 7936 14596 7964
rect 15212 7948 15240 7976
rect 14513 7908 14596 7936
rect 14645 7939 14703 7945
rect 14513 7905 14525 7908
rect 14467 7899 14525 7905
rect 14645 7905 14657 7939
rect 14691 7905 14703 7939
rect 14645 7899 14703 7905
rect 13722 7828 13728 7880
rect 13780 7828 13786 7880
rect 13354 7760 13360 7812
rect 13412 7800 13418 7812
rect 14660 7800 14688 7899
rect 14734 7896 14740 7948
rect 14792 7896 14798 7948
rect 14826 7896 14832 7948
rect 14884 7896 14890 7948
rect 15194 7896 15200 7948
rect 15252 7945 15258 7948
rect 15396 7945 15424 8044
rect 18782 8032 18788 8084
rect 18840 8032 18846 8084
rect 20162 8032 20168 8084
rect 20220 8072 20226 8084
rect 20530 8072 20536 8084
rect 20220 8044 20536 8072
rect 20220 8032 20226 8044
rect 20530 8032 20536 8044
rect 20588 8032 20594 8084
rect 22189 8075 22247 8081
rect 22189 8072 22201 8075
rect 20916 8044 22201 8072
rect 16574 8004 16580 8016
rect 16132 7976 16580 8004
rect 15252 7936 15261 7945
rect 15381 7939 15439 7945
rect 15252 7908 15297 7936
rect 15252 7899 15261 7908
rect 15381 7905 15393 7939
rect 15427 7905 15439 7939
rect 15381 7899 15439 7905
rect 15252 7896 15258 7899
rect 15470 7896 15476 7948
rect 15528 7896 15534 7948
rect 16132 7945 16160 7976
rect 16574 7964 16580 7976
rect 16632 8004 16638 8016
rect 17586 8004 17592 8016
rect 16632 7976 17592 8004
rect 16632 7964 16638 7976
rect 17586 7964 17592 7976
rect 17644 7964 17650 8016
rect 20806 8004 20812 8016
rect 19444 7976 20812 8004
rect 15565 7939 15623 7945
rect 15565 7905 15577 7939
rect 15611 7905 15623 7939
rect 15565 7899 15623 7905
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7905 16175 7939
rect 16373 7939 16431 7945
rect 16373 7936 16385 7939
rect 16117 7899 16175 7905
rect 16224 7908 16385 7936
rect 13412 7772 14688 7800
rect 13412 7760 13418 7772
rect 14734 7760 14740 7812
rect 14792 7800 14798 7812
rect 15488 7800 15516 7896
rect 14792 7772 15516 7800
rect 14792 7760 14798 7772
rect 3418 7692 3424 7744
rect 3476 7692 3482 7744
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 4249 7735 4307 7741
rect 4249 7732 4261 7735
rect 4212 7704 4261 7732
rect 4212 7692 4218 7704
rect 4249 7701 4261 7704
rect 4295 7701 4307 7735
rect 4249 7695 4307 7701
rect 7561 7735 7619 7741
rect 7561 7701 7573 7735
rect 7607 7732 7619 7735
rect 7742 7732 7748 7744
rect 7607 7704 7748 7732
rect 7607 7701 7619 7704
rect 7561 7695 7619 7701
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 8110 7692 8116 7744
rect 8168 7692 8174 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 10229 7735 10287 7741
rect 10229 7732 10241 7735
rect 8720 7704 10241 7732
rect 8720 7692 8726 7704
rect 10229 7701 10241 7704
rect 10275 7732 10287 7735
rect 11330 7732 11336 7744
rect 10275 7704 11336 7732
rect 10275 7701 10287 7704
rect 10229 7695 10287 7701
rect 11330 7692 11336 7704
rect 11388 7692 11394 7744
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 13170 7732 13176 7744
rect 11940 7704 13176 7732
rect 11940 7692 11946 7704
rect 13170 7692 13176 7704
rect 13228 7692 13234 7744
rect 15105 7735 15163 7741
rect 15105 7701 15117 7735
rect 15151 7732 15163 7735
rect 15378 7732 15384 7744
rect 15151 7704 15384 7732
rect 15151 7701 15163 7704
rect 15105 7695 15163 7701
rect 15378 7692 15384 7704
rect 15436 7692 15442 7744
rect 15580 7732 15608 7899
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7868 15899 7871
rect 16224 7868 16252 7908
rect 16373 7905 16385 7908
rect 16419 7905 16431 7939
rect 16373 7899 16431 7905
rect 18598 7896 18604 7948
rect 18656 7896 18662 7948
rect 19444 7945 19472 7976
rect 20806 7964 20812 7976
rect 20864 7964 20870 8016
rect 20916 8013 20944 8044
rect 22189 8041 22201 8044
rect 22235 8041 22247 8075
rect 24026 8072 24032 8084
rect 22189 8035 22247 8041
rect 23768 8044 24032 8072
rect 20901 8007 20959 8013
rect 20901 7973 20913 8007
rect 20947 7973 20959 8007
rect 20901 7967 20959 7973
rect 21008 7976 21956 8004
rect 19429 7939 19487 7945
rect 19429 7905 19441 7939
rect 19475 7905 19487 7939
rect 19429 7899 19487 7905
rect 19518 7896 19524 7948
rect 19576 7896 19582 7948
rect 19705 7939 19763 7945
rect 19705 7905 19717 7939
rect 19751 7936 19763 7939
rect 20070 7936 20076 7948
rect 19751 7908 20076 7936
rect 19751 7905 19763 7908
rect 19705 7899 19763 7905
rect 20070 7896 20076 7908
rect 20128 7896 20134 7948
rect 21008 7945 21036 7976
rect 20533 7939 20591 7945
rect 20533 7905 20545 7939
rect 20579 7905 20591 7939
rect 20533 7899 20591 7905
rect 20625 7939 20683 7945
rect 20625 7905 20637 7939
rect 20671 7936 20683 7939
rect 20993 7939 21051 7945
rect 20671 7908 20769 7936
rect 20671 7905 20683 7908
rect 20625 7899 20683 7905
rect 15887 7840 16252 7868
rect 15887 7837 15899 7840
rect 15841 7831 15899 7837
rect 18322 7828 18328 7880
rect 18380 7868 18386 7880
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 18380 7840 19257 7868
rect 18380 7828 18386 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7868 19671 7871
rect 19794 7868 19800 7880
rect 19659 7840 19800 7868
rect 19659 7837 19671 7840
rect 19613 7831 19671 7837
rect 19794 7828 19800 7840
rect 19852 7828 19858 7880
rect 20548 7868 20576 7899
rect 20548 7840 20668 7868
rect 20640 7812 20668 7840
rect 18690 7760 18696 7812
rect 18748 7800 18754 7812
rect 20622 7800 20628 7812
rect 18748 7772 20628 7800
rect 18748 7760 18754 7772
rect 20622 7760 20628 7772
rect 20680 7760 20686 7812
rect 20741 7800 20769 7908
rect 20993 7905 21005 7939
rect 21039 7905 21051 7939
rect 20993 7899 21051 7905
rect 21358 7896 21364 7948
rect 21416 7936 21422 7948
rect 21453 7939 21511 7945
rect 21453 7936 21465 7939
rect 21416 7908 21465 7936
rect 21416 7896 21422 7908
rect 21453 7905 21465 7908
rect 21499 7905 21511 7939
rect 21453 7899 21511 7905
rect 21634 7896 21640 7948
rect 21692 7896 21698 7948
rect 21729 7939 21787 7945
rect 21729 7905 21741 7939
rect 21775 7905 21787 7939
rect 21729 7899 21787 7905
rect 21821 7939 21879 7945
rect 21821 7905 21833 7939
rect 21867 7905 21879 7939
rect 21928 7936 21956 7976
rect 22002 7964 22008 8016
rect 22060 7964 22066 8016
rect 23382 8004 23388 8016
rect 22204 7976 23388 8004
rect 22204 7936 22232 7976
rect 23382 7964 23388 7976
rect 23440 7964 23446 8016
rect 21928 7908 22232 7936
rect 22281 7939 22339 7945
rect 21821 7899 21879 7905
rect 22281 7905 22293 7939
rect 22327 7936 22339 7939
rect 22554 7936 22560 7948
rect 22327 7908 22560 7936
rect 22327 7905 22339 7908
rect 22281 7899 22339 7905
rect 21082 7828 21088 7880
rect 21140 7828 21146 7880
rect 21269 7803 21327 7809
rect 21269 7800 21281 7803
rect 20741 7772 21281 7800
rect 21269 7769 21281 7772
rect 21315 7800 21327 7803
rect 21744 7800 21772 7899
rect 21836 7868 21864 7899
rect 22554 7896 22560 7908
rect 22612 7896 22618 7948
rect 23017 7939 23075 7945
rect 23017 7905 23029 7939
rect 23063 7936 23075 7939
rect 23566 7936 23572 7948
rect 23063 7908 23572 7936
rect 23063 7905 23075 7908
rect 23017 7899 23075 7905
rect 23566 7896 23572 7908
rect 23624 7936 23630 7948
rect 23661 7939 23719 7945
rect 23661 7936 23673 7939
rect 23624 7908 23673 7936
rect 23624 7896 23630 7908
rect 23661 7905 23673 7908
rect 23707 7936 23719 7939
rect 23768 7936 23796 8044
rect 24026 8032 24032 8044
rect 24084 8032 24090 8084
rect 24121 8075 24179 8081
rect 24121 8041 24133 8075
rect 24167 8072 24179 8075
rect 24486 8072 24492 8084
rect 24167 8044 24492 8072
rect 24167 8041 24179 8044
rect 24121 8035 24179 8041
rect 24486 8032 24492 8044
rect 24544 8032 24550 8084
rect 24857 8075 24915 8081
rect 24857 8041 24869 8075
rect 24903 8072 24915 8075
rect 24946 8072 24952 8084
rect 24903 8044 24952 8072
rect 24903 8041 24915 8044
rect 24857 8035 24915 8041
rect 24946 8032 24952 8044
rect 25004 8032 25010 8084
rect 24305 8007 24363 8013
rect 24305 8004 24317 8007
rect 23860 7976 24317 8004
rect 23860 7948 23888 7976
rect 24305 7973 24317 7976
rect 24351 7973 24363 8007
rect 24305 7967 24363 7973
rect 24762 7964 24768 8016
rect 24820 7964 24826 8016
rect 23707 7908 23796 7936
rect 23707 7905 23719 7908
rect 23661 7899 23719 7905
rect 23842 7896 23848 7948
rect 23900 7896 23906 7948
rect 24210 7896 24216 7948
rect 24268 7896 24274 7948
rect 24397 7929 24455 7935
rect 24397 7926 24409 7929
rect 24396 7895 24409 7926
rect 24443 7895 24455 7929
rect 24670 7896 24676 7948
rect 24728 7896 24734 7948
rect 24396 7889 24455 7895
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 21836 7840 22385 7868
rect 22373 7837 22385 7840
rect 22419 7868 22431 7871
rect 22646 7868 22652 7880
rect 22419 7840 22652 7868
rect 22419 7837 22431 7840
rect 22373 7831 22431 7837
rect 22646 7828 22652 7840
rect 22704 7828 22710 7880
rect 23750 7828 23756 7880
rect 23808 7868 23814 7880
rect 24121 7871 24179 7877
rect 24121 7868 24133 7871
rect 23808 7840 24133 7868
rect 23808 7828 23814 7840
rect 24121 7837 24133 7840
rect 24167 7837 24179 7871
rect 24121 7831 24179 7837
rect 22462 7800 22468 7812
rect 21315 7772 22468 7800
rect 21315 7769 21327 7772
rect 21269 7763 21327 7769
rect 22462 7760 22468 7772
rect 22520 7760 22526 7812
rect 23474 7760 23480 7812
rect 23532 7800 23538 7812
rect 23937 7803 23995 7809
rect 23937 7800 23949 7803
rect 23532 7772 23949 7800
rect 23532 7760 23538 7772
rect 23937 7769 23949 7772
rect 23983 7769 23995 7803
rect 24396 7800 24424 7889
rect 24780 7800 24808 7964
rect 25130 7896 25136 7948
rect 25188 7896 25194 7948
rect 25222 7896 25228 7948
rect 25280 7896 25286 7948
rect 23937 7763 23995 7769
rect 24325 7772 24808 7800
rect 24325 7744 24353 7772
rect 17497 7735 17555 7741
rect 17497 7732 17509 7735
rect 15580 7704 17509 7732
rect 17497 7701 17509 7704
rect 17543 7732 17555 7735
rect 17770 7732 17776 7744
rect 17543 7704 17776 7732
rect 17543 7701 17555 7704
rect 17497 7695 17555 7701
rect 17770 7692 17776 7704
rect 17828 7692 17834 7744
rect 22002 7692 22008 7744
rect 22060 7692 22066 7744
rect 23106 7692 23112 7744
rect 23164 7692 23170 7744
rect 24302 7692 24308 7744
rect 24360 7692 24366 7744
rect 24762 7692 24768 7744
rect 24820 7732 24826 7744
rect 24949 7735 25007 7741
rect 24949 7732 24961 7735
rect 24820 7704 24961 7732
rect 24820 7692 24826 7704
rect 24949 7701 24961 7704
rect 24995 7701 25007 7735
rect 24949 7695 25007 7701
rect 552 7642 27416 7664
rect 552 7590 3756 7642
rect 3808 7590 3820 7642
rect 3872 7590 3884 7642
rect 3936 7590 3948 7642
rect 4000 7590 4012 7642
rect 4064 7590 10472 7642
rect 10524 7590 10536 7642
rect 10588 7590 10600 7642
rect 10652 7590 10664 7642
rect 10716 7590 10728 7642
rect 10780 7590 17188 7642
rect 17240 7590 17252 7642
rect 17304 7590 17316 7642
rect 17368 7590 17380 7642
rect 17432 7590 17444 7642
rect 17496 7590 23904 7642
rect 23956 7590 23968 7642
rect 24020 7590 24032 7642
rect 24084 7590 24096 7642
rect 24148 7590 24160 7642
rect 24212 7590 27416 7642
rect 552 7568 27416 7590
rect 3973 7531 4031 7537
rect 3973 7497 3985 7531
rect 4019 7528 4031 7531
rect 4246 7528 4252 7540
rect 4019 7500 4252 7528
rect 4019 7497 4031 7500
rect 3973 7491 4031 7497
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 5353 7531 5411 7537
rect 5353 7497 5365 7531
rect 5399 7528 5411 7531
rect 5626 7528 5632 7540
rect 5399 7500 5632 7528
rect 5399 7497 5411 7500
rect 5353 7491 5411 7497
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 5721 7531 5779 7537
rect 5721 7497 5733 7531
rect 5767 7528 5779 7531
rect 5767 7500 6408 7528
rect 5767 7497 5779 7500
rect 5721 7491 5779 7497
rect 3234 7420 3240 7472
rect 3292 7460 3298 7472
rect 3786 7460 3792 7472
rect 3292 7432 3792 7460
rect 3292 7420 3298 7432
rect 3786 7420 3792 7432
rect 3844 7420 3850 7472
rect 3329 7395 3387 7401
rect 3329 7392 3341 7395
rect 2884 7364 3341 7392
rect 2884 7333 2912 7364
rect 3329 7361 3341 7364
rect 3375 7361 3387 7395
rect 4154 7392 4160 7404
rect 3329 7355 3387 7361
rect 3436 7364 4160 7392
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7293 2927 7327
rect 2869 7287 2927 7293
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7324 3111 7327
rect 3436 7324 3464 7364
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 6380 7392 6408 7500
rect 6454 7488 6460 7540
rect 6512 7488 6518 7540
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 11054 7528 11060 7540
rect 9180 7500 11060 7528
rect 9180 7488 9186 7500
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 11790 7488 11796 7540
rect 11848 7528 11854 7540
rect 11885 7531 11943 7537
rect 11885 7528 11897 7531
rect 11848 7500 11897 7528
rect 11848 7488 11854 7500
rect 11885 7497 11897 7500
rect 11931 7497 11943 7531
rect 11885 7491 11943 7497
rect 13354 7488 13360 7540
rect 13412 7488 13418 7540
rect 13541 7531 13599 7537
rect 13541 7497 13553 7531
rect 13587 7528 13599 7531
rect 13722 7528 13728 7540
rect 13587 7500 13728 7528
rect 13587 7497 13599 7500
rect 13541 7491 13599 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 15286 7488 15292 7540
rect 15344 7528 15350 7540
rect 16669 7531 16727 7537
rect 16669 7528 16681 7531
rect 15344 7500 16681 7528
rect 15344 7488 15350 7500
rect 16669 7497 16681 7500
rect 16715 7497 16727 7531
rect 18966 7528 18972 7540
rect 16669 7491 16727 7497
rect 16768 7500 18972 7528
rect 11149 7463 11207 7469
rect 11149 7429 11161 7463
rect 11195 7460 11207 7463
rect 13630 7460 13636 7472
rect 11195 7432 13636 7460
rect 11195 7429 11207 7432
rect 11149 7423 11207 7429
rect 13630 7420 13636 7432
rect 13688 7420 13694 7472
rect 16768 7460 16796 7500
rect 18966 7488 18972 7500
rect 19024 7488 19030 7540
rect 19794 7488 19800 7540
rect 19852 7528 19858 7540
rect 20257 7531 20315 7537
rect 20257 7528 20269 7531
rect 19852 7500 20269 7528
rect 19852 7488 19858 7500
rect 20257 7497 20269 7500
rect 20303 7528 20315 7531
rect 21174 7528 21180 7540
rect 20303 7500 21180 7528
rect 20303 7497 20315 7500
rect 20257 7491 20315 7497
rect 21174 7488 21180 7500
rect 21232 7488 21238 7540
rect 23017 7531 23075 7537
rect 23017 7497 23029 7531
rect 23063 7528 23075 7531
rect 23474 7528 23480 7540
rect 23063 7500 23480 7528
rect 23063 7497 23075 7500
rect 23017 7491 23075 7497
rect 23474 7488 23480 7500
rect 23532 7488 23538 7540
rect 24118 7488 24124 7540
rect 24176 7528 24182 7540
rect 24397 7531 24455 7537
rect 24397 7528 24409 7531
rect 24176 7500 24409 7528
rect 24176 7488 24182 7500
rect 24397 7497 24409 7500
rect 24443 7497 24455 7531
rect 24397 7491 24455 7497
rect 26878 7488 26884 7540
rect 26936 7488 26942 7540
rect 16684 7432 16796 7460
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6380 7364 7021 7392
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 7742 7352 7748 7404
rect 7800 7352 7806 7404
rect 8846 7352 8852 7404
rect 8904 7352 8910 7404
rect 12342 7392 12348 7404
rect 10612 7364 11192 7392
rect 3099 7296 3464 7324
rect 3099 7293 3111 7296
rect 3053 7287 3111 7293
rect 3510 7284 3516 7336
rect 3568 7284 3574 7336
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7293 3663 7327
rect 3605 7287 3663 7293
rect 3418 7216 3424 7268
rect 3476 7256 3482 7268
rect 3620 7256 3648 7287
rect 3694 7284 3700 7336
rect 3752 7284 3758 7336
rect 3786 7284 3792 7336
rect 3844 7284 3850 7336
rect 4614 7284 4620 7336
rect 4672 7284 4678 7336
rect 4982 7284 4988 7336
rect 5040 7284 5046 7336
rect 5626 7324 5632 7336
rect 5092 7296 5632 7324
rect 5092 7256 5120 7296
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 5997 7327 6055 7333
rect 5997 7293 6009 7327
rect 6043 7293 6055 7327
rect 5997 7287 6055 7293
rect 3476 7228 5120 7256
rect 5353 7259 5411 7265
rect 3476 7216 3482 7228
rect 5353 7225 5365 7259
rect 5399 7256 5411 7259
rect 5810 7256 5816 7268
rect 5399 7228 5816 7256
rect 5399 7225 5411 7228
rect 5353 7219 5411 7225
rect 5810 7216 5816 7228
rect 5868 7216 5874 7268
rect 6012 7256 6040 7287
rect 6086 7284 6092 7336
rect 6144 7284 6150 7336
rect 6181 7327 6239 7333
rect 6181 7293 6193 7327
rect 6227 7324 6239 7327
rect 6365 7327 6423 7333
rect 6227 7296 6316 7324
rect 6227 7293 6239 7296
rect 6181 7287 6239 7293
rect 6012 7228 6132 7256
rect 6104 7200 6132 7228
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 2961 7191 3019 7197
rect 2961 7188 2973 7191
rect 2832 7160 2973 7188
rect 2832 7148 2838 7160
rect 2961 7157 2973 7160
rect 3007 7157 3019 7191
rect 2961 7151 3019 7157
rect 3326 7148 3332 7200
rect 3384 7188 3390 7200
rect 4246 7188 4252 7200
rect 3384 7160 4252 7188
rect 3384 7148 3390 7160
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 5537 7191 5595 7197
rect 5537 7157 5549 7191
rect 5583 7188 5595 7191
rect 5994 7188 6000 7200
rect 5583 7160 6000 7188
rect 5583 7157 5595 7160
rect 5537 7151 5595 7157
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 6086 7148 6092 7200
rect 6144 7148 6150 7200
rect 6288 7188 6316 7296
rect 6365 7293 6377 7327
rect 6411 7324 6423 7327
rect 6730 7324 6736 7336
rect 6411 7296 6736 7324
rect 6411 7293 6423 7296
rect 6365 7287 6423 7293
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 8110 7284 8116 7336
rect 8168 7324 8174 7336
rect 10612 7333 10640 7364
rect 11164 7336 11192 7364
rect 11624 7364 12348 7392
rect 9105 7327 9163 7333
rect 9105 7324 9117 7327
rect 8168 7296 9117 7324
rect 8168 7284 8174 7296
rect 9105 7293 9117 7296
rect 9151 7293 9163 7327
rect 9105 7287 9163 7293
rect 10597 7327 10655 7333
rect 10597 7293 10609 7327
rect 10643 7293 10655 7327
rect 10597 7287 10655 7293
rect 10689 7327 10747 7333
rect 10689 7293 10701 7327
rect 10735 7324 10747 7327
rect 10778 7324 10784 7336
rect 10735 7296 10784 7324
rect 10735 7293 10747 7296
rect 10689 7287 10747 7293
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7293 10931 7327
rect 10873 7287 10931 7293
rect 10965 7327 11023 7333
rect 10965 7293 10977 7327
rect 11011 7324 11023 7327
rect 11054 7324 11060 7336
rect 11011 7296 11060 7324
rect 11011 7293 11023 7296
rect 10965 7287 11023 7293
rect 10318 7216 10324 7268
rect 10376 7256 10382 7268
rect 10888 7256 10916 7287
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 11146 7284 11152 7336
rect 11204 7284 11210 7336
rect 11241 7327 11299 7333
rect 11241 7293 11253 7327
rect 11287 7293 11299 7327
rect 11241 7287 11299 7293
rect 10376 7228 10916 7256
rect 11256 7256 11284 7287
rect 11422 7284 11428 7336
rect 11480 7284 11486 7336
rect 11514 7284 11520 7336
rect 11572 7284 11578 7336
rect 11624 7333 11652 7364
rect 12342 7352 12348 7364
rect 12400 7392 12406 7404
rect 12400 7364 13124 7392
rect 12400 7352 12406 7364
rect 11609 7327 11667 7333
rect 11609 7293 11621 7327
rect 11655 7293 11667 7327
rect 11609 7287 11667 7293
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 13096 7333 13124 7364
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 12124 7296 12725 7324
rect 12124 7284 12130 7296
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 12861 7327 12919 7333
rect 12861 7293 12873 7327
rect 12907 7324 12919 7327
rect 13081 7327 13139 7333
rect 12907 7293 12940 7324
rect 12861 7287 12940 7293
rect 13081 7293 13093 7327
rect 13127 7293 13139 7327
rect 13081 7287 13139 7293
rect 12618 7256 12624 7268
rect 11256 7228 12624 7256
rect 10376 7216 10382 7228
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 7006 7188 7012 7200
rect 6288 7160 7012 7188
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 7193 7191 7251 7197
rect 7193 7157 7205 7191
rect 7239 7188 7251 7191
rect 7466 7188 7472 7200
rect 7239 7160 7472 7188
rect 7239 7157 7251 7160
rect 7193 7151 7251 7157
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 10229 7191 10287 7197
rect 10229 7188 10241 7191
rect 8352 7160 10241 7188
rect 8352 7148 8358 7160
rect 10229 7157 10241 7160
rect 10275 7188 10287 7191
rect 12912 7188 12940 7287
rect 13170 7284 13176 7336
rect 13228 7333 13234 7336
rect 13228 7324 13236 7333
rect 13228 7296 13273 7324
rect 13228 7287 13236 7296
rect 13228 7284 13234 7287
rect 14182 7284 14188 7336
rect 14240 7324 14246 7336
rect 14654 7327 14712 7333
rect 14654 7324 14666 7327
rect 14240 7296 14666 7324
rect 14240 7284 14246 7296
rect 14654 7293 14666 7296
rect 14700 7293 14712 7327
rect 14654 7287 14712 7293
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7324 14979 7327
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 14967 7296 15117 7324
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 15105 7293 15117 7296
rect 15151 7324 15163 7327
rect 16574 7324 16580 7336
rect 15151 7296 16580 7324
rect 15151 7293 15163 7296
rect 15105 7287 15163 7293
rect 16574 7284 16580 7296
rect 16632 7284 16638 7336
rect 12989 7259 13047 7265
rect 12989 7225 13001 7259
rect 13035 7256 13047 7259
rect 13262 7256 13268 7268
rect 13035 7228 13268 7256
rect 13035 7225 13047 7228
rect 12989 7219 13047 7225
rect 13262 7216 13268 7228
rect 13320 7216 13326 7268
rect 15378 7265 15384 7268
rect 15372 7219 15384 7265
rect 15436 7256 15442 7268
rect 16684 7256 16712 7432
rect 18046 7420 18052 7472
rect 18104 7460 18110 7472
rect 20717 7463 20775 7469
rect 20717 7460 20729 7463
rect 18104 7432 20729 7460
rect 18104 7420 18110 7432
rect 20717 7429 20729 7432
rect 20763 7429 20775 7463
rect 20717 7423 20775 7429
rect 22833 7463 22891 7469
rect 22833 7429 22845 7463
rect 22879 7460 22891 7463
rect 23566 7460 23572 7472
rect 22879 7432 23572 7460
rect 22879 7429 22891 7432
rect 22833 7423 22891 7429
rect 23566 7420 23572 7432
rect 23624 7420 23630 7472
rect 24578 7420 24584 7472
rect 24636 7460 24642 7472
rect 25314 7460 25320 7472
rect 24636 7432 25320 7460
rect 24636 7420 24642 7432
rect 25314 7420 25320 7432
rect 25372 7460 25378 7472
rect 25372 7432 25544 7460
rect 25372 7420 25378 7432
rect 17862 7352 17868 7404
rect 17920 7392 17926 7404
rect 18230 7392 18236 7404
rect 17920 7364 18236 7392
rect 17920 7352 17926 7364
rect 18230 7352 18236 7364
rect 18288 7352 18294 7404
rect 19334 7352 19340 7404
rect 19392 7352 19398 7404
rect 24029 7395 24087 7401
rect 24029 7361 24041 7395
rect 24075 7392 24087 7395
rect 24762 7392 24768 7404
rect 24075 7364 24768 7392
rect 24075 7361 24087 7364
rect 24029 7355 24087 7361
rect 24762 7352 24768 7364
rect 24820 7352 24826 7404
rect 25516 7401 25544 7432
rect 25501 7395 25559 7401
rect 25501 7361 25513 7395
rect 25547 7361 25559 7395
rect 25501 7355 25559 7361
rect 16850 7284 16856 7336
rect 16908 7284 16914 7336
rect 16942 7284 16948 7336
rect 17000 7324 17006 7336
rect 17589 7327 17647 7333
rect 17589 7324 17601 7327
rect 17000 7296 17601 7324
rect 17000 7284 17006 7296
rect 17589 7293 17601 7296
rect 17635 7324 17647 7327
rect 18785 7327 18843 7333
rect 18785 7324 18797 7327
rect 17635 7296 18797 7324
rect 17635 7293 17647 7296
rect 17589 7287 17647 7293
rect 18785 7293 18797 7296
rect 18831 7293 18843 7327
rect 18785 7287 18843 7293
rect 19610 7284 19616 7336
rect 19668 7324 19674 7336
rect 20625 7327 20683 7333
rect 20625 7324 20637 7327
rect 19668 7296 20637 7324
rect 19668 7284 19674 7296
rect 20625 7293 20637 7296
rect 20671 7293 20683 7327
rect 20625 7287 20683 7293
rect 20809 7327 20867 7333
rect 20809 7293 20821 7327
rect 20855 7293 20867 7327
rect 20809 7287 20867 7293
rect 21453 7327 21511 7333
rect 21453 7293 21465 7327
rect 21499 7293 21511 7327
rect 21453 7287 21511 7293
rect 21720 7327 21778 7333
rect 21720 7293 21732 7327
rect 21766 7324 21778 7327
rect 22002 7324 22008 7336
rect 21766 7296 22008 7324
rect 21766 7293 21778 7296
rect 21720 7287 21778 7293
rect 15436 7228 15472 7256
rect 16408 7228 16712 7256
rect 20165 7259 20223 7265
rect 15378 7216 15384 7219
rect 15436 7216 15442 7228
rect 13354 7188 13360 7200
rect 10275 7160 13360 7188
rect 10275 7157 10287 7160
rect 10229 7151 10287 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 15010 7148 15016 7200
rect 15068 7188 15074 7200
rect 16408 7188 16436 7228
rect 20165 7225 20177 7259
rect 20211 7256 20223 7259
rect 20211 7228 20300 7256
rect 20211 7225 20223 7228
rect 20165 7219 20223 7225
rect 15068 7160 16436 7188
rect 15068 7148 15074 7160
rect 16482 7148 16488 7200
rect 16540 7148 16546 7200
rect 19981 7191 20039 7197
rect 19981 7157 19993 7191
rect 20027 7188 20039 7191
rect 20070 7188 20076 7200
rect 20027 7160 20076 7188
rect 20027 7157 20039 7160
rect 19981 7151 20039 7157
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 20272 7188 20300 7228
rect 20346 7216 20352 7268
rect 20404 7256 20410 7268
rect 20824 7256 20852 7287
rect 20404 7228 20852 7256
rect 21468 7256 21496 7287
rect 22002 7284 22008 7296
rect 22060 7284 22066 7336
rect 22922 7284 22928 7336
rect 22980 7284 22986 7336
rect 23106 7284 23112 7336
rect 23164 7284 23170 7336
rect 23474 7284 23480 7336
rect 23532 7324 23538 7336
rect 23937 7327 23995 7333
rect 23937 7324 23949 7327
rect 23532 7296 23949 7324
rect 23532 7284 23538 7296
rect 23937 7293 23949 7296
rect 23983 7293 23995 7327
rect 23937 7287 23995 7293
rect 24121 7327 24179 7333
rect 24121 7293 24133 7327
rect 24167 7324 24179 7327
rect 24210 7324 24216 7336
rect 24167 7296 24216 7324
rect 24167 7293 24179 7296
rect 24121 7287 24179 7293
rect 24210 7284 24216 7296
rect 24268 7284 24274 7336
rect 24854 7324 24860 7336
rect 24412 7296 24860 7324
rect 24412 7268 24440 7296
rect 24854 7284 24860 7296
rect 24912 7284 24918 7336
rect 25774 7333 25780 7336
rect 25409 7327 25467 7333
rect 25409 7293 25421 7327
rect 25455 7293 25467 7327
rect 25768 7324 25780 7333
rect 25735 7296 25780 7324
rect 25409 7287 25467 7293
rect 25768 7287 25780 7296
rect 21818 7256 21824 7268
rect 21468 7228 21824 7256
rect 20404 7216 20410 7228
rect 21818 7216 21824 7228
rect 21876 7216 21882 7268
rect 23658 7216 23664 7268
rect 23716 7256 23722 7268
rect 24394 7265 24400 7268
rect 24381 7259 24400 7265
rect 23716 7228 24348 7256
rect 23716 7216 23722 7228
rect 20530 7188 20536 7200
rect 20272 7160 20536 7188
rect 20530 7148 20536 7160
rect 20588 7188 20594 7200
rect 21358 7188 21364 7200
rect 20588 7160 21364 7188
rect 20588 7148 20594 7160
rect 21358 7148 21364 7160
rect 21416 7148 21422 7200
rect 23750 7148 23756 7200
rect 23808 7188 23814 7200
rect 24213 7191 24271 7197
rect 24213 7188 24225 7191
rect 23808 7160 24225 7188
rect 23808 7148 23814 7160
rect 24213 7157 24225 7160
rect 24259 7157 24271 7191
rect 24320 7188 24348 7228
rect 24381 7225 24393 7259
rect 24381 7219 24400 7225
rect 24394 7216 24400 7219
rect 24452 7216 24458 7268
rect 24486 7216 24492 7268
rect 24544 7256 24550 7268
rect 24581 7259 24639 7265
rect 24581 7256 24593 7259
rect 24544 7228 24593 7256
rect 24544 7216 24550 7228
rect 24581 7225 24593 7228
rect 24627 7256 24639 7259
rect 25038 7256 25044 7268
rect 24627 7228 25044 7256
rect 24627 7225 24639 7228
rect 24581 7219 24639 7225
rect 25038 7216 25044 7228
rect 25096 7216 25102 7268
rect 25424 7256 25452 7287
rect 25774 7284 25780 7287
rect 25832 7284 25838 7336
rect 25866 7256 25872 7268
rect 25424 7228 25872 7256
rect 25866 7216 25872 7228
rect 25924 7216 25930 7268
rect 24765 7191 24823 7197
rect 24765 7188 24777 7191
rect 24320 7160 24777 7188
rect 24213 7151 24271 7157
rect 24765 7157 24777 7160
rect 24811 7157 24823 7191
rect 24765 7151 24823 7157
rect 552 7098 27576 7120
rect 552 7046 7114 7098
rect 7166 7046 7178 7098
rect 7230 7046 7242 7098
rect 7294 7046 7306 7098
rect 7358 7046 7370 7098
rect 7422 7046 13830 7098
rect 13882 7046 13894 7098
rect 13946 7046 13958 7098
rect 14010 7046 14022 7098
rect 14074 7046 14086 7098
rect 14138 7046 20546 7098
rect 20598 7046 20610 7098
rect 20662 7046 20674 7098
rect 20726 7046 20738 7098
rect 20790 7046 20802 7098
rect 20854 7046 27262 7098
rect 27314 7046 27326 7098
rect 27378 7046 27390 7098
rect 27442 7046 27454 7098
rect 27506 7046 27518 7098
rect 27570 7046 27576 7098
rect 552 7024 27576 7046
rect 3694 6944 3700 6996
rect 3752 6984 3758 6996
rect 3881 6987 3939 6993
rect 3881 6984 3893 6987
rect 3752 6956 3893 6984
rect 3752 6944 3758 6956
rect 3881 6953 3893 6956
rect 3927 6984 3939 6987
rect 4614 6984 4620 6996
rect 3927 6956 4620 6984
rect 3927 6953 3939 6956
rect 3881 6947 3939 6953
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 6086 6944 6092 6996
rect 6144 6984 6150 6996
rect 6144 6956 7512 6984
rect 6144 6944 6150 6956
rect 7484 6928 7512 6956
rect 8202 6944 8208 6996
rect 8260 6944 8266 6996
rect 9398 6944 9404 6996
rect 9456 6984 9462 6996
rect 9456 6956 10824 6984
rect 9456 6944 9462 6956
rect 10796 6928 10824 6956
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 11112 6956 11376 6984
rect 11112 6944 11118 6956
rect 6178 6916 6184 6928
rect 2608 6888 3004 6916
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 2501 6851 2559 6857
rect 2501 6848 2513 6851
rect 1636 6820 2513 6848
rect 1636 6808 1642 6820
rect 2501 6817 2513 6820
rect 2547 6848 2559 6851
rect 2608 6848 2636 6888
rect 2774 6857 2780 6860
rect 2547 6820 2636 6848
rect 2547 6817 2559 6820
rect 2501 6811 2559 6817
rect 2768 6811 2780 6857
rect 2832 6848 2838 6860
rect 2976 6848 3004 6888
rect 4172 6888 6184 6916
rect 4172 6860 4200 6888
rect 6178 6876 6184 6888
rect 6236 6876 6242 6928
rect 7466 6876 7472 6928
rect 7524 6916 7530 6928
rect 8481 6919 8539 6925
rect 8481 6916 8493 6919
rect 7524 6888 8493 6916
rect 7524 6876 7530 6888
rect 8481 6885 8493 6888
rect 8527 6885 8539 6919
rect 9737 6919 9795 6925
rect 9737 6916 9749 6919
rect 8481 6879 8539 6885
rect 9048 6888 9749 6916
rect 4154 6848 4160 6860
rect 2832 6820 2868 6848
rect 2976 6820 4160 6848
rect 2774 6808 2780 6811
rect 2832 6808 2838 6820
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 4424 6851 4482 6857
rect 4424 6817 4436 6851
rect 4470 6848 4482 6851
rect 5718 6848 5724 6860
rect 4470 6820 5724 6848
rect 4470 6817 4482 6820
rect 4424 6811 4482 6817
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 7834 6808 7840 6860
rect 7892 6808 7898 6860
rect 8386 6857 8392 6860
rect 8384 6848 8392 6857
rect 8347 6820 8392 6848
rect 8384 6811 8392 6820
rect 8386 6808 8392 6811
rect 8444 6808 8450 6860
rect 8570 6808 8576 6860
rect 8628 6808 8634 6860
rect 8662 6808 8668 6860
rect 8720 6857 8726 6860
rect 8720 6851 8759 6857
rect 8747 6817 8759 6851
rect 8720 6811 8759 6817
rect 8720 6808 8726 6811
rect 8846 6808 8852 6860
rect 8904 6808 8910 6860
rect 8938 6808 8944 6860
rect 8996 6848 9002 6860
rect 9048 6848 9076 6888
rect 9737 6885 9749 6888
rect 9783 6885 9795 6919
rect 9737 6879 9795 6885
rect 9950 6876 9956 6928
rect 10008 6876 10014 6928
rect 10778 6876 10784 6928
rect 10836 6916 10842 6928
rect 10836 6888 11100 6916
rect 10836 6876 10842 6888
rect 8996 6820 9076 6848
rect 8996 6808 9002 6820
rect 9122 6808 9128 6860
rect 9180 6808 9186 6860
rect 9217 6851 9275 6857
rect 9217 6817 9229 6851
rect 9263 6817 9275 6851
rect 9217 6811 9275 6817
rect 9232 6780 9260 6811
rect 9398 6808 9404 6860
rect 9456 6808 9462 6860
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 9048 6752 9260 6780
rect 7006 6672 7012 6724
rect 7064 6712 7070 6724
rect 8941 6715 8999 6721
rect 8941 6712 8953 6715
rect 7064 6684 8953 6712
rect 7064 6672 7070 6684
rect 8941 6681 8953 6684
rect 8987 6681 8999 6715
rect 8941 6675 8999 6681
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 6270 6644 6276 6656
rect 5592 6616 6276 6644
rect 5592 6604 5598 6616
rect 6270 6604 6276 6616
rect 6328 6644 6334 6656
rect 9048 6644 9076 6752
rect 9214 6672 9220 6724
rect 9272 6712 9278 6724
rect 9508 6712 9536 6811
rect 10042 6808 10048 6860
rect 10100 6808 10106 6860
rect 11072 6857 11100 6888
rect 11348 6857 11376 6956
rect 11422 6944 11428 6996
rect 11480 6984 11486 6996
rect 11517 6987 11575 6993
rect 11517 6984 11529 6987
rect 11480 6956 11529 6984
rect 11480 6944 11486 6956
rect 11517 6953 11529 6956
rect 11563 6953 11575 6987
rect 11517 6947 11575 6953
rect 12161 6987 12219 6993
rect 12161 6953 12173 6987
rect 12207 6984 12219 6987
rect 12250 6984 12256 6996
rect 12207 6956 12256 6984
rect 12207 6953 12219 6956
rect 12161 6947 12219 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 16482 6984 16488 6996
rect 12860 6956 16488 6984
rect 12860 6944 12866 6956
rect 16482 6944 16488 6956
rect 16540 6944 16546 6996
rect 20254 6944 20260 6996
rect 20312 6984 20318 6996
rect 20622 6984 20628 6996
rect 20312 6956 20628 6984
rect 20312 6944 20318 6956
rect 20622 6944 20628 6956
rect 20680 6984 20686 6996
rect 24029 6987 24087 6993
rect 20680 6956 21128 6984
rect 20680 6944 20686 6956
rect 12710 6876 12716 6928
rect 12768 6916 12774 6928
rect 12989 6919 13047 6925
rect 12989 6916 13001 6919
rect 12768 6888 13001 6916
rect 12768 6876 12774 6888
rect 12989 6885 13001 6888
rect 13035 6916 13047 6919
rect 13170 6916 13176 6928
rect 13035 6888 13176 6916
rect 13035 6885 13047 6888
rect 12989 6879 13047 6885
rect 13170 6876 13176 6888
rect 13228 6916 13234 6928
rect 17770 6916 17776 6928
rect 13228 6888 17776 6916
rect 13228 6876 13234 6888
rect 17770 6876 17776 6888
rect 17828 6876 17834 6928
rect 19610 6876 19616 6928
rect 19668 6916 19674 6928
rect 20717 6919 20775 6925
rect 19668 6888 20024 6916
rect 19668 6876 19674 6888
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 10152 6820 10977 6848
rect 9858 6740 9864 6792
rect 9916 6780 9922 6792
rect 10152 6780 10180 6820
rect 10965 6817 10977 6820
rect 11011 6817 11023 6851
rect 10965 6811 11023 6817
rect 11057 6851 11115 6857
rect 11057 6817 11069 6851
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 11241 6851 11299 6857
rect 11241 6817 11253 6851
rect 11287 6817 11299 6851
rect 11241 6811 11299 6817
rect 11333 6851 11391 6857
rect 11333 6817 11345 6851
rect 11379 6848 11391 6851
rect 12253 6851 12311 6857
rect 11379 6820 11560 6848
rect 11379 6817 11391 6820
rect 11333 6811 11391 6817
rect 9916 6752 10180 6780
rect 10321 6783 10379 6789
rect 9916 6740 9922 6752
rect 10321 6749 10333 6783
rect 10367 6780 10379 6783
rect 10410 6780 10416 6792
rect 10367 6752 10416 6780
rect 10367 6749 10379 6752
rect 10321 6743 10379 6749
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 11256 6780 11284 6811
rect 11422 6780 11428 6792
rect 11256 6752 11428 6780
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11532 6780 11560 6820
rect 12253 6817 12265 6851
rect 12299 6848 12311 6851
rect 12894 6848 12900 6860
rect 12299 6820 12900 6848
rect 12299 6817 12311 6820
rect 12253 6811 12311 6817
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 17856 6851 17914 6857
rect 17856 6817 17868 6851
rect 17902 6848 17914 6851
rect 19061 6851 19119 6857
rect 19061 6848 19073 6851
rect 17902 6820 19073 6848
rect 17902 6817 17914 6820
rect 17856 6811 17914 6817
rect 19061 6817 19073 6820
rect 19107 6817 19119 6851
rect 19061 6811 19119 6817
rect 19334 6808 19340 6860
rect 19392 6848 19398 6860
rect 19996 6857 20024 6888
rect 20717 6885 20729 6919
rect 20763 6916 20775 6919
rect 20990 6916 20996 6928
rect 20763 6888 20996 6916
rect 20763 6885 20775 6888
rect 20717 6879 20775 6885
rect 19797 6851 19855 6857
rect 19797 6848 19809 6851
rect 19392 6820 19809 6848
rect 19392 6808 19398 6820
rect 19797 6817 19809 6820
rect 19843 6817 19855 6851
rect 19797 6811 19855 6817
rect 19981 6851 20039 6857
rect 19981 6817 19993 6851
rect 20027 6817 20039 6851
rect 19981 6811 20039 6817
rect 20070 6808 20076 6860
rect 20128 6848 20134 6860
rect 20257 6851 20315 6857
rect 20257 6848 20269 6851
rect 20128 6820 20269 6848
rect 20128 6808 20134 6820
rect 20257 6817 20269 6820
rect 20303 6817 20315 6851
rect 20732 6848 20760 6879
rect 20990 6876 20996 6888
rect 21048 6876 21054 6928
rect 20257 6811 20315 6817
rect 20364 6820 20760 6848
rect 12437 6783 12495 6789
rect 12437 6780 12449 6783
rect 11532 6752 12449 6780
rect 12437 6749 12449 6752
rect 12483 6780 12495 6783
rect 12483 6752 13032 6780
rect 12483 6749 12495 6752
rect 12437 6743 12495 6749
rect 9272 6684 9536 6712
rect 9272 6672 9278 6684
rect 9582 6672 9588 6724
rect 9640 6712 9646 6724
rect 11238 6712 11244 6724
rect 9640 6684 11244 6712
rect 9640 6672 9646 6684
rect 11238 6672 11244 6684
rect 11296 6672 11302 6724
rect 11698 6672 11704 6724
rect 11756 6712 11762 6724
rect 11793 6715 11851 6721
rect 11793 6712 11805 6715
rect 11756 6684 11805 6712
rect 11756 6672 11762 6684
rect 11793 6681 11805 6684
rect 11839 6681 11851 6715
rect 13004 6712 13032 6752
rect 13078 6740 13084 6792
rect 13136 6740 13142 6792
rect 13265 6783 13323 6789
rect 13265 6749 13277 6783
rect 13311 6780 13323 6783
rect 13446 6780 13452 6792
rect 13311 6752 13452 6780
rect 13311 6749 13323 6752
rect 13265 6743 13323 6749
rect 13280 6712 13308 6743
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 17586 6740 17592 6792
rect 17644 6740 17650 6792
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 20165 6783 20223 6789
rect 20165 6749 20177 6783
rect 20211 6780 20223 6783
rect 20364 6780 20392 6820
rect 20806 6808 20812 6860
rect 20864 6808 20870 6860
rect 20898 6808 20904 6860
rect 20956 6808 20962 6860
rect 21100 6857 21128 6956
rect 24029 6953 24041 6987
rect 24075 6984 24087 6987
rect 24394 6984 24400 6996
rect 24075 6956 24400 6984
rect 24075 6953 24087 6956
rect 24029 6947 24087 6953
rect 24394 6944 24400 6956
rect 24452 6944 24458 6996
rect 25866 6984 25872 6996
rect 24596 6956 25872 6984
rect 23845 6919 23903 6925
rect 23845 6885 23857 6919
rect 23891 6916 23903 6919
rect 24302 6916 24308 6928
rect 23891 6888 24308 6916
rect 23891 6885 23903 6888
rect 23845 6879 23903 6885
rect 24302 6876 24308 6888
rect 24360 6876 24366 6928
rect 24596 6916 24624 6956
rect 25866 6944 25872 6956
rect 25924 6944 25930 6996
rect 24412 6888 24624 6916
rect 21085 6851 21143 6857
rect 21085 6817 21097 6851
rect 21131 6817 21143 6851
rect 21085 6811 21143 6817
rect 21729 6851 21787 6857
rect 21729 6817 21741 6851
rect 21775 6817 21787 6851
rect 23566 6848 23572 6860
rect 21729 6811 21787 6817
rect 22066 6820 23572 6848
rect 20211 6752 20392 6780
rect 20211 6749 20223 6752
rect 20165 6743 20223 6749
rect 20438 6740 20444 6792
rect 20496 6780 20502 6792
rect 21744 6780 21772 6811
rect 20496 6752 21772 6780
rect 20496 6740 20502 6752
rect 20349 6715 20407 6721
rect 20349 6712 20361 6715
rect 11793 6675 11851 6681
rect 11900 6684 12940 6712
rect 13004 6684 13308 6712
rect 18524 6684 20361 6712
rect 6328 6616 9076 6644
rect 6328 6604 6334 6616
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 9769 6647 9827 6653
rect 9769 6644 9781 6647
rect 9548 6616 9781 6644
rect 9548 6604 9554 6616
rect 9769 6613 9781 6616
rect 9815 6613 9827 6647
rect 9769 6607 9827 6613
rect 10134 6604 10140 6656
rect 10192 6604 10198 6656
rect 10226 6604 10232 6656
rect 10284 6604 10290 6656
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 11054 6644 11060 6656
rect 10468 6616 11060 6644
rect 10468 6604 10474 6616
rect 11054 6604 11060 6616
rect 11112 6644 11118 6656
rect 11900 6644 11928 6684
rect 11112 6616 11928 6644
rect 11112 6604 11118 6616
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 12621 6647 12679 6653
rect 12621 6644 12633 6647
rect 12216 6616 12633 6644
rect 12216 6604 12222 6616
rect 12621 6613 12633 6616
rect 12667 6613 12679 6647
rect 12912 6644 12940 6684
rect 16298 6644 16304 6656
rect 12912 6616 16304 6644
rect 12621 6607 12679 6613
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 18322 6604 18328 6656
rect 18380 6644 18386 6656
rect 18524 6644 18552 6684
rect 20349 6681 20361 6684
rect 20395 6681 20407 6715
rect 22066 6712 22094 6820
rect 23566 6808 23572 6820
rect 23624 6848 23630 6860
rect 24118 6848 24124 6860
rect 23624 6820 24124 6848
rect 23624 6808 23630 6820
rect 24118 6808 24124 6820
rect 24176 6808 24182 6860
rect 24412 6857 24440 6888
rect 24213 6851 24271 6857
rect 24213 6817 24225 6851
rect 24259 6817 24271 6851
rect 24213 6811 24271 6817
rect 24397 6851 24455 6857
rect 24397 6817 24409 6851
rect 24443 6817 24455 6851
rect 24397 6811 24455 6817
rect 24489 6851 24547 6857
rect 24489 6817 24501 6851
rect 24535 6848 24547 6851
rect 24578 6848 24584 6860
rect 24535 6820 24584 6848
rect 24535 6817 24547 6820
rect 24489 6811 24547 6817
rect 20349 6675 20407 6681
rect 21192 6684 22094 6712
rect 24228 6712 24256 6811
rect 24578 6808 24584 6820
rect 24636 6808 24642 6860
rect 24762 6857 24768 6860
rect 24756 6811 24768 6857
rect 24820 6848 24826 6860
rect 26145 6851 26203 6857
rect 24820 6820 24856 6848
rect 24762 6808 24768 6811
rect 24820 6808 24826 6820
rect 26145 6817 26157 6851
rect 26191 6848 26203 6851
rect 26421 6851 26479 6857
rect 26421 6848 26433 6851
rect 26191 6820 26433 6848
rect 26191 6817 26203 6820
rect 26145 6811 26203 6817
rect 26421 6817 26433 6820
rect 26467 6817 26479 6851
rect 26421 6811 26479 6817
rect 25866 6740 25872 6792
rect 25924 6780 25930 6792
rect 26973 6783 27031 6789
rect 26973 6780 26985 6783
rect 25924 6752 26985 6780
rect 25924 6740 25930 6752
rect 26973 6749 26985 6752
rect 27019 6749 27031 6783
rect 26973 6743 27031 6749
rect 24394 6712 24400 6724
rect 24228 6684 24400 6712
rect 18380 6616 18552 6644
rect 18969 6647 19027 6653
rect 18380 6604 18386 6616
rect 18969 6613 18981 6647
rect 19015 6644 19027 6647
rect 19334 6644 19340 6656
rect 19015 6616 19340 6644
rect 19015 6613 19027 6616
rect 18969 6607 19027 6613
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 19702 6604 19708 6656
rect 19760 6644 19766 6656
rect 20070 6644 20076 6656
rect 19760 6616 20076 6644
rect 19760 6604 19766 6616
rect 20070 6604 20076 6616
rect 20128 6604 20134 6656
rect 20254 6604 20260 6656
rect 20312 6644 20318 6656
rect 20533 6647 20591 6653
rect 20533 6644 20545 6647
rect 20312 6616 20545 6644
rect 20312 6604 20318 6616
rect 20533 6613 20545 6616
rect 20579 6644 20591 6647
rect 21192 6644 21220 6684
rect 24394 6672 24400 6684
rect 24452 6672 24458 6724
rect 26053 6715 26111 6721
rect 26053 6712 26065 6715
rect 25424 6684 26065 6712
rect 20579 6616 21220 6644
rect 20579 6613 20591 6616
rect 20533 6607 20591 6613
rect 22370 6604 22376 6656
rect 22428 6644 22434 6656
rect 23017 6647 23075 6653
rect 23017 6644 23029 6647
rect 22428 6616 23029 6644
rect 22428 6604 22434 6616
rect 23017 6613 23029 6616
rect 23063 6613 23075 6647
rect 23017 6607 23075 6613
rect 24302 6604 24308 6656
rect 24360 6644 24366 6656
rect 25424 6644 25452 6684
rect 26053 6681 26065 6684
rect 26099 6681 26111 6715
rect 26053 6675 26111 6681
rect 24360 6616 25452 6644
rect 24360 6604 24366 6616
rect 552 6554 27416 6576
rect 552 6502 3756 6554
rect 3808 6502 3820 6554
rect 3872 6502 3884 6554
rect 3936 6502 3948 6554
rect 4000 6502 4012 6554
rect 4064 6502 10472 6554
rect 10524 6502 10536 6554
rect 10588 6502 10600 6554
rect 10652 6502 10664 6554
rect 10716 6502 10728 6554
rect 10780 6502 17188 6554
rect 17240 6502 17252 6554
rect 17304 6502 17316 6554
rect 17368 6502 17380 6554
rect 17432 6502 17444 6554
rect 17496 6502 23904 6554
rect 23956 6502 23968 6554
rect 24020 6502 24032 6554
rect 24084 6502 24096 6554
rect 24148 6502 24160 6554
rect 24212 6502 27416 6554
rect 552 6480 27416 6502
rect 4982 6400 4988 6452
rect 5040 6400 5046 6452
rect 5442 6400 5448 6452
rect 5500 6440 5506 6452
rect 5500 6412 5672 6440
rect 5500 6400 5506 6412
rect 5534 6332 5540 6384
rect 5592 6332 5598 6384
rect 5644 6372 5672 6412
rect 5810 6400 5816 6452
rect 5868 6400 5874 6452
rect 9030 6440 9036 6452
rect 6104 6412 9036 6440
rect 6104 6372 6132 6412
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 9401 6443 9459 6449
rect 9401 6409 9413 6443
rect 9447 6440 9459 6443
rect 10042 6440 10048 6452
rect 9447 6412 10048 6440
rect 9447 6409 9459 6412
rect 9401 6403 9459 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10318 6400 10324 6452
rect 10376 6400 10382 6452
rect 11238 6400 11244 6452
rect 11296 6400 11302 6452
rect 11330 6400 11336 6452
rect 11388 6440 11394 6452
rect 14550 6440 14556 6452
rect 11388 6412 14556 6440
rect 11388 6400 11394 6412
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 17678 6400 17684 6452
rect 17736 6400 17742 6452
rect 18509 6443 18567 6449
rect 18509 6409 18521 6443
rect 18555 6440 18567 6443
rect 19610 6440 19616 6452
rect 18555 6412 19616 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 19610 6400 19616 6412
rect 19668 6400 19674 6452
rect 21266 6440 21272 6452
rect 20640 6412 21272 6440
rect 5644 6344 6132 6372
rect 6104 6313 6132 6344
rect 6178 6332 6184 6384
rect 6236 6372 6242 6384
rect 9582 6372 9588 6384
rect 6236 6344 6592 6372
rect 6236 6332 6242 6344
rect 6089 6307 6147 6313
rect 6089 6273 6101 6307
rect 6135 6273 6147 6307
rect 6089 6267 6147 6273
rect 6270 6264 6276 6316
rect 6328 6264 6334 6316
rect 6564 6313 6592 6344
rect 8588 6344 9588 6372
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 3510 6196 3516 6248
rect 3568 6236 3574 6248
rect 5169 6239 5227 6245
rect 5169 6236 5181 6239
rect 3568 6208 5181 6236
rect 3568 6196 3574 6208
rect 5169 6205 5181 6208
rect 5215 6236 5227 6239
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 5215 6208 6009 6236
rect 5215 6205 5227 6208
rect 5169 6199 5227 6205
rect 5997 6205 6009 6208
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 6181 6239 6239 6245
rect 6181 6205 6193 6239
rect 6227 6236 6239 6239
rect 7558 6236 7564 6248
rect 6227 6208 7564 6236
rect 6227 6205 6239 6208
rect 6181 6199 6239 6205
rect 4614 6128 4620 6180
rect 4672 6168 4678 6180
rect 4672 6140 5396 6168
rect 4672 6128 4678 6140
rect 5258 6060 5264 6112
rect 5316 6060 5322 6112
rect 5368 6109 5396 6140
rect 5353 6103 5411 6109
rect 5353 6069 5365 6103
rect 5399 6100 5411 6103
rect 6196 6100 6224 6199
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 7742 6196 7748 6248
rect 7800 6236 7806 6248
rect 8021 6239 8079 6245
rect 8021 6236 8033 6239
rect 7800 6208 8033 6236
rect 7800 6196 7806 6208
rect 8021 6205 8033 6208
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 8202 6196 8208 6248
rect 8260 6196 8266 6248
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6236 8539 6239
rect 8588 6236 8616 6344
rect 9582 6332 9588 6344
rect 9640 6332 9646 6384
rect 10965 6375 11023 6381
rect 10965 6341 10977 6375
rect 11011 6372 11023 6375
rect 19978 6372 19984 6384
rect 11011 6344 11652 6372
rect 11011 6341 11023 6344
rect 10965 6335 11023 6341
rect 10226 6304 10232 6316
rect 8680 6276 10232 6304
rect 8680 6245 8708 6276
rect 10226 6264 10232 6276
rect 10284 6264 10290 6316
rect 10318 6264 10324 6316
rect 10376 6304 10382 6316
rect 11054 6304 11060 6316
rect 10376 6276 11060 6304
rect 10376 6264 10382 6276
rect 11054 6264 11060 6276
rect 11112 6264 11118 6316
rect 8527 6208 8616 6236
rect 8665 6239 8723 6245
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 8665 6205 8677 6239
rect 8711 6205 8723 6239
rect 8665 6199 8723 6205
rect 8849 6239 8907 6245
rect 8849 6205 8861 6239
rect 8895 6236 8907 6239
rect 9677 6239 9735 6245
rect 9677 6236 9689 6239
rect 8895 6208 9689 6236
rect 8895 6205 8907 6208
rect 8849 6199 8907 6205
rect 9677 6205 9689 6208
rect 9723 6236 9735 6239
rect 9950 6236 9956 6248
rect 9723 6208 9956 6236
rect 9723 6205 9735 6208
rect 9677 6199 9735 6205
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 10042 6196 10048 6248
rect 10100 6236 10106 6248
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 10100 6208 10425 6236
rect 10100 6196 10106 6208
rect 10413 6205 10425 6208
rect 10459 6236 10471 6239
rect 10962 6236 10968 6248
rect 10459 6208 10968 6236
rect 10459 6205 10471 6208
rect 10413 6199 10471 6205
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 11330 6196 11336 6248
rect 11388 6196 11394 6248
rect 11624 6245 11652 6344
rect 12406 6344 19984 6372
rect 11425 6239 11483 6245
rect 11425 6205 11437 6239
rect 11471 6205 11483 6239
rect 11425 6199 11483 6205
rect 11609 6239 11667 6245
rect 11609 6205 11621 6239
rect 11655 6236 11667 6239
rect 12406 6236 12434 6344
rect 19978 6332 19984 6344
rect 20036 6332 20042 6384
rect 16390 6304 16396 6316
rect 13924 6276 16396 6304
rect 11655 6208 12434 6236
rect 13725 6239 13783 6245
rect 11655 6205 11667 6208
rect 11609 6199 11667 6205
rect 13725 6205 13737 6239
rect 13771 6236 13783 6239
rect 13814 6236 13820 6248
rect 13771 6208 13820 6236
rect 13771 6205 13783 6208
rect 13725 6199 13783 6205
rect 6816 6171 6874 6177
rect 6816 6137 6828 6171
rect 6862 6168 6874 6171
rect 8113 6171 8171 6177
rect 8113 6168 8125 6171
rect 6862 6140 8125 6168
rect 6862 6137 6874 6140
rect 6816 6131 6874 6137
rect 8113 6137 8125 6140
rect 8159 6137 8171 6171
rect 9968 6168 9996 6196
rect 10597 6171 10655 6177
rect 10597 6168 10609 6171
rect 8113 6131 8171 6137
rect 8496 6140 9536 6168
rect 9968 6140 10609 6168
rect 5399 6072 6224 6100
rect 7929 6103 7987 6109
rect 5399 6069 5411 6072
rect 5353 6063 5411 6069
rect 7929 6069 7941 6103
rect 7975 6100 7987 6103
rect 8496 6100 8524 6140
rect 9508 6112 9536 6140
rect 10597 6137 10609 6140
rect 10643 6137 10655 6171
rect 10597 6131 10655 6137
rect 10689 6171 10747 6177
rect 10689 6137 10701 6171
rect 10735 6168 10747 6171
rect 11057 6171 11115 6177
rect 10735 6140 10916 6168
rect 10735 6137 10747 6140
rect 10689 6131 10747 6137
rect 7975 6072 8524 6100
rect 7975 6069 7987 6072
rect 7929 6063 7987 6069
rect 8570 6060 8576 6112
rect 8628 6060 8634 6112
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 10704 6100 10732 6131
rect 9548 6072 10732 6100
rect 9548 6060 9554 6072
rect 10778 6060 10784 6112
rect 10836 6060 10842 6112
rect 10888 6100 10916 6140
rect 11057 6137 11069 6171
rect 11103 6168 11115 6171
rect 11440 6168 11468 6199
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 13924 6177 13952 6276
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 17586 6264 17592 6316
rect 17644 6304 17650 6316
rect 18138 6304 18144 6316
rect 17644 6276 18144 6304
rect 17644 6264 17650 6276
rect 18138 6264 18144 6276
rect 18196 6304 18202 6316
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 18196 6276 18705 6304
rect 18196 6264 18202 6276
rect 18693 6273 18705 6276
rect 18739 6273 18751 6307
rect 19996 6304 20024 6332
rect 20640 6313 20668 6412
rect 21266 6400 21272 6412
rect 21324 6440 21330 6452
rect 21324 6412 23428 6440
rect 21324 6400 21330 6412
rect 20717 6375 20775 6381
rect 20717 6341 20729 6375
rect 20763 6372 20775 6375
rect 20898 6372 20904 6384
rect 20763 6344 20904 6372
rect 20763 6341 20775 6344
rect 20717 6335 20775 6341
rect 20898 6332 20904 6344
rect 20956 6332 20962 6384
rect 23400 6316 23428 6412
rect 23474 6400 23480 6452
rect 23532 6400 23538 6452
rect 23569 6443 23627 6449
rect 23569 6409 23581 6443
rect 23615 6440 23627 6443
rect 23750 6440 23756 6452
rect 23615 6412 23756 6440
rect 23615 6409 23627 6412
rect 23569 6403 23627 6409
rect 23750 6400 23756 6412
rect 23808 6440 23814 6452
rect 24121 6443 24179 6449
rect 24121 6440 24133 6443
rect 23808 6412 24133 6440
rect 23808 6400 23814 6412
rect 24121 6409 24133 6412
rect 24167 6409 24179 6443
rect 24121 6403 24179 6409
rect 25222 6400 25228 6452
rect 25280 6440 25286 6452
rect 25866 6440 25872 6452
rect 25280 6412 25872 6440
rect 25280 6400 25286 6412
rect 25866 6400 25872 6412
rect 25924 6400 25930 6452
rect 20625 6307 20683 6313
rect 19996 6276 20576 6304
rect 18693 6267 18751 6273
rect 14093 6239 14151 6245
rect 14093 6205 14105 6239
rect 14139 6236 14151 6239
rect 14274 6236 14280 6248
rect 14139 6208 14280 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 14274 6196 14280 6208
rect 14332 6196 14338 6248
rect 16117 6239 16175 6245
rect 16117 6205 16129 6239
rect 16163 6236 16175 6239
rect 16942 6236 16948 6248
rect 16163 6208 16948 6236
rect 16163 6205 16175 6208
rect 16117 6199 16175 6205
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 18046 6196 18052 6248
rect 18104 6196 18110 6248
rect 18322 6236 18328 6248
rect 18156 6208 18328 6236
rect 13909 6171 13967 6177
rect 13909 6168 13921 6171
rect 11103 6140 11468 6168
rect 11624 6140 13921 6168
rect 11103 6137 11115 6140
rect 11057 6131 11115 6137
rect 11624 6112 11652 6140
rect 13909 6137 13921 6140
rect 13955 6137 13967 6171
rect 13909 6131 13967 6137
rect 14001 6171 14059 6177
rect 14001 6137 14013 6171
rect 14047 6137 14059 6171
rect 14001 6131 14059 6137
rect 11422 6100 11428 6112
rect 10888 6072 11428 6100
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 11514 6060 11520 6112
rect 11572 6060 11578 6112
rect 11606 6060 11612 6112
rect 11664 6060 11670 6112
rect 12250 6060 12256 6112
rect 12308 6100 12314 6112
rect 14016 6100 14044 6131
rect 15654 6128 15660 6180
rect 15712 6168 15718 6180
rect 15712 6140 15976 6168
rect 15712 6128 15718 6140
rect 12308 6072 14044 6100
rect 14277 6103 14335 6109
rect 12308 6060 12314 6072
rect 14277 6069 14289 6103
rect 14323 6100 14335 6103
rect 15838 6100 15844 6112
rect 14323 6072 15844 6100
rect 14323 6069 14335 6072
rect 14277 6063 14335 6069
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 15948 6109 15976 6140
rect 16850 6128 16856 6180
rect 16908 6168 16914 6180
rect 17497 6171 17555 6177
rect 17497 6168 17509 6171
rect 16908 6140 17509 6168
rect 16908 6128 16914 6140
rect 17497 6137 17509 6140
rect 17543 6137 17555 6171
rect 17497 6131 17555 6137
rect 17713 6171 17771 6177
rect 17713 6137 17725 6171
rect 17759 6168 17771 6171
rect 18064 6168 18092 6196
rect 18156 6177 18184 6208
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 18414 6196 18420 6248
rect 18472 6196 18478 6248
rect 18509 6239 18567 6245
rect 18509 6205 18521 6239
rect 18555 6236 18567 6239
rect 18598 6236 18604 6248
rect 18555 6208 18604 6236
rect 18555 6205 18567 6208
rect 18509 6199 18567 6205
rect 18598 6196 18604 6208
rect 18656 6196 18662 6248
rect 20438 6196 20444 6248
rect 20496 6196 20502 6248
rect 20548 6236 20576 6276
rect 20625 6273 20637 6307
rect 20671 6273 20683 6307
rect 21266 6304 21272 6316
rect 20625 6267 20683 6273
rect 20824 6276 21272 6304
rect 20824 6248 20852 6276
rect 21266 6264 21272 6276
rect 21324 6264 21330 6316
rect 23382 6264 23388 6316
rect 23440 6264 23446 6316
rect 24486 6304 24492 6316
rect 23492 6276 24492 6304
rect 23492 6248 23520 6276
rect 24486 6264 24492 6276
rect 24544 6264 24550 6316
rect 20806 6236 20812 6248
rect 20548 6208 20812 6236
rect 20806 6196 20812 6208
rect 20864 6196 20870 6248
rect 20901 6239 20959 6245
rect 20901 6205 20913 6239
rect 20947 6236 20959 6239
rect 21358 6236 21364 6248
rect 20947 6208 21364 6236
rect 20947 6205 20959 6208
rect 20901 6199 20959 6205
rect 21358 6196 21364 6208
rect 21416 6196 21422 6248
rect 21818 6196 21824 6248
rect 21876 6236 21882 6248
rect 22370 6236 22376 6248
rect 21876 6208 22376 6236
rect 21876 6196 21882 6208
rect 22370 6196 22376 6208
rect 22428 6236 22434 6248
rect 23474 6236 23480 6248
rect 22428 6208 23480 6236
rect 22428 6196 22434 6208
rect 23474 6196 23480 6208
rect 23532 6196 23538 6248
rect 23658 6196 23664 6248
rect 23716 6196 23722 6248
rect 24029 6239 24087 6245
rect 24029 6236 24041 6239
rect 23768 6208 24041 6236
rect 17759 6140 18092 6168
rect 18141 6171 18199 6177
rect 17759 6137 17771 6140
rect 17713 6131 17771 6137
rect 18141 6137 18153 6171
rect 18187 6137 18199 6171
rect 18141 6131 18199 6137
rect 18233 6171 18291 6177
rect 18233 6137 18245 6171
rect 18279 6168 18291 6171
rect 21082 6168 21088 6180
rect 18279 6140 21088 6168
rect 18279 6137 18291 6140
rect 18233 6131 18291 6137
rect 21082 6128 21088 6140
rect 21140 6128 21146 6180
rect 21266 6128 21272 6180
rect 21324 6168 21330 6180
rect 22002 6168 22008 6180
rect 21324 6140 22008 6168
rect 21324 6128 21330 6140
rect 22002 6128 22008 6140
rect 22060 6128 22066 6180
rect 22128 6171 22186 6177
rect 22128 6137 22140 6171
rect 22174 6168 22186 6171
rect 22738 6168 22744 6180
rect 22174 6140 22744 6168
rect 22174 6137 22186 6140
rect 22128 6131 22186 6137
rect 22738 6128 22744 6140
rect 22796 6128 22802 6180
rect 22830 6128 22836 6180
rect 22888 6168 22894 6180
rect 23768 6168 23796 6208
rect 24029 6205 24041 6208
rect 24075 6205 24087 6239
rect 24029 6199 24087 6205
rect 24302 6196 24308 6248
rect 24360 6196 24366 6248
rect 22888 6140 23796 6168
rect 23937 6171 23995 6177
rect 22888 6128 22894 6140
rect 23937 6137 23949 6171
rect 23983 6168 23995 6171
rect 24210 6168 24216 6180
rect 23983 6140 24216 6168
rect 23983 6137 23995 6140
rect 23937 6131 23995 6137
rect 24210 6128 24216 6140
rect 24268 6128 24274 6180
rect 24397 6171 24455 6177
rect 24397 6137 24409 6171
rect 24443 6168 24455 6171
rect 24578 6168 24584 6180
rect 24443 6140 24584 6168
rect 24443 6137 24455 6140
rect 24397 6131 24455 6137
rect 24578 6128 24584 6140
rect 24636 6128 24642 6180
rect 24762 6177 24768 6180
rect 24756 6131 24768 6177
rect 24762 6128 24768 6131
rect 24820 6128 24826 6180
rect 15933 6103 15991 6109
rect 15933 6069 15945 6103
rect 15979 6069 15991 6103
rect 15933 6063 15991 6069
rect 17865 6103 17923 6109
rect 17865 6069 17877 6103
rect 17911 6100 17923 6103
rect 17954 6100 17960 6112
rect 17911 6072 17960 6100
rect 17911 6069 17923 6072
rect 17865 6063 17923 6069
rect 17954 6060 17960 6072
rect 18012 6060 18018 6112
rect 20622 6060 20628 6112
rect 20680 6100 20686 6112
rect 20993 6103 21051 6109
rect 20993 6100 21005 6103
rect 20680 6072 21005 6100
rect 20680 6060 20686 6072
rect 20993 6069 21005 6072
rect 21039 6100 21051 6103
rect 22554 6100 22560 6112
rect 21039 6072 22560 6100
rect 21039 6069 21051 6072
rect 20993 6063 21051 6069
rect 22554 6060 22560 6072
rect 22612 6060 22618 6112
rect 552 6010 27576 6032
rect 552 5958 7114 6010
rect 7166 5958 7178 6010
rect 7230 5958 7242 6010
rect 7294 5958 7306 6010
rect 7358 5958 7370 6010
rect 7422 5958 13830 6010
rect 13882 5958 13894 6010
rect 13946 5958 13958 6010
rect 14010 5958 14022 6010
rect 14074 5958 14086 6010
rect 14138 5958 20546 6010
rect 20598 5958 20610 6010
rect 20662 5958 20674 6010
rect 20726 5958 20738 6010
rect 20790 5958 20802 6010
rect 20854 5958 27262 6010
rect 27314 5958 27326 6010
rect 27378 5958 27390 6010
rect 27442 5958 27454 6010
rect 27506 5958 27518 6010
rect 27570 5958 27576 6010
rect 552 5936 27576 5958
rect 4338 5896 4344 5908
rect 4080 5868 4344 5896
rect 4080 5769 4108 5868
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 5718 5856 5724 5908
rect 5776 5896 5782 5908
rect 5813 5899 5871 5905
rect 5813 5896 5825 5899
rect 5776 5868 5825 5896
rect 5776 5856 5782 5868
rect 5813 5865 5825 5868
rect 5859 5865 5871 5899
rect 5813 5859 5871 5865
rect 7742 5856 7748 5908
rect 7800 5856 7806 5908
rect 9493 5899 9551 5905
rect 9493 5865 9505 5899
rect 9539 5896 9551 5899
rect 9674 5896 9680 5908
rect 9539 5868 9680 5896
rect 9539 5865 9551 5868
rect 9493 5859 9551 5865
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 11609 5899 11667 5905
rect 11609 5896 11621 5899
rect 11388 5868 11621 5896
rect 11388 5856 11394 5868
rect 11609 5865 11621 5868
rect 11655 5865 11667 5899
rect 11609 5859 11667 5865
rect 12069 5899 12127 5905
rect 12069 5865 12081 5899
rect 12115 5896 12127 5899
rect 12158 5896 12164 5908
rect 12115 5868 12164 5896
rect 12115 5865 12127 5868
rect 12069 5859 12127 5865
rect 12158 5856 12164 5868
rect 12216 5856 12222 5908
rect 12250 5856 12256 5908
rect 12308 5856 12314 5908
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 13081 5899 13139 5905
rect 13081 5896 13093 5899
rect 13044 5868 13093 5896
rect 13044 5856 13050 5868
rect 13081 5865 13093 5868
rect 13127 5865 13139 5899
rect 13081 5859 13139 5865
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 13909 5899 13967 5905
rect 13909 5896 13921 5899
rect 13872 5868 13921 5896
rect 13872 5856 13878 5868
rect 13909 5865 13921 5868
rect 13955 5865 13967 5899
rect 13909 5859 13967 5865
rect 14182 5856 14188 5908
rect 14240 5896 14246 5908
rect 14737 5899 14795 5905
rect 14737 5896 14749 5899
rect 14240 5868 14749 5896
rect 14240 5856 14246 5868
rect 14737 5865 14749 5868
rect 14783 5865 14795 5899
rect 14737 5859 14795 5865
rect 15102 5856 15108 5908
rect 15160 5896 15166 5908
rect 16114 5896 16120 5908
rect 15160 5868 16120 5896
rect 15160 5856 15166 5868
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 17678 5856 17684 5908
rect 17736 5896 17742 5908
rect 19245 5899 19303 5905
rect 19245 5896 19257 5899
rect 17736 5868 19257 5896
rect 17736 5856 17742 5868
rect 19245 5865 19257 5868
rect 19291 5865 19303 5899
rect 19886 5896 19892 5908
rect 19245 5859 19303 5865
rect 19628 5868 19892 5896
rect 6730 5828 6736 5840
rect 4172 5800 6736 5828
rect 4172 5769 4200 5800
rect 6730 5788 6736 5800
rect 6788 5788 6794 5840
rect 8202 5788 8208 5840
rect 8260 5828 8266 5840
rect 8573 5831 8631 5837
rect 8573 5828 8585 5831
rect 8260 5800 8585 5828
rect 8260 5788 8266 5800
rect 8573 5797 8585 5800
rect 8619 5828 8631 5831
rect 10134 5828 10140 5840
rect 8619 5800 10140 5828
rect 8619 5797 8631 5800
rect 8573 5791 8631 5797
rect 10134 5788 10140 5800
rect 10192 5788 10198 5840
rect 10781 5831 10839 5837
rect 10781 5797 10793 5831
rect 10827 5828 10839 5831
rect 10870 5828 10876 5840
rect 10827 5800 10876 5828
rect 10827 5797 10839 5800
rect 10781 5791 10839 5797
rect 10870 5788 10876 5800
rect 10928 5788 10934 5840
rect 12526 5828 12532 5840
rect 11900 5800 12532 5828
rect 3973 5763 4031 5769
rect 3973 5729 3985 5763
rect 4019 5729 4031 5763
rect 3973 5723 4031 5729
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 4157 5763 4215 5769
rect 4157 5729 4169 5763
rect 4203 5729 4215 5763
rect 4157 5723 4215 5729
rect 3988 5692 4016 5723
rect 4246 5720 4252 5772
rect 4304 5760 4310 5772
rect 4341 5763 4399 5769
rect 4341 5760 4353 5763
rect 4304 5732 4353 5760
rect 4304 5720 4310 5732
rect 4341 5729 4353 5732
rect 4387 5760 4399 5763
rect 5166 5760 5172 5772
rect 4387 5732 5172 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 5258 5720 5264 5772
rect 5316 5760 5322 5772
rect 5353 5763 5411 5769
rect 5353 5760 5365 5763
rect 5316 5732 5365 5760
rect 5316 5720 5322 5732
rect 5353 5729 5365 5732
rect 5399 5760 5411 5763
rect 5442 5760 5448 5772
rect 5399 5732 5448 5760
rect 5399 5729 5411 5732
rect 5353 5723 5411 5729
rect 5442 5720 5448 5732
rect 5500 5720 5506 5772
rect 5994 5720 6000 5772
rect 6052 5720 6058 5772
rect 7469 5763 7527 5769
rect 7469 5729 7481 5763
rect 7515 5760 7527 5763
rect 7837 5763 7895 5769
rect 7837 5760 7849 5763
rect 7515 5732 7849 5760
rect 7515 5729 7527 5732
rect 7469 5723 7527 5729
rect 7837 5729 7849 5732
rect 7883 5729 7895 5763
rect 8757 5763 8815 5769
rect 8757 5760 8769 5763
rect 7837 5723 7895 5729
rect 7944 5732 8769 5760
rect 4433 5695 4491 5701
rect 4433 5692 4445 5695
rect 3988 5664 4445 5692
rect 4433 5661 4445 5664
rect 4479 5661 4491 5695
rect 4433 5655 4491 5661
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 4985 5695 5043 5701
rect 4985 5692 4997 5695
rect 4580 5664 4997 5692
rect 4580 5652 4586 5664
rect 4985 5661 4997 5664
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 5074 5652 5080 5704
rect 5132 5692 5138 5704
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 5132 5664 7573 5692
rect 5132 5652 5138 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 7561 5655 7619 5661
rect 5350 5584 5356 5636
rect 5408 5624 5414 5636
rect 7576 5624 7604 5655
rect 7742 5652 7748 5704
rect 7800 5652 7806 5704
rect 7944 5624 7972 5732
rect 8757 5729 8769 5732
rect 8803 5760 8815 5763
rect 8846 5760 8852 5772
rect 8803 5732 8852 5760
rect 8803 5729 8815 5732
rect 8757 5723 8815 5729
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5760 8999 5763
rect 9490 5760 9496 5772
rect 8987 5732 9496 5760
rect 8987 5729 8999 5732
rect 8941 5723 8999 5729
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8956 5692 8984 5723
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 10962 5720 10968 5772
rect 11020 5720 11026 5772
rect 11900 5769 11928 5800
rect 12526 5788 12532 5800
rect 12584 5788 12590 5840
rect 13354 5788 13360 5840
rect 13412 5828 13418 5840
rect 15010 5828 15016 5840
rect 13412 5800 15016 5828
rect 13412 5788 13418 5800
rect 15010 5788 15016 5800
rect 15068 5788 15074 5840
rect 18414 5788 18420 5840
rect 18472 5828 18478 5840
rect 19628 5837 19656 5868
rect 19886 5856 19892 5868
rect 19944 5896 19950 5908
rect 20257 5899 20315 5905
rect 20257 5896 20269 5899
rect 19944 5868 20269 5896
rect 19944 5856 19950 5868
rect 20257 5865 20269 5868
rect 20303 5896 20315 5899
rect 20346 5896 20352 5908
rect 20303 5868 20352 5896
rect 20303 5865 20315 5868
rect 20257 5859 20315 5865
rect 20346 5856 20352 5868
rect 20404 5856 20410 5908
rect 21174 5896 21180 5908
rect 20456 5868 21180 5896
rect 19613 5831 19671 5837
rect 19613 5828 19625 5831
rect 18472 5800 19625 5828
rect 18472 5788 18478 5800
rect 19613 5797 19625 5800
rect 19659 5797 19671 5831
rect 20456 5828 20484 5868
rect 21174 5856 21180 5868
rect 21232 5856 21238 5908
rect 21358 5856 21364 5908
rect 21416 5856 21422 5908
rect 22097 5899 22155 5905
rect 22097 5865 22109 5899
rect 22143 5865 22155 5899
rect 22097 5859 22155 5865
rect 19613 5791 19671 5797
rect 19904 5800 20484 5828
rect 20717 5831 20775 5837
rect 11885 5763 11943 5769
rect 11885 5729 11897 5763
rect 11931 5729 11943 5763
rect 11885 5723 11943 5729
rect 12161 5763 12219 5769
rect 12161 5729 12173 5763
rect 12207 5760 12219 5763
rect 12621 5763 12679 5769
rect 12207 5732 12434 5760
rect 12207 5729 12219 5732
rect 12161 5723 12219 5729
rect 8527 5664 8984 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 9030 5652 9036 5704
rect 9088 5692 9094 5704
rect 9088 5664 11836 5692
rect 9088 5652 9094 5664
rect 5408 5596 5672 5624
rect 7576 5596 7972 5624
rect 5408 5584 5414 5596
rect 3326 5516 3332 5568
rect 3384 5556 3390 5568
rect 3697 5559 3755 5565
rect 3697 5556 3709 5559
rect 3384 5528 3709 5556
rect 3384 5516 3390 5528
rect 3697 5525 3709 5528
rect 3743 5525 3755 5559
rect 3697 5519 3755 5525
rect 5534 5516 5540 5568
rect 5592 5516 5598 5568
rect 5644 5556 5672 5596
rect 8846 5584 8852 5636
rect 8904 5624 8910 5636
rect 10778 5624 10784 5636
rect 8904 5596 10784 5624
rect 8904 5584 8910 5596
rect 10778 5584 10784 5596
rect 10836 5584 10842 5636
rect 11606 5556 11612 5568
rect 5644 5528 11612 5556
rect 11606 5516 11612 5528
rect 11664 5516 11670 5568
rect 11698 5516 11704 5568
rect 11756 5516 11762 5568
rect 11808 5556 11836 5664
rect 12406 5624 12434 5732
rect 12621 5729 12633 5763
rect 12667 5760 12679 5763
rect 12802 5760 12808 5772
rect 12667 5732 12808 5760
rect 12667 5729 12679 5732
rect 12621 5723 12679 5729
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 13446 5720 13452 5772
rect 13504 5720 13510 5772
rect 13541 5763 13599 5769
rect 13541 5729 13553 5763
rect 13587 5760 13599 5763
rect 14182 5760 14188 5772
rect 13587 5732 14188 5760
rect 13587 5729 13599 5732
rect 13541 5723 13599 5729
rect 14182 5720 14188 5732
rect 14240 5720 14246 5772
rect 14277 5763 14335 5769
rect 14277 5729 14289 5763
rect 14323 5760 14335 5763
rect 14550 5760 14556 5772
rect 14323 5732 14556 5760
rect 14323 5729 14335 5732
rect 14277 5723 14335 5729
rect 14550 5720 14556 5732
rect 14608 5760 14614 5772
rect 15378 5760 15384 5772
rect 14608 5732 15384 5760
rect 14608 5720 14614 5732
rect 15378 5720 15384 5732
rect 15436 5720 15442 5772
rect 15838 5720 15844 5772
rect 15896 5760 15902 5772
rect 18046 5769 18052 5772
rect 16301 5763 16359 5769
rect 16301 5760 16313 5763
rect 15896 5732 16313 5760
rect 15896 5720 15902 5732
rect 16301 5729 16313 5732
rect 16347 5729 16359 5763
rect 16301 5723 16359 5729
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5760 16543 5763
rect 16577 5763 16635 5769
rect 16577 5760 16589 5763
rect 16531 5732 16589 5760
rect 16531 5729 16543 5732
rect 16485 5723 16543 5729
rect 16577 5729 16589 5732
rect 16623 5729 16635 5763
rect 16577 5723 16635 5729
rect 18040 5723 18052 5769
rect 18046 5720 18052 5723
rect 18104 5720 18110 5772
rect 19429 5763 19487 5769
rect 19429 5729 19441 5763
rect 19475 5760 19487 5763
rect 19518 5760 19524 5772
rect 19475 5732 19524 5760
rect 19475 5729 19487 5732
rect 19429 5723 19487 5729
rect 12710 5652 12716 5704
rect 12768 5652 12774 5704
rect 12897 5695 12955 5701
rect 12897 5661 12909 5695
rect 12943 5692 12955 5695
rect 12986 5692 12992 5704
rect 12943 5664 12992 5692
rect 12943 5661 12955 5664
rect 12897 5655 12955 5661
rect 12912 5624 12940 5655
rect 12986 5652 12992 5664
rect 13044 5692 13050 5704
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13044 5664 13737 5692
rect 13044 5652 13050 5664
rect 13725 5661 13737 5664
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 12406 5596 12940 5624
rect 13740 5624 13768 5655
rect 14366 5652 14372 5704
rect 14424 5652 14430 5704
rect 14461 5695 14519 5701
rect 14461 5661 14473 5695
rect 14507 5661 14519 5695
rect 14461 5655 14519 5661
rect 14476 5624 14504 5655
rect 15194 5652 15200 5704
rect 15252 5652 15258 5704
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5692 15347 5695
rect 15654 5692 15660 5704
rect 15335 5664 15660 5692
rect 15335 5661 15347 5664
rect 15289 5655 15347 5661
rect 15304 5624 15332 5655
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5692 16175 5695
rect 16850 5692 16856 5704
rect 16163 5664 16856 5692
rect 16163 5661 16175 5664
rect 16117 5655 16175 5661
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 13740 5596 15332 5624
rect 14274 5556 14280 5568
rect 11808 5528 14280 5556
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 16761 5559 16819 5565
rect 16761 5525 16773 5559
rect 16807 5556 16819 5559
rect 16850 5556 16856 5568
rect 16807 5528 16856 5556
rect 16807 5525 16819 5528
rect 16761 5519 16819 5525
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 17788 5556 17816 5655
rect 19153 5627 19211 5633
rect 19153 5593 19165 5627
rect 19199 5624 19211 5627
rect 19444 5624 19472 5723
rect 19518 5720 19524 5732
rect 19576 5720 19582 5772
rect 19904 5769 19932 5800
rect 20717 5797 20729 5831
rect 20763 5828 20775 5831
rect 22112 5828 22140 5859
rect 22738 5856 22744 5908
rect 22796 5856 22802 5908
rect 24762 5856 24768 5908
rect 24820 5896 24826 5908
rect 25041 5899 25099 5905
rect 25041 5896 25053 5899
rect 24820 5868 25053 5896
rect 24820 5856 24826 5868
rect 25041 5865 25053 5868
rect 25087 5865 25099 5899
rect 25041 5859 25099 5865
rect 25130 5856 25136 5908
rect 25188 5896 25194 5908
rect 25188 5868 25820 5896
rect 25188 5856 25194 5868
rect 20763 5800 22140 5828
rect 20763 5797 20775 5800
rect 20717 5791 20775 5797
rect 24578 5788 24584 5840
rect 24636 5828 24642 5840
rect 25685 5831 25743 5837
rect 25685 5828 25697 5831
rect 24636 5800 25697 5828
rect 24636 5788 24642 5800
rect 25685 5797 25697 5800
rect 25731 5797 25743 5831
rect 25685 5791 25743 5797
rect 19889 5763 19947 5769
rect 19889 5729 19901 5763
rect 19935 5729 19947 5763
rect 19889 5723 19947 5729
rect 19978 5720 19984 5772
rect 20036 5760 20042 5772
rect 20073 5763 20131 5769
rect 20073 5760 20085 5763
rect 20036 5732 20085 5760
rect 20036 5720 20042 5732
rect 20073 5729 20085 5732
rect 20119 5729 20131 5763
rect 20073 5723 20131 5729
rect 20254 5720 20260 5772
rect 20312 5760 20318 5772
rect 20349 5763 20407 5769
rect 20349 5760 20361 5763
rect 20312 5732 20361 5760
rect 20312 5720 20318 5732
rect 20349 5729 20361 5732
rect 20395 5729 20407 5763
rect 22925 5763 22983 5769
rect 22925 5760 22937 5763
rect 20349 5723 20407 5729
rect 20916 5732 22937 5760
rect 20916 5633 20944 5732
rect 22925 5729 22937 5732
rect 22971 5729 22983 5763
rect 22925 5723 22983 5729
rect 23566 5720 23572 5772
rect 23624 5760 23630 5772
rect 24121 5763 24179 5769
rect 24121 5760 24133 5763
rect 23624 5732 24133 5760
rect 23624 5720 23630 5732
rect 24121 5729 24133 5732
rect 24167 5729 24179 5763
rect 24121 5723 24179 5729
rect 24210 5720 24216 5772
rect 24268 5760 24274 5772
rect 24397 5763 24455 5769
rect 24397 5760 24409 5763
rect 24268 5732 24409 5760
rect 24268 5720 24274 5732
rect 24397 5729 24409 5732
rect 24443 5729 24455 5763
rect 24397 5723 24455 5729
rect 25130 5720 25136 5772
rect 25188 5760 25194 5772
rect 25792 5769 25820 5868
rect 25317 5763 25375 5769
rect 25317 5760 25329 5763
rect 25188 5732 25329 5760
rect 25188 5720 25194 5732
rect 25317 5729 25329 5732
rect 25363 5729 25375 5763
rect 25317 5723 25375 5729
rect 25501 5763 25559 5769
rect 25501 5729 25513 5763
rect 25547 5760 25559 5763
rect 25593 5763 25651 5769
rect 25593 5760 25605 5763
rect 25547 5732 25605 5760
rect 25547 5729 25559 5732
rect 25501 5723 25559 5729
rect 25593 5729 25605 5732
rect 25639 5729 25651 5763
rect 25593 5723 25651 5729
rect 25777 5763 25835 5769
rect 25777 5729 25789 5763
rect 25823 5760 25835 5763
rect 26050 5760 26056 5772
rect 25823 5732 26056 5760
rect 25823 5729 25835 5732
rect 25777 5723 25835 5729
rect 21174 5652 21180 5704
rect 21232 5692 21238 5704
rect 21910 5692 21916 5704
rect 21232 5664 21916 5692
rect 21232 5652 21238 5664
rect 21910 5652 21916 5664
rect 21968 5652 21974 5704
rect 22281 5695 22339 5701
rect 22281 5692 22293 5695
rect 22204 5664 22293 5692
rect 19199 5596 19472 5624
rect 20901 5627 20959 5633
rect 19199 5593 19211 5596
rect 19153 5587 19211 5593
rect 20901 5593 20913 5627
rect 20947 5593 20959 5627
rect 20901 5587 20959 5593
rect 20990 5584 20996 5636
rect 21048 5624 21054 5636
rect 22204 5624 22232 5664
rect 22281 5661 22293 5664
rect 22327 5661 22339 5695
rect 22281 5655 22339 5661
rect 22370 5652 22376 5704
rect 22428 5652 22434 5704
rect 22465 5695 22523 5701
rect 22465 5661 22477 5695
rect 22511 5661 22523 5695
rect 22465 5655 22523 5661
rect 21048 5596 22232 5624
rect 21048 5584 21054 5596
rect 18138 5556 18144 5568
rect 17788 5528 18144 5556
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 20717 5559 20775 5565
rect 20717 5525 20729 5559
rect 20763 5556 20775 5559
rect 21450 5556 21456 5568
rect 20763 5528 21456 5556
rect 20763 5525 20775 5528
rect 20717 5519 20775 5525
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 22094 5516 22100 5568
rect 22152 5556 22158 5568
rect 22480 5556 22508 5655
rect 22554 5652 22560 5704
rect 22612 5652 22618 5704
rect 23937 5695 23995 5701
rect 23937 5661 23949 5695
rect 23983 5661 23995 5695
rect 25516 5692 25544 5723
rect 26050 5720 26056 5732
rect 26108 5720 26114 5772
rect 23937 5655 23995 5661
rect 24320 5664 25544 5692
rect 23952 5624 23980 5655
rect 24210 5624 24216 5636
rect 23952 5596 24216 5624
rect 24210 5584 24216 5596
rect 24268 5584 24274 5636
rect 22152 5528 22508 5556
rect 22152 5516 22158 5528
rect 23750 5516 23756 5568
rect 23808 5556 23814 5568
rect 24320 5565 24348 5664
rect 24305 5559 24363 5565
rect 24305 5556 24317 5559
rect 23808 5528 24317 5556
rect 23808 5516 23814 5528
rect 24305 5525 24317 5528
rect 24351 5525 24363 5559
rect 24305 5519 24363 5525
rect 25130 5516 25136 5568
rect 25188 5516 25194 5568
rect 552 5466 27416 5488
rect 552 5414 3756 5466
rect 3808 5414 3820 5466
rect 3872 5414 3884 5466
rect 3936 5414 3948 5466
rect 4000 5414 4012 5466
rect 4064 5414 10472 5466
rect 10524 5414 10536 5466
rect 10588 5414 10600 5466
rect 10652 5414 10664 5466
rect 10716 5414 10728 5466
rect 10780 5414 17188 5466
rect 17240 5414 17252 5466
rect 17304 5414 17316 5466
rect 17368 5414 17380 5466
rect 17432 5414 17444 5466
rect 17496 5414 23904 5466
rect 23956 5414 23968 5466
rect 24020 5414 24032 5466
rect 24084 5414 24096 5466
rect 24148 5414 24160 5466
rect 24212 5414 27416 5466
rect 552 5392 27416 5414
rect 6730 5312 6736 5364
rect 6788 5352 6794 5364
rect 7009 5355 7067 5361
rect 7009 5352 7021 5355
rect 6788 5324 7021 5352
rect 6788 5312 6794 5324
rect 7009 5321 7021 5324
rect 7055 5321 7067 5355
rect 8662 5352 8668 5364
rect 7009 5315 7067 5321
rect 7392 5324 8668 5352
rect 4154 5176 4160 5228
rect 4212 5176 4218 5228
rect 5166 5176 5172 5228
rect 5224 5216 5230 5228
rect 5224 5188 7328 5216
rect 5224 5176 5230 5188
rect 6181 5151 6239 5157
rect 6181 5148 6193 5151
rect 5552 5120 6193 5148
rect 4424 5083 4482 5089
rect 4424 5049 4436 5083
rect 4470 5080 4482 5083
rect 4706 5080 4712 5092
rect 4470 5052 4712 5080
rect 4470 5049 4482 5052
rect 4424 5043 4482 5049
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 5552 5024 5580 5120
rect 6181 5117 6193 5120
rect 6227 5117 6239 5151
rect 6181 5111 6239 5117
rect 6362 5108 6368 5160
rect 6420 5148 6426 5160
rect 7193 5151 7251 5157
rect 7193 5148 7205 5151
rect 6420 5120 7205 5148
rect 6420 5108 6426 5120
rect 7193 5117 7205 5120
rect 7239 5117 7251 5151
rect 7193 5111 7251 5117
rect 5534 4972 5540 5024
rect 5592 4972 5598 5024
rect 5626 4972 5632 5024
rect 5684 4972 5690 5024
rect 7208 5012 7236 5111
rect 7300 5080 7328 5188
rect 7392 5157 7420 5324
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 9950 5352 9956 5364
rect 9907 5324 9956 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 10042 5312 10048 5364
rect 10100 5312 10106 5364
rect 12894 5312 12900 5364
rect 12952 5352 12958 5364
rect 13541 5355 13599 5361
rect 13541 5352 13553 5355
rect 12952 5324 13553 5352
rect 12952 5312 12958 5324
rect 13541 5321 13553 5324
rect 13587 5321 13599 5355
rect 13541 5315 13599 5321
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 14553 5355 14611 5361
rect 14553 5352 14565 5355
rect 13780 5324 14565 5352
rect 13780 5312 13786 5324
rect 14553 5321 14565 5324
rect 14599 5321 14611 5355
rect 14553 5315 14611 5321
rect 15105 5355 15163 5361
rect 15105 5321 15117 5355
rect 15151 5352 15163 5355
rect 15746 5352 15752 5364
rect 15151 5324 15752 5352
rect 15151 5321 15163 5324
rect 15105 5315 15163 5321
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 16592 5324 17540 5352
rect 16206 5284 16212 5296
rect 11813 5256 16212 5284
rect 7484 5188 8064 5216
rect 7484 5157 7512 5188
rect 8036 5157 8064 5188
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5117 7435 5151
rect 7377 5111 7435 5117
rect 7469 5151 7527 5157
rect 7469 5117 7481 5151
rect 7515 5117 7527 5151
rect 7469 5111 7527 5117
rect 7745 5151 7803 5157
rect 7745 5117 7757 5151
rect 7791 5117 7803 5151
rect 7745 5111 7803 5117
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5148 8079 5151
rect 8386 5148 8392 5160
rect 8067 5120 8392 5148
rect 8067 5117 8079 5120
rect 8021 5111 8079 5117
rect 7561 5083 7619 5089
rect 7561 5080 7573 5083
rect 7300 5052 7573 5080
rect 7561 5049 7573 5052
rect 7607 5049 7619 5083
rect 7561 5043 7619 5049
rect 7760 5024 7788 5111
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 8481 5151 8539 5157
rect 8481 5117 8493 5151
rect 8527 5148 8539 5151
rect 9122 5148 9128 5160
rect 8527 5120 9128 5148
rect 8527 5117 8539 5120
rect 8481 5111 8539 5117
rect 9122 5108 9128 5120
rect 9180 5148 9186 5160
rect 9674 5148 9680 5160
rect 9180 5120 9680 5148
rect 9180 5108 9186 5120
rect 9674 5108 9680 5120
rect 9732 5148 9738 5160
rect 10870 5148 10876 5160
rect 9732 5120 10876 5148
rect 9732 5108 9738 5120
rect 10870 5108 10876 5120
rect 10928 5148 10934 5160
rect 11425 5151 11483 5157
rect 11425 5148 11437 5151
rect 10928 5120 11437 5148
rect 10928 5108 10934 5120
rect 11425 5117 11437 5120
rect 11471 5117 11483 5151
rect 11425 5111 11483 5117
rect 7929 5083 7987 5089
rect 7929 5049 7941 5083
rect 7975 5080 7987 5083
rect 8294 5080 8300 5092
rect 7975 5052 8300 5080
rect 7975 5049 7987 5052
rect 7929 5043 7987 5049
rect 8294 5040 8300 5052
rect 8352 5040 8358 5092
rect 8570 5040 8576 5092
rect 8628 5080 8634 5092
rect 8726 5083 8784 5089
rect 8726 5080 8738 5083
rect 8628 5052 8738 5080
rect 8628 5040 8634 5052
rect 8726 5049 8738 5052
rect 8772 5049 8784 5083
rect 8726 5043 8784 5049
rect 11180 5083 11238 5089
rect 11180 5049 11192 5083
rect 11226 5080 11238 5083
rect 11514 5080 11520 5092
rect 11226 5052 11520 5080
rect 11226 5049 11238 5052
rect 11180 5043 11238 5049
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 7742 5012 7748 5024
rect 7208 4984 7748 5012
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 8478 4972 8484 5024
rect 8536 5012 8542 5024
rect 9398 5012 9404 5024
rect 8536 4984 9404 5012
rect 8536 4972 8542 4984
rect 9398 4972 9404 4984
rect 9456 5012 9462 5024
rect 11813 5012 11841 5256
rect 14185 5219 14243 5225
rect 14185 5185 14197 5219
rect 14231 5216 14243 5219
rect 15396 5216 15424 5256
rect 16206 5244 16212 5256
rect 16264 5244 16270 5296
rect 14231 5188 15056 5216
rect 15396 5188 15516 5216
rect 14231 5185 14243 5188
rect 14185 5179 14243 5185
rect 15028 5160 15056 5188
rect 12618 5108 12624 5160
rect 12676 5148 12682 5160
rect 12713 5151 12771 5157
rect 12713 5148 12725 5151
rect 12676 5120 12725 5148
rect 12676 5108 12682 5120
rect 12713 5117 12725 5120
rect 12759 5117 12771 5151
rect 12713 5111 12771 5117
rect 14274 5108 14280 5160
rect 14332 5148 14338 5160
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 14332 5120 14381 5148
rect 14332 5108 14338 5120
rect 14369 5117 14381 5120
rect 14415 5117 14427 5151
rect 14369 5111 14427 5117
rect 14458 5108 14464 5160
rect 14516 5108 14522 5160
rect 15010 5108 15016 5160
rect 15068 5148 15074 5160
rect 15488 5157 15516 5188
rect 15654 5176 15660 5228
rect 15712 5176 15718 5228
rect 15473 5151 15531 5157
rect 15068 5120 15424 5148
rect 15068 5108 15074 5120
rect 12986 5040 12992 5092
rect 13044 5080 13050 5092
rect 14001 5083 14059 5089
rect 14001 5080 14013 5083
rect 13044 5052 14013 5080
rect 13044 5040 13050 5052
rect 14001 5049 14013 5052
rect 14047 5049 14059 5083
rect 14476 5080 14504 5108
rect 15396 5080 15424 5120
rect 15473 5117 15485 5151
rect 15519 5117 15531 5151
rect 15473 5111 15531 5117
rect 15565 5151 15623 5157
rect 15565 5117 15577 5151
rect 15611 5148 15623 5151
rect 16022 5148 16028 5160
rect 15611 5120 16028 5148
rect 15611 5117 15623 5120
rect 15565 5111 15623 5117
rect 16022 5108 16028 5120
rect 16080 5108 16086 5160
rect 16592 5157 16620 5324
rect 17512 5284 17540 5324
rect 18046 5312 18052 5364
rect 18104 5352 18110 5364
rect 18233 5355 18291 5361
rect 18233 5352 18245 5355
rect 18104 5324 18245 5352
rect 18104 5312 18110 5324
rect 18233 5321 18245 5324
rect 18279 5321 18291 5355
rect 20806 5352 20812 5364
rect 18233 5315 18291 5321
rect 20364 5324 20812 5352
rect 18138 5284 18144 5296
rect 17512 5256 18144 5284
rect 18138 5244 18144 5256
rect 18196 5244 18202 5296
rect 17954 5176 17960 5228
rect 18012 5216 18018 5228
rect 18012 5188 18460 5216
rect 18012 5176 18018 5188
rect 16850 5157 16856 5160
rect 16577 5151 16635 5157
rect 16577 5117 16589 5151
rect 16623 5117 16635 5151
rect 16844 5148 16856 5157
rect 16811 5120 16856 5148
rect 16577 5111 16635 5117
rect 16844 5111 16856 5120
rect 16850 5108 16856 5111
rect 16908 5108 16914 5160
rect 18432 5157 18460 5188
rect 18417 5151 18475 5157
rect 18417 5117 18429 5151
rect 18463 5117 18475 5151
rect 18417 5111 18475 5117
rect 19886 5108 19892 5160
rect 19944 5108 19950 5160
rect 20073 5151 20131 5157
rect 20073 5117 20085 5151
rect 20119 5148 20131 5151
rect 20364 5148 20392 5324
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 21821 5355 21879 5361
rect 21821 5321 21833 5355
rect 21867 5352 21879 5355
rect 21910 5352 21916 5364
rect 21867 5324 21916 5352
rect 21867 5321 21879 5324
rect 21821 5315 21879 5321
rect 21910 5312 21916 5324
rect 21968 5312 21974 5364
rect 23566 5312 23572 5364
rect 23624 5312 23630 5364
rect 24486 5312 24492 5364
rect 24544 5352 24550 5364
rect 25225 5355 25283 5361
rect 25225 5352 25237 5355
rect 24544 5324 25237 5352
rect 24544 5312 24550 5324
rect 25225 5321 25237 5324
rect 25271 5321 25283 5355
rect 25225 5315 25283 5321
rect 26050 5312 26056 5364
rect 26108 5352 26114 5364
rect 26697 5355 26755 5361
rect 26697 5352 26709 5355
rect 26108 5324 26709 5352
rect 26108 5312 26114 5324
rect 26697 5321 26709 5324
rect 26743 5321 26755 5355
rect 26697 5315 26755 5321
rect 23750 5284 23756 5296
rect 23124 5256 23756 5284
rect 20119 5120 20392 5148
rect 20441 5151 20499 5157
rect 20119 5117 20131 5120
rect 20073 5111 20131 5117
rect 20441 5117 20453 5151
rect 20487 5148 20499 5151
rect 20990 5148 20996 5160
rect 20487 5120 20996 5148
rect 20487 5117 20499 5120
rect 20441 5111 20499 5117
rect 20990 5108 20996 5120
rect 21048 5148 21054 5160
rect 21818 5148 21824 5160
rect 21048 5120 21824 5148
rect 21048 5108 21054 5120
rect 21818 5108 21824 5120
rect 21876 5108 21882 5160
rect 23124 5157 23152 5256
rect 23750 5244 23756 5256
rect 23808 5244 23814 5296
rect 23382 5176 23388 5228
rect 23440 5176 23446 5228
rect 23474 5176 23480 5228
rect 23532 5216 23538 5228
rect 23845 5219 23903 5225
rect 23845 5216 23857 5219
rect 23532 5188 23857 5216
rect 23532 5176 23538 5188
rect 23845 5185 23857 5188
rect 23891 5185 23903 5219
rect 23845 5179 23903 5185
rect 23109 5151 23167 5157
rect 23109 5117 23121 5151
rect 23155 5117 23167 5151
rect 23109 5111 23167 5117
rect 23293 5151 23351 5157
rect 23293 5117 23305 5151
rect 23339 5117 23351 5151
rect 23293 5111 23351 5117
rect 23661 5151 23719 5157
rect 23661 5117 23673 5151
rect 23707 5148 23719 5151
rect 23750 5148 23756 5160
rect 23707 5120 23756 5148
rect 23707 5117 23719 5120
rect 23661 5111 23719 5117
rect 16666 5080 16672 5092
rect 14001 5043 14059 5049
rect 14384 5052 15240 5080
rect 15396 5052 16672 5080
rect 9456 4984 11841 5012
rect 9456 4972 9462 4984
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 11940 4984 12173 5012
rect 11940 4972 11946 4984
rect 12161 4981 12173 4984
rect 12207 4981 12219 5015
rect 12161 4975 12219 4981
rect 13909 5015 13967 5021
rect 13909 4981 13921 5015
rect 13955 5012 13967 5015
rect 14384 5012 14412 5052
rect 13955 4984 14412 5012
rect 15212 5012 15240 5052
rect 16666 5040 16672 5052
rect 16724 5040 16730 5092
rect 19981 5083 20039 5089
rect 19981 5049 19993 5083
rect 20027 5080 20039 5083
rect 20686 5083 20744 5089
rect 20686 5080 20698 5083
rect 20027 5052 20698 5080
rect 20027 5049 20039 5052
rect 19981 5043 20039 5049
rect 20686 5049 20698 5052
rect 20732 5049 20744 5083
rect 23308 5080 23336 5111
rect 23750 5108 23756 5120
rect 23808 5108 23814 5160
rect 23860 5148 23888 5179
rect 25317 5151 25375 5157
rect 25317 5148 25329 5151
rect 23860 5120 25329 5148
rect 25317 5117 25329 5120
rect 25363 5117 25375 5151
rect 25317 5111 25375 5117
rect 23385 5083 23443 5089
rect 23385 5080 23397 5083
rect 23308 5052 23397 5080
rect 20686 5043 20744 5049
rect 23385 5049 23397 5052
rect 23431 5049 23443 5083
rect 24090 5083 24148 5089
rect 24090 5080 24102 5083
rect 23385 5043 23443 5049
rect 23676 5052 24102 5080
rect 17957 5015 18015 5021
rect 17957 5012 17969 5015
rect 15212 4984 17969 5012
rect 13955 4981 13967 4984
rect 13909 4975 13967 4981
rect 17957 4981 17969 4984
rect 18003 5012 18015 5015
rect 19150 5012 19156 5024
rect 18003 4984 19156 5012
rect 18003 4981 18015 4984
rect 17957 4975 18015 4981
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 23201 5015 23259 5021
rect 23201 4981 23213 5015
rect 23247 5012 23259 5015
rect 23676 5012 23704 5052
rect 24090 5049 24102 5052
rect 24136 5049 24148 5083
rect 24090 5043 24148 5049
rect 25406 5040 25412 5092
rect 25464 5080 25470 5092
rect 25562 5083 25620 5089
rect 25562 5080 25574 5083
rect 25464 5052 25574 5080
rect 25464 5040 25470 5052
rect 25562 5049 25574 5052
rect 25608 5049 25620 5083
rect 25562 5043 25620 5049
rect 23247 4984 23704 5012
rect 23247 4981 23259 4984
rect 23201 4975 23259 4981
rect 552 4922 27576 4944
rect 552 4870 7114 4922
rect 7166 4870 7178 4922
rect 7230 4870 7242 4922
rect 7294 4870 7306 4922
rect 7358 4870 7370 4922
rect 7422 4870 13830 4922
rect 13882 4870 13894 4922
rect 13946 4870 13958 4922
rect 14010 4870 14022 4922
rect 14074 4870 14086 4922
rect 14138 4870 20546 4922
rect 20598 4870 20610 4922
rect 20662 4870 20674 4922
rect 20726 4870 20738 4922
rect 20790 4870 20802 4922
rect 20854 4870 27262 4922
rect 27314 4870 27326 4922
rect 27378 4870 27390 4922
rect 27442 4870 27454 4922
rect 27506 4870 27518 4922
rect 27570 4870 27576 4922
rect 552 4848 27576 4870
rect 4433 4811 4491 4817
rect 4433 4777 4445 4811
rect 4479 4808 4491 4811
rect 4522 4808 4528 4820
rect 4479 4780 4528 4808
rect 4479 4777 4491 4780
rect 4433 4771 4491 4777
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 4706 4768 4712 4820
rect 4764 4768 4770 4820
rect 7926 4768 7932 4820
rect 7984 4768 7990 4820
rect 8478 4768 8484 4820
rect 8536 4768 8542 4820
rect 12345 4811 12403 4817
rect 8588 4780 12296 4808
rect 4154 4740 4160 4752
rect 3068 4712 4160 4740
rect 3068 4681 3096 4712
rect 4154 4700 4160 4712
rect 4212 4700 4218 4752
rect 5626 4740 5632 4752
rect 5000 4712 5632 4740
rect 3326 4681 3332 4684
rect 3053 4675 3111 4681
rect 3053 4641 3065 4675
rect 3099 4641 3111 4675
rect 3320 4672 3332 4681
rect 3287 4644 3332 4672
rect 3053 4635 3111 4641
rect 3320 4635 3332 4644
rect 3326 4632 3332 4635
rect 3384 4632 3390 4684
rect 5000 4681 5028 4712
rect 5626 4700 5632 4712
rect 5684 4700 5690 4752
rect 8386 4740 8392 4752
rect 8036 4712 8392 4740
rect 4985 4675 5043 4681
rect 4985 4641 4997 4675
rect 5031 4641 5043 4675
rect 4985 4635 5043 4641
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4641 5135 4675
rect 5077 4635 5135 4641
rect 4338 4564 4344 4616
rect 4396 4604 4402 4616
rect 5092 4604 5120 4635
rect 5166 4632 5172 4684
rect 5224 4632 5230 4684
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 5353 4675 5411 4681
rect 5353 4672 5365 4675
rect 5316 4644 5365 4672
rect 5316 4632 5322 4644
rect 5353 4641 5365 4644
rect 5399 4672 5411 4675
rect 5399 4644 7696 4672
rect 5399 4641 5411 4644
rect 5353 4635 5411 4641
rect 6730 4604 6736 4616
rect 4396 4576 6736 4604
rect 4396 4564 4402 4576
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 7561 4471 7619 4477
rect 7561 4468 7573 4471
rect 7524 4440 7573 4468
rect 7524 4428 7530 4440
rect 7561 4437 7573 4440
rect 7607 4437 7619 4471
rect 7668 4468 7696 4644
rect 7742 4632 7748 4684
rect 7800 4632 7806 4684
rect 8036 4681 8064 4712
rect 8386 4700 8392 4712
rect 8444 4740 8450 4752
rect 8588 4740 8616 4780
rect 12066 4740 12072 4752
rect 8444 4712 8616 4740
rect 8444 4700 8450 4712
rect 8588 4681 8616 4712
rect 10612 4712 12072 4740
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4641 8079 4675
rect 8021 4635 8079 4641
rect 8297 4675 8355 4681
rect 8297 4641 8309 4675
rect 8343 4641 8355 4675
rect 8297 4635 8355 4641
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4641 8631 4675
rect 8573 4635 8631 4641
rect 7760 4604 7788 4632
rect 8312 4604 8340 4635
rect 10042 4632 10048 4684
rect 10100 4672 10106 4684
rect 10612 4681 10640 4712
rect 12066 4700 12072 4712
rect 12124 4700 12130 4752
rect 12268 4740 12296 4780
rect 12345 4777 12357 4811
rect 12391 4808 12403 4811
rect 12618 4808 12624 4820
rect 12391 4780 12624 4808
rect 12391 4777 12403 4780
rect 12345 4771 12403 4777
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 12805 4811 12863 4817
rect 12805 4777 12817 4811
rect 12851 4808 12863 4811
rect 13170 4808 13176 4820
rect 12851 4780 13176 4808
rect 12851 4777 12863 4780
rect 12805 4771 12863 4777
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 13817 4811 13875 4817
rect 13817 4777 13829 4811
rect 13863 4808 13875 4811
rect 14182 4808 14188 4820
rect 13863 4780 14188 4808
rect 13863 4777 13875 4780
rect 13817 4771 13875 4777
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 14645 4811 14703 4817
rect 14645 4808 14657 4811
rect 14424 4780 14657 4808
rect 14424 4768 14430 4780
rect 14645 4777 14657 4780
rect 14691 4777 14703 4811
rect 19610 4808 19616 4820
rect 14645 4771 14703 4777
rect 14956 4780 19616 4808
rect 13354 4740 13360 4752
rect 12268 4712 13360 4740
rect 13354 4700 13360 4712
rect 13412 4700 13418 4752
rect 14956 4740 14984 4780
rect 14200 4712 14984 4740
rect 15013 4743 15071 4749
rect 10413 4675 10471 4681
rect 10413 4672 10425 4675
rect 10100 4644 10425 4672
rect 10100 4632 10106 4644
rect 10413 4641 10425 4644
rect 10459 4641 10471 4675
rect 10413 4635 10471 4641
rect 10505 4675 10563 4681
rect 10505 4641 10517 4675
rect 10551 4641 10563 4675
rect 10505 4635 10563 4641
rect 10597 4675 10655 4681
rect 10597 4641 10609 4675
rect 10643 4641 10655 4675
rect 10597 4635 10655 4641
rect 8662 4604 8668 4616
rect 7760 4576 8668 4604
rect 8662 4564 8668 4576
rect 8720 4564 8726 4616
rect 9858 4564 9864 4616
rect 9916 4604 9922 4616
rect 10520 4604 10548 4635
rect 10778 4632 10784 4684
rect 10836 4632 10842 4684
rect 10870 4632 10876 4684
rect 10928 4672 10934 4684
rect 10965 4675 11023 4681
rect 10965 4672 10977 4675
rect 10928 4644 10977 4672
rect 10928 4632 10934 4644
rect 10965 4641 10977 4644
rect 11011 4641 11023 4675
rect 10965 4635 11023 4641
rect 11232 4675 11290 4681
rect 11232 4641 11244 4675
rect 11278 4672 11290 4675
rect 12158 4672 12164 4684
rect 11278 4644 12164 4672
rect 11278 4641 11290 4644
rect 11232 4635 11290 4641
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 12526 4632 12532 4684
rect 12584 4672 12590 4684
rect 12621 4675 12679 4681
rect 12621 4672 12633 4675
rect 12584 4644 12633 4672
rect 12584 4632 12590 4644
rect 12621 4641 12633 4644
rect 12667 4641 12679 4675
rect 12621 4635 12679 4641
rect 12894 4632 12900 4684
rect 12952 4632 12958 4684
rect 14200 4681 14228 4712
rect 15013 4709 15025 4743
rect 15059 4740 15071 4743
rect 15059 4712 15332 4740
rect 15059 4709 15071 4712
rect 15013 4703 15071 4709
rect 14185 4675 14243 4681
rect 14185 4641 14197 4675
rect 14231 4641 14243 4675
rect 14185 4635 14243 4641
rect 14366 4632 14372 4684
rect 14424 4672 14430 4684
rect 15105 4675 15163 4681
rect 15105 4672 15117 4675
rect 14424 4644 15117 4672
rect 14424 4632 14430 4644
rect 15105 4641 15117 4644
rect 15151 4641 15163 4675
rect 15304 4672 15332 4712
rect 15378 4700 15384 4752
rect 15436 4740 15442 4752
rect 15436 4712 16344 4740
rect 15436 4700 15442 4712
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 15304 4644 16221 4672
rect 15105 4635 15163 4641
rect 16209 4641 16221 4644
rect 16255 4641 16267 4675
rect 16316 4672 16344 4712
rect 16390 4700 16396 4752
rect 16448 4700 16454 4752
rect 16485 4675 16543 4681
rect 16485 4672 16497 4675
rect 16316 4644 16497 4672
rect 16209 4635 16267 4641
rect 16485 4641 16497 4644
rect 16531 4641 16543 4675
rect 16485 4635 16543 4641
rect 9916 4576 10548 4604
rect 9916 4564 9922 4576
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 14458 4564 14464 4616
rect 14516 4604 14522 4616
rect 15010 4604 15016 4616
rect 14516 4576 15016 4604
rect 14516 4564 14522 4576
rect 15010 4564 15016 4576
rect 15068 4604 15074 4616
rect 15197 4607 15255 4613
rect 15197 4604 15209 4607
rect 15068 4576 15209 4604
rect 15068 4564 15074 4576
rect 15197 4573 15209 4576
rect 15243 4573 15255 4607
rect 16224 4604 16252 4635
rect 16574 4632 16580 4684
rect 16632 4632 16638 4684
rect 16859 4681 16887 4780
rect 19610 4768 19616 4780
rect 19668 4768 19674 4820
rect 23750 4768 23756 4820
rect 23808 4768 23814 4820
rect 24670 4768 24676 4820
rect 24728 4808 24734 4820
rect 24781 4811 24839 4817
rect 24781 4808 24793 4811
rect 24728 4780 24793 4808
rect 24728 4768 24734 4780
rect 24781 4777 24793 4780
rect 24827 4777 24839 4811
rect 24781 4771 24839 4777
rect 24949 4811 25007 4817
rect 24949 4777 24961 4811
rect 24995 4777 25007 4811
rect 24949 4771 25007 4777
rect 25225 4811 25283 4817
rect 25225 4777 25237 4811
rect 25271 4808 25283 4811
rect 25406 4808 25412 4820
rect 25271 4780 25412 4808
rect 25271 4777 25283 4780
rect 25225 4771 25283 4777
rect 17034 4700 17040 4752
rect 17092 4700 17098 4752
rect 17126 4700 17132 4752
rect 17184 4700 17190 4752
rect 24578 4700 24584 4752
rect 24636 4700 24642 4752
rect 16853 4675 16911 4681
rect 16853 4641 16865 4675
rect 16899 4641 16911 4675
rect 16853 4635 16911 4641
rect 17221 4675 17279 4681
rect 17221 4641 17233 4675
rect 17267 4641 17279 4675
rect 17221 4635 17279 4641
rect 18785 4675 18843 4681
rect 18785 4641 18797 4675
rect 18831 4641 18843 4675
rect 18785 4635 18843 4641
rect 16592 4604 16620 4632
rect 17236 4604 17264 4635
rect 16224 4576 16344 4604
rect 16592 4576 17264 4604
rect 15197 4567 15255 4573
rect 8110 4496 8116 4548
rect 8168 4496 8174 4548
rect 10778 4536 10784 4548
rect 8220 4508 10784 4536
rect 8220 4468 8248 4508
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 16316 4536 16344 4576
rect 18598 4564 18604 4616
rect 18656 4564 18662 4616
rect 17405 4539 17463 4545
rect 16316 4508 16887 4536
rect 7668 4440 8248 4468
rect 7561 4431 7619 4437
rect 10134 4428 10140 4480
rect 10192 4428 10198 4480
rect 10962 4428 10968 4480
rect 11020 4468 11026 4480
rect 12437 4471 12495 4477
rect 12437 4468 12449 4471
rect 11020 4440 12449 4468
rect 11020 4428 11026 4440
rect 12437 4437 12449 4440
rect 12483 4437 12495 4471
rect 12437 4431 12495 4437
rect 16758 4428 16764 4480
rect 16816 4428 16822 4480
rect 16859 4468 16887 4508
rect 17405 4505 17417 4539
rect 17451 4536 17463 4539
rect 18800 4536 18828 4635
rect 24394 4632 24400 4684
rect 24452 4632 24458 4684
rect 24964 4672 24992 4771
rect 25406 4768 25412 4780
rect 25464 4768 25470 4820
rect 25041 4675 25099 4681
rect 25041 4672 25053 4675
rect 24964 4644 25053 4672
rect 25041 4641 25053 4644
rect 25087 4641 25099 4675
rect 25041 4635 25099 4641
rect 19518 4536 19524 4548
rect 17451 4508 18828 4536
rect 18892 4508 19524 4536
rect 17451 4505 17463 4508
rect 17405 4499 17463 4505
rect 18892 4468 18920 4508
rect 19518 4496 19524 4508
rect 19576 4496 19582 4548
rect 16859 4440 18920 4468
rect 18969 4471 19027 4477
rect 18969 4437 18981 4471
rect 19015 4468 19027 4471
rect 19334 4468 19340 4480
rect 19015 4440 19340 4468
rect 19015 4437 19027 4440
rect 18969 4431 19027 4437
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 24765 4471 24823 4477
rect 24765 4437 24777 4471
rect 24811 4468 24823 4471
rect 25130 4468 25136 4480
rect 24811 4440 25136 4468
rect 24811 4437 24823 4440
rect 24765 4431 24823 4437
rect 25130 4428 25136 4440
rect 25188 4428 25194 4480
rect 552 4378 27416 4400
rect 552 4326 3756 4378
rect 3808 4326 3820 4378
rect 3872 4326 3884 4378
rect 3936 4326 3948 4378
rect 4000 4326 4012 4378
rect 4064 4326 10472 4378
rect 10524 4326 10536 4378
rect 10588 4326 10600 4378
rect 10652 4326 10664 4378
rect 10716 4326 10728 4378
rect 10780 4326 17188 4378
rect 17240 4326 17252 4378
rect 17304 4326 17316 4378
rect 17368 4326 17380 4378
rect 17432 4326 17444 4378
rect 17496 4326 23904 4378
rect 23956 4326 23968 4378
rect 24020 4326 24032 4378
rect 24084 4326 24096 4378
rect 24148 4326 24160 4378
rect 24212 4326 27416 4378
rect 552 4304 27416 4326
rect 5534 4264 5540 4276
rect 4908 4236 5540 4264
rect 3053 4199 3111 4205
rect 3053 4165 3065 4199
rect 3099 4196 3111 4199
rect 3099 4168 4660 4196
rect 3099 4165 3111 4168
rect 3053 4159 3111 4165
rect 4154 4128 4160 4140
rect 2746 4100 4160 4128
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4060 1731 4063
rect 2746 4060 2774 4100
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4522 4128 4528 4140
rect 4356 4100 4528 4128
rect 1719 4032 2774 4060
rect 3605 4063 3663 4069
rect 1719 4029 1731 4032
rect 1673 4023 1731 4029
rect 3605 4029 3617 4063
rect 3651 4029 3663 4063
rect 3605 4023 3663 4029
rect 1940 3995 1998 4001
rect 1940 3961 1952 3995
rect 1986 3992 1998 3995
rect 2774 3992 2780 4004
rect 1986 3964 2780 3992
rect 1986 3961 1998 3964
rect 1940 3955 1998 3961
rect 2774 3952 2780 3964
rect 2832 3952 2838 4004
rect 3620 3992 3648 4023
rect 3786 4020 3792 4072
rect 3844 4020 3850 4072
rect 4062 4020 4068 4072
rect 4120 4020 4126 4072
rect 4356 4060 4384 4100
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 4632 4072 4660 4168
rect 4908 4128 4936 4236
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 10042 4224 10048 4276
rect 10100 4224 10106 4276
rect 12158 4224 12164 4276
rect 12216 4224 12222 4276
rect 16574 4224 16580 4276
rect 16632 4264 16638 4276
rect 17034 4264 17040 4276
rect 16632 4236 17040 4264
rect 16632 4224 16638 4236
rect 17034 4224 17040 4236
rect 17092 4224 17098 4276
rect 19610 4224 19616 4276
rect 19668 4264 19674 4276
rect 19978 4264 19984 4276
rect 19668 4236 19984 4264
rect 19668 4224 19674 4236
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 6914 4156 6920 4208
rect 6972 4196 6978 4208
rect 8110 4196 8116 4208
rect 6972 4168 8116 4196
rect 6972 4156 6978 4168
rect 8110 4156 8116 4168
rect 8168 4156 8174 4208
rect 8662 4156 8668 4208
rect 8720 4196 8726 4208
rect 12526 4196 12532 4208
rect 8720 4168 12532 4196
rect 8720 4156 8726 4168
rect 12526 4156 12532 4168
rect 12584 4196 12590 4208
rect 12584 4168 13768 4196
rect 12584 4156 12590 4168
rect 5534 4128 5540 4140
rect 4816 4100 4936 4128
rect 5000 4100 5540 4128
rect 4172 4032 4384 4060
rect 4433 4063 4491 4069
rect 4172 4001 4200 4032
rect 4433 4029 4445 4063
rect 4479 4060 4491 4063
rect 4614 4060 4620 4072
rect 4479 4032 4620 4060
rect 4479 4029 4491 4032
rect 4433 4023 4491 4029
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 4706 4020 4712 4072
rect 4764 4020 4770 4072
rect 4816 4069 4844 4100
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4029 4859 4063
rect 4801 4023 4859 4029
rect 4893 4063 4951 4069
rect 4893 4029 4905 4063
rect 4939 4060 4951 4063
rect 5000 4060 5028 4100
rect 5534 4088 5540 4100
rect 5592 4128 5598 4140
rect 5902 4128 5908 4140
rect 5592 4100 5908 4128
rect 5592 4088 5598 4100
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 12253 4131 12311 4137
rect 12253 4128 12265 4131
rect 11440 4100 12265 4128
rect 4939 4032 5028 4060
rect 4939 4029 4951 4032
rect 4893 4023 4951 4029
rect 4157 3995 4215 4001
rect 3620 3964 3924 3992
rect 3418 3884 3424 3936
rect 3476 3884 3482 3936
rect 3896 3933 3924 3964
rect 4157 3961 4169 3995
rect 4203 3961 4215 3995
rect 4157 3955 4215 3961
rect 4249 3995 4307 4001
rect 4249 3961 4261 3995
rect 4295 3992 4307 3995
rect 4908 3992 4936 4023
rect 5074 4020 5080 4072
rect 5132 4020 5138 4072
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4029 6699 4063
rect 6641 4023 6699 4029
rect 4295 3964 4936 3992
rect 4295 3961 4307 3964
rect 4249 3955 4307 3961
rect 4982 3952 4988 4004
rect 5040 3992 5046 4004
rect 5353 3995 5411 4001
rect 5353 3992 5365 3995
rect 5040 3964 5365 3992
rect 5040 3952 5046 3964
rect 5353 3961 5365 3964
rect 5399 3961 5411 3995
rect 6656 3992 6684 4023
rect 6730 4020 6736 4072
rect 6788 4020 6794 4072
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 6914 4060 6920 4072
rect 6871 4032 6920 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 6914 4020 6920 4032
rect 6972 4020 6978 4072
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4060 7067 4063
rect 7558 4060 7564 4072
rect 7055 4032 7564 4060
rect 7055 4029 7067 4032
rect 7009 4023 7067 4029
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 7650 4020 7656 4072
rect 7708 4020 7714 4072
rect 8386 4020 8392 4072
rect 8444 4020 8450 4072
rect 8662 4020 8668 4072
rect 8720 4020 8726 4072
rect 10686 4020 10692 4072
rect 10744 4020 10750 4072
rect 10778 4020 10784 4072
rect 10836 4020 10842 4072
rect 10962 4020 10968 4072
rect 11020 4020 11026 4072
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 11195 4063 11253 4069
rect 11112 4032 11157 4060
rect 11112 4020 11118 4032
rect 11195 4029 11207 4063
rect 11241 4060 11253 4063
rect 11440 4060 11468 4100
rect 12253 4097 12265 4100
rect 12299 4097 12311 4131
rect 12253 4091 12311 4097
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 13541 4131 13599 4137
rect 13541 4128 13553 4131
rect 12400 4100 13553 4128
rect 12400 4088 12406 4100
rect 13541 4097 13553 4100
rect 13587 4097 13599 4131
rect 13541 4091 13599 4097
rect 11241 4032 11468 4060
rect 11241 4029 11253 4032
rect 11195 4023 11253 4029
rect 11514 4020 11520 4072
rect 11572 4020 11578 4072
rect 11698 4020 11704 4072
rect 11756 4020 11762 4072
rect 11790 4020 11796 4072
rect 11848 4020 11854 4072
rect 11882 4020 11888 4072
rect 11940 4020 11946 4072
rect 13740 4069 13768 4168
rect 16758 4156 16764 4208
rect 16816 4196 16822 4208
rect 16816 4168 16896 4196
rect 16816 4156 16822 4168
rect 16390 4088 16396 4140
rect 16448 4128 16454 4140
rect 16868 4128 16896 4168
rect 16942 4156 16948 4208
rect 17000 4196 17006 4208
rect 17310 4196 17316 4208
rect 17000 4168 17316 4196
rect 17000 4156 17006 4168
rect 17310 4156 17316 4168
rect 17368 4196 17374 4208
rect 17678 4196 17684 4208
rect 17368 4168 17684 4196
rect 17368 4156 17374 4168
rect 17678 4156 17684 4168
rect 17736 4196 17742 4208
rect 18598 4196 18604 4208
rect 17736 4168 18604 4196
rect 17736 4156 17742 4168
rect 18598 4156 18604 4168
rect 18656 4196 18662 4208
rect 18656 4168 18736 4196
rect 18656 4156 18662 4168
rect 18708 4137 18736 4168
rect 18693 4131 18751 4137
rect 16448 4100 16796 4128
rect 16868 4100 17448 4128
rect 16448 4088 16454 4100
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12268 4032 12817 4060
rect 12268 4004 12296 4032
rect 12805 4029 12817 4032
rect 12851 4029 12863 4063
rect 12805 4023 12863 4029
rect 13725 4063 13783 4069
rect 13725 4029 13737 4063
rect 13771 4029 13783 4063
rect 13725 4023 13783 4029
rect 14001 4063 14059 4069
rect 14001 4029 14013 4063
rect 14047 4060 14059 4063
rect 14182 4060 14188 4072
rect 14047 4032 14188 4060
rect 14047 4029 14059 4032
rect 14001 4023 14059 4029
rect 14182 4020 14188 4032
rect 14240 4060 14246 4072
rect 14240 4032 14504 4060
rect 14240 4020 14246 4032
rect 7101 3995 7159 4001
rect 7101 3992 7113 3995
rect 6656 3964 7113 3992
rect 5353 3955 5411 3961
rect 7101 3961 7113 3964
rect 7147 3961 7159 3995
rect 7101 3955 7159 3961
rect 8481 3995 8539 4001
rect 8481 3961 8493 3995
rect 8527 3992 8539 3995
rect 12066 3992 12072 4004
rect 8527 3964 12072 3992
rect 8527 3961 8539 3964
rect 8481 3955 8539 3961
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 12250 3952 12256 4004
rect 12308 3952 12314 4004
rect 12342 3952 12348 4004
rect 12400 3992 12406 4004
rect 14366 3992 14372 4004
rect 12400 3964 14372 3992
rect 12400 3952 12406 3964
rect 14366 3952 14372 3964
rect 14424 3952 14430 4004
rect 14476 3992 14504 4032
rect 15102 4020 15108 4072
rect 15160 4060 15166 4072
rect 16669 4063 16727 4069
rect 15160 4054 16620 4060
rect 16669 4054 16681 4063
rect 15160 4032 16681 4054
rect 15160 4020 15166 4032
rect 16592 4029 16681 4032
rect 16715 4029 16727 4063
rect 16768 4060 16796 4100
rect 16853 4063 16911 4069
rect 16853 4060 16865 4063
rect 16768 4032 16865 4060
rect 16592 4026 16727 4029
rect 16669 4023 16727 4026
rect 16853 4029 16865 4032
rect 16899 4029 16911 4063
rect 16853 4023 16911 4029
rect 15286 3992 15292 4004
rect 14476 3964 15292 3992
rect 15286 3952 15292 3964
rect 15344 3992 15350 4004
rect 15654 3992 15660 4004
rect 15344 3964 15660 3992
rect 15344 3952 15350 3964
rect 15654 3952 15660 3964
rect 15712 3952 15718 4004
rect 16684 3992 16712 4023
rect 17034 4020 17040 4072
rect 17092 4020 17098 4072
rect 17310 4020 17316 4072
rect 17368 4020 17374 4072
rect 17420 4060 17448 4100
rect 18693 4097 18705 4131
rect 18739 4128 18751 4131
rect 18739 4100 19472 4128
rect 18739 4097 18751 4100
rect 18693 4091 18751 4097
rect 17497 4063 17555 4069
rect 17497 4060 17509 4063
rect 17420 4032 17509 4060
rect 17497 4029 17509 4032
rect 17543 4029 17555 4063
rect 17497 4023 17555 4029
rect 17681 4063 17739 4069
rect 17681 4029 17693 4063
rect 17727 4060 17739 4063
rect 17865 4063 17923 4069
rect 17865 4060 17877 4063
rect 17727 4032 17877 4060
rect 17727 4029 17739 4032
rect 17681 4023 17739 4029
rect 17865 4029 17877 4032
rect 17911 4029 17923 4063
rect 17865 4023 17923 4029
rect 18877 4063 18935 4069
rect 18877 4029 18889 4063
rect 18923 4029 18935 4063
rect 18877 4023 18935 4029
rect 16758 3992 16764 4004
rect 16684 3964 16764 3992
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 16945 3995 17003 4001
rect 16945 3961 16957 3995
rect 16991 3961 17003 3995
rect 18892 3992 18920 4023
rect 19334 4020 19340 4072
rect 19392 4020 19398 4072
rect 19444 4060 19472 4100
rect 20990 4088 20996 4140
rect 21048 4088 21054 4140
rect 23937 4063 23995 4069
rect 23937 4060 23949 4063
rect 19444 4032 23949 4060
rect 23937 4029 23949 4032
rect 23983 4060 23995 4063
rect 24578 4060 24584 4072
rect 23983 4032 24584 4060
rect 23983 4029 23995 4032
rect 23937 4023 23995 4029
rect 24578 4020 24584 4032
rect 24636 4020 24642 4072
rect 20726 3995 20784 4001
rect 20726 3992 20738 3995
rect 16945 3955 17003 3961
rect 17236 3964 18920 3992
rect 19536 3964 20738 3992
rect 3881 3927 3939 3933
rect 3881 3893 3893 3927
rect 3927 3893 3939 3927
rect 3881 3887 3939 3893
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4525 3927 4583 3933
rect 4525 3924 4537 3927
rect 4028 3896 4537 3924
rect 4028 3884 4034 3896
rect 4525 3893 4537 3896
rect 4571 3893 4583 3927
rect 4525 3887 4583 3893
rect 5258 3884 5264 3936
rect 5316 3884 5322 3936
rect 6362 3884 6368 3936
rect 6420 3884 6426 3936
rect 8849 3927 8907 3933
rect 8849 3893 8861 3927
rect 8895 3924 8907 3927
rect 9582 3924 9588 3936
rect 8895 3896 9588 3924
rect 8895 3893 8907 3896
rect 8849 3887 8907 3893
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 10778 3884 10784 3936
rect 10836 3924 10842 3936
rect 11330 3924 11336 3936
rect 10836 3896 11336 3924
rect 10836 3884 10842 3896
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11422 3884 11428 3936
rect 11480 3884 11486 3936
rect 12802 3884 12808 3936
rect 12860 3924 12866 3936
rect 13909 3927 13967 3933
rect 13909 3924 13921 3927
rect 12860 3896 13921 3924
rect 12860 3884 12866 3896
rect 13909 3893 13921 3896
rect 13955 3924 13967 3927
rect 16960 3924 16988 3955
rect 17236 3933 17264 3964
rect 13955 3896 16988 3924
rect 17221 3927 17279 3933
rect 13955 3893 13967 3896
rect 13909 3887 13967 3893
rect 17221 3893 17233 3927
rect 17267 3893 17279 3927
rect 17221 3887 17279 3893
rect 18046 3884 18052 3936
rect 18104 3884 18110 3936
rect 19061 3927 19119 3933
rect 19061 3893 19073 3927
rect 19107 3924 19119 3927
rect 19426 3924 19432 3936
rect 19107 3896 19432 3924
rect 19107 3893 19119 3896
rect 19061 3887 19119 3893
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 19536 3933 19564 3964
rect 20726 3961 20738 3964
rect 20772 3961 20784 3995
rect 20726 3955 20784 3961
rect 23014 3952 23020 4004
rect 23072 3992 23078 4004
rect 24121 3995 24179 4001
rect 24121 3992 24133 3995
rect 23072 3964 24133 3992
rect 23072 3952 23078 3964
rect 24121 3961 24133 3964
rect 24167 3961 24179 3995
rect 24121 3955 24179 3961
rect 19521 3927 19579 3933
rect 19521 3893 19533 3927
rect 19567 3893 19579 3927
rect 19521 3887 19579 3893
rect 552 3834 27576 3856
rect 552 3782 7114 3834
rect 7166 3782 7178 3834
rect 7230 3782 7242 3834
rect 7294 3782 7306 3834
rect 7358 3782 7370 3834
rect 7422 3782 13830 3834
rect 13882 3782 13894 3834
rect 13946 3782 13958 3834
rect 14010 3782 14022 3834
rect 14074 3782 14086 3834
rect 14138 3782 20546 3834
rect 20598 3782 20610 3834
rect 20662 3782 20674 3834
rect 20726 3782 20738 3834
rect 20790 3782 20802 3834
rect 20854 3782 27262 3834
rect 27314 3782 27326 3834
rect 27378 3782 27390 3834
rect 27442 3782 27454 3834
rect 27506 3782 27518 3834
rect 27570 3782 27576 3834
rect 552 3760 27576 3782
rect 2774 3680 2780 3732
rect 2832 3680 2838 3732
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 4706 3720 4712 3732
rect 4120 3692 4712 3720
rect 4120 3680 4126 3692
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 7834 3720 7840 3732
rect 4856 3692 7840 3720
rect 4856 3680 4862 3692
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 10781 3723 10839 3729
rect 10781 3720 10793 3723
rect 10744 3692 10793 3720
rect 10744 3680 10750 3692
rect 10781 3689 10793 3692
rect 10827 3720 10839 3723
rect 10962 3720 10968 3732
rect 10827 3692 10968 3720
rect 10827 3689 10839 3692
rect 10781 3683 10839 3689
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 12345 3723 12403 3729
rect 12345 3720 12357 3723
rect 12308 3692 12357 3720
rect 12308 3680 12314 3692
rect 12345 3689 12357 3692
rect 12391 3689 12403 3723
rect 12345 3683 12403 3689
rect 12710 3680 12716 3732
rect 12768 3720 12774 3732
rect 13173 3723 13231 3729
rect 13173 3720 13185 3723
rect 12768 3692 13185 3720
rect 12768 3680 12774 3692
rect 13173 3689 13185 3692
rect 13219 3689 13231 3723
rect 13173 3683 13231 3689
rect 13541 3723 13599 3729
rect 13541 3689 13553 3723
rect 13587 3720 13599 3723
rect 15102 3720 15108 3732
rect 13587 3692 15108 3720
rect 13587 3689 13599 3692
rect 13541 3683 13599 3689
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 15194 3680 15200 3732
rect 15252 3680 15258 3732
rect 16022 3680 16028 3732
rect 16080 3720 16086 3732
rect 16117 3723 16175 3729
rect 16117 3720 16129 3723
rect 16080 3692 16129 3720
rect 16080 3680 16086 3692
rect 16117 3689 16129 3692
rect 16163 3689 16175 3723
rect 16117 3683 16175 3689
rect 16482 3680 16488 3732
rect 16540 3680 16546 3732
rect 16758 3680 16764 3732
rect 16816 3720 16822 3732
rect 16816 3692 19334 3720
rect 16816 3680 16822 3692
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 5442 3652 5448 3664
rect 4212 3624 5448 3652
rect 4212 3612 4218 3624
rect 5442 3612 5448 3624
rect 5500 3652 5506 3664
rect 6172 3655 6230 3661
rect 5500 3624 5948 3652
rect 5500 3612 5506 3624
rect 2961 3587 3019 3593
rect 2961 3553 2973 3587
rect 3007 3584 3019 3587
rect 3418 3584 3424 3596
rect 3007 3556 3424 3584
rect 3007 3553 3019 3556
rect 2961 3547 3019 3553
rect 3418 3544 3424 3556
rect 3476 3544 3482 3596
rect 3970 3544 3976 3596
rect 4028 3544 4034 3596
rect 4172 3584 4200 3612
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 4172 3556 4261 3584
rect 4249 3553 4261 3556
rect 4295 3553 4307 3587
rect 4249 3547 4307 3553
rect 4516 3587 4574 3593
rect 4516 3553 4528 3587
rect 4562 3584 4574 3587
rect 5810 3584 5816 3596
rect 4562 3556 5816 3584
rect 4562 3553 4574 3556
rect 4516 3547 4574 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 5920 3593 5948 3624
rect 6172 3621 6184 3655
rect 6218 3652 6230 3655
rect 6362 3652 6368 3664
rect 6218 3624 6368 3652
rect 6218 3621 6230 3624
rect 6172 3615 6230 3621
rect 6362 3612 6368 3624
rect 6420 3612 6426 3664
rect 11232 3655 11290 3661
rect 9416 3624 11008 3652
rect 9416 3596 9444 3624
rect 5905 3587 5963 3593
rect 5905 3553 5917 3587
rect 5951 3553 5963 3587
rect 5905 3547 5963 3553
rect 8869 3587 8927 3593
rect 8869 3553 8881 3587
rect 8915 3584 8927 3587
rect 9030 3584 9036 3596
rect 8915 3556 9036 3584
rect 8915 3553 8927 3556
rect 8869 3547 8927 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 9398 3584 9404 3596
rect 9180 3556 9404 3584
rect 9180 3544 9186 3556
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 9668 3587 9726 3593
rect 9668 3553 9680 3587
rect 9714 3584 9726 3587
rect 10134 3584 10140 3596
rect 9714 3556 10140 3584
rect 9714 3553 9726 3556
rect 9668 3547 9726 3553
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10980 3593 11008 3624
rect 11232 3621 11244 3655
rect 11278 3652 11290 3655
rect 11422 3652 11428 3664
rect 11278 3624 11428 3652
rect 11278 3621 11290 3624
rect 11232 3615 11290 3621
rect 11422 3612 11428 3624
rect 11480 3612 11486 3664
rect 12066 3612 12072 3664
rect 12124 3652 12130 3664
rect 13262 3652 13268 3664
rect 12124 3624 13268 3652
rect 12124 3612 12130 3624
rect 13262 3612 13268 3624
rect 13320 3652 13326 3664
rect 13630 3652 13636 3664
rect 13320 3624 13636 3652
rect 13320 3612 13326 3624
rect 13630 3612 13636 3624
rect 13688 3652 13694 3664
rect 14369 3655 14427 3661
rect 14369 3652 14381 3655
rect 13688 3624 14381 3652
rect 13688 3612 13694 3624
rect 14369 3621 14381 3624
rect 14415 3621 14427 3655
rect 14369 3615 14427 3621
rect 15565 3655 15623 3661
rect 15565 3621 15577 3655
rect 15611 3652 15623 3655
rect 15838 3652 15844 3664
rect 15611 3624 15844 3652
rect 15611 3621 15623 3624
rect 15565 3615 15623 3621
rect 15838 3612 15844 3624
rect 15896 3612 15902 3664
rect 17034 3612 17040 3664
rect 17092 3652 17098 3664
rect 17770 3652 17776 3664
rect 17092 3624 17356 3652
rect 17092 3612 17098 3624
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3553 11023 3587
rect 10965 3547 11023 3553
rect 11514 3544 11520 3596
rect 11572 3584 11578 3596
rect 11572 3556 12020 3584
rect 11572 3544 11578 3556
rect 3786 3476 3792 3528
rect 3844 3516 3850 3528
rect 4157 3519 4215 3525
rect 4157 3516 4169 3519
rect 3844 3488 4169 3516
rect 3844 3476 3850 3488
rect 4157 3485 4169 3488
rect 4203 3485 4215 3519
rect 11992 3516 12020 3556
rect 12250 3544 12256 3596
rect 12308 3584 12314 3596
rect 12621 3587 12679 3593
rect 12621 3584 12633 3587
rect 12308 3556 12633 3584
rect 12308 3544 12314 3556
rect 12621 3553 12633 3556
rect 12667 3553 12679 3587
rect 12621 3547 12679 3553
rect 12710 3544 12716 3596
rect 12768 3544 12774 3596
rect 12802 3544 12808 3596
rect 12860 3544 12866 3596
rect 12986 3544 12992 3596
rect 13044 3544 13050 3596
rect 15856 3556 16804 3584
rect 13633 3519 13691 3525
rect 13633 3516 13645 3519
rect 11992 3488 13645 3516
rect 4157 3479 4215 3485
rect 13633 3485 13645 3488
rect 13679 3485 13691 3519
rect 13633 3479 13691 3485
rect 13817 3519 13875 3525
rect 13817 3485 13829 3519
rect 13863 3516 13875 3519
rect 13998 3516 14004 3528
rect 13863 3488 14004 3516
rect 13863 3485 13875 3488
rect 13817 3479 13875 3485
rect 3602 3340 3608 3392
rect 3660 3380 3666 3392
rect 3789 3383 3847 3389
rect 3789 3380 3801 3383
rect 3660 3352 3801 3380
rect 3660 3340 3666 3352
rect 3789 3349 3801 3352
rect 3835 3349 3847 3383
rect 4172 3380 4200 3479
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 14182 3476 14188 3528
rect 14240 3476 14246 3528
rect 14274 3476 14280 3528
rect 14332 3476 14338 3528
rect 15654 3476 15660 3528
rect 15712 3476 15718 3528
rect 15856 3525 15884 3556
rect 16776 3525 16804 3556
rect 16942 3544 16948 3596
rect 17000 3544 17006 3596
rect 17328 3593 17356 3624
rect 17420 3624 17776 3652
rect 17129 3587 17187 3593
rect 17129 3584 17141 3587
rect 17052 3556 17141 3584
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3485 15899 3519
rect 16577 3519 16635 3525
rect 16577 3516 16589 3519
rect 15841 3479 15899 3485
rect 15948 3488 16589 3516
rect 7834 3408 7840 3460
rect 7892 3448 7898 3460
rect 14737 3451 14795 3457
rect 7892 3420 8064 3448
rect 7892 3408 7898 3420
rect 5350 3380 5356 3392
rect 4172 3352 5356 3380
rect 3789 3343 3847 3349
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 5626 3340 5632 3392
rect 5684 3340 5690 3392
rect 7285 3383 7343 3389
rect 7285 3349 7297 3383
rect 7331 3380 7343 3383
rect 7650 3380 7656 3392
rect 7331 3352 7656 3380
rect 7331 3349 7343 3352
rect 7285 3343 7343 3349
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 7745 3383 7803 3389
rect 7745 3349 7757 3383
rect 7791 3380 7803 3383
rect 7926 3380 7932 3392
rect 7791 3352 7932 3380
rect 7791 3349 7803 3352
rect 7745 3343 7803 3349
rect 7926 3340 7932 3352
rect 7984 3340 7990 3392
rect 8036 3380 8064 3420
rect 14737 3417 14749 3451
rect 14783 3448 14795 3451
rect 15470 3448 15476 3460
rect 14783 3420 15476 3448
rect 14783 3417 14795 3420
rect 14737 3411 14795 3417
rect 15470 3408 15476 3420
rect 15528 3408 15534 3460
rect 15948 3448 15976 3488
rect 16577 3485 16589 3488
rect 16623 3485 16635 3519
rect 16577 3479 16635 3485
rect 16761 3519 16819 3525
rect 16761 3485 16773 3519
rect 16807 3516 16819 3519
rect 16850 3516 16856 3528
rect 16807 3488 16856 3516
rect 16807 3485 16819 3488
rect 16761 3479 16819 3485
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 15580 3420 15976 3448
rect 12342 3380 12348 3392
rect 8036 3352 12348 3380
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 12437 3383 12495 3389
rect 12437 3349 12449 3383
rect 12483 3380 12495 3383
rect 12526 3380 12532 3392
rect 12483 3352 12532 3380
rect 12483 3349 12495 3352
rect 12437 3343 12495 3349
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 13170 3340 13176 3392
rect 13228 3380 13234 3392
rect 15580 3380 15608 3420
rect 16022 3408 16028 3460
rect 16080 3448 16086 3460
rect 16390 3448 16396 3460
rect 16080 3420 16396 3448
rect 16080 3408 16086 3420
rect 16390 3408 16396 3420
rect 16448 3448 16454 3460
rect 16666 3448 16672 3460
rect 16448 3420 16672 3448
rect 16448 3408 16454 3420
rect 16666 3408 16672 3420
rect 16724 3448 16730 3460
rect 17052 3448 17080 3556
rect 17129 3553 17141 3556
rect 17175 3553 17187 3587
rect 17129 3547 17187 3553
rect 17221 3587 17279 3593
rect 17221 3553 17233 3587
rect 17267 3553 17279 3587
rect 17221 3547 17279 3553
rect 17313 3587 17371 3593
rect 17313 3553 17325 3587
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 17236 3516 17264 3547
rect 17420 3516 17448 3624
rect 17770 3612 17776 3624
rect 17828 3612 17834 3664
rect 18046 3612 18052 3664
rect 18104 3652 18110 3664
rect 18386 3655 18444 3661
rect 18386 3652 18398 3655
rect 18104 3624 18398 3652
rect 18104 3612 18110 3624
rect 18386 3621 18398 3624
rect 18432 3621 18444 3655
rect 19306 3652 19334 3692
rect 19518 3680 19524 3732
rect 19576 3680 19582 3732
rect 19613 3723 19671 3729
rect 19613 3689 19625 3723
rect 19659 3689 19671 3723
rect 19613 3683 19671 3689
rect 19628 3652 19656 3683
rect 19886 3652 19892 3664
rect 19306 3624 19892 3652
rect 18386 3615 18444 3621
rect 19886 3612 19892 3624
rect 19944 3612 19950 3664
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 17236 3488 17448 3516
rect 17512 3556 17877 3584
rect 17512 3457 17540 3556
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 17954 3544 17960 3596
rect 18012 3584 18018 3596
rect 19794 3584 19800 3596
rect 18012 3556 19800 3584
rect 18012 3544 18018 3556
rect 19794 3544 19800 3556
rect 19852 3544 19858 3596
rect 20438 3544 20444 3596
rect 20496 3584 20502 3596
rect 20726 3587 20784 3593
rect 20726 3584 20738 3587
rect 20496 3556 20738 3584
rect 20496 3544 20502 3556
rect 20726 3553 20738 3556
rect 20772 3553 20784 3587
rect 20726 3547 20784 3553
rect 20990 3544 20996 3596
rect 21048 3544 21054 3596
rect 17678 3476 17684 3528
rect 17736 3476 17742 3528
rect 18138 3476 18144 3528
rect 18196 3476 18202 3528
rect 16724 3420 17080 3448
rect 17497 3451 17555 3457
rect 16724 3408 16730 3420
rect 17497 3417 17509 3451
rect 17543 3417 17555 3451
rect 17497 3411 17555 3417
rect 13228 3352 15608 3380
rect 18049 3383 18107 3389
rect 13228 3340 13234 3352
rect 18049 3349 18061 3383
rect 18095 3380 18107 3383
rect 18322 3380 18328 3392
rect 18095 3352 18328 3380
rect 18095 3349 18107 3352
rect 18049 3343 18107 3349
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 552 3290 27416 3312
rect 552 3238 3756 3290
rect 3808 3238 3820 3290
rect 3872 3238 3884 3290
rect 3936 3238 3948 3290
rect 4000 3238 4012 3290
rect 4064 3238 10472 3290
rect 10524 3238 10536 3290
rect 10588 3238 10600 3290
rect 10652 3238 10664 3290
rect 10716 3238 10728 3290
rect 10780 3238 17188 3290
rect 17240 3238 17252 3290
rect 17304 3238 17316 3290
rect 17368 3238 17380 3290
rect 17432 3238 17444 3290
rect 17496 3238 23904 3290
rect 23956 3238 23968 3290
rect 24020 3238 24032 3290
rect 24084 3238 24096 3290
rect 24148 3238 24160 3290
rect 24212 3238 27416 3290
rect 552 3216 27416 3238
rect 4154 3176 4160 3188
rect 3252 3148 4160 3176
rect 3252 3049 3280 3148
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 5074 3176 5080 3188
rect 4663 3148 5080 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 6641 3179 6699 3185
rect 6641 3176 6653 3179
rect 5868 3148 6653 3176
rect 5868 3136 5874 3148
rect 6641 3145 6653 3148
rect 6687 3145 6699 3179
rect 6641 3139 6699 3145
rect 6730 3136 6736 3188
rect 6788 3176 6794 3188
rect 8938 3176 8944 3188
rect 6788 3148 8944 3176
rect 6788 3136 6794 3148
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9030 3136 9036 3188
rect 9088 3176 9094 3188
rect 9125 3179 9183 3185
rect 9125 3176 9137 3179
rect 9088 3148 9137 3176
rect 9088 3136 9094 3148
rect 9125 3145 9137 3148
rect 9171 3145 9183 3179
rect 12250 3176 12256 3188
rect 9125 3139 9183 3145
rect 10888 3148 12256 3176
rect 4706 3068 4712 3120
rect 4764 3108 4770 3120
rect 5718 3108 5724 3120
rect 4764 3080 5724 3108
rect 4764 3068 4770 3080
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 5460 3040 5488 3080
rect 5718 3068 5724 3080
rect 5776 3108 5782 3120
rect 7653 3111 7711 3117
rect 5776 3080 7144 3108
rect 5776 3068 5782 3080
rect 5905 3043 5963 3049
rect 5905 3040 5917 3043
rect 3237 3003 3295 3009
rect 5368 3012 5488 3040
rect 5644 3012 5917 3040
rect 5368 2981 5396 3012
rect 5644 2984 5672 3012
rect 5905 3009 5917 3012
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 7116 3040 7144 3080
rect 7653 3077 7665 3111
rect 7699 3108 7711 3111
rect 8846 3108 8852 3120
rect 7699 3080 8852 3108
rect 7699 3077 7711 3080
rect 7653 3071 7711 3077
rect 8846 3068 8852 3080
rect 8904 3068 8910 3120
rect 9306 3068 9312 3120
rect 9364 3108 9370 3120
rect 9364 3080 9996 3108
rect 9364 3068 9370 3080
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 6788 3012 7052 3040
rect 7116 3012 7880 3040
rect 6788 3000 6794 3012
rect 5353 2975 5411 2981
rect 5353 2941 5365 2975
rect 5399 2941 5411 2975
rect 5353 2935 5411 2941
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2972 5503 2975
rect 5626 2972 5632 2984
rect 5491 2944 5632 2972
rect 5491 2941 5503 2944
rect 5445 2935 5503 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 5718 2932 5724 2984
rect 5776 2932 5782 2984
rect 7024 2981 7052 3012
rect 6549 2975 6607 2981
rect 6549 2941 6561 2975
rect 6595 2972 6607 2975
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 6595 2944 6929 2972
rect 6595 2941 6607 2944
rect 6549 2935 6607 2941
rect 6917 2941 6929 2944
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2941 7067 2975
rect 7009 2935 7067 2941
rect 7101 2975 7159 2981
rect 7101 2941 7113 2975
rect 7147 2972 7159 2975
rect 7190 2972 7196 2984
rect 7147 2944 7196 2972
rect 7147 2941 7159 2944
rect 7101 2935 7159 2941
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 7285 2975 7343 2981
rect 7285 2941 7297 2975
rect 7331 2972 7343 2975
rect 7558 2972 7564 2984
rect 7331 2944 7564 2972
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 7558 2932 7564 2944
rect 7616 2932 7622 2984
rect 7852 2981 7880 3012
rect 7944 3012 8401 3040
rect 7944 2984 7972 3012
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 8938 3000 8944 3052
rect 8996 3040 9002 3052
rect 9858 3040 9864 3052
rect 8996 3012 9864 3040
rect 8996 3000 9002 3012
rect 7837 2975 7895 2981
rect 7837 2941 7849 2975
rect 7883 2941 7895 2975
rect 7837 2935 7895 2941
rect 7926 2932 7932 2984
rect 7984 2932 7990 2984
rect 8205 2975 8263 2981
rect 8205 2941 8217 2975
rect 8251 2972 8263 2975
rect 8294 2972 8300 2984
rect 8251 2944 8300 2972
rect 8251 2941 8263 2944
rect 8205 2935 8263 2941
rect 8294 2932 8300 2944
rect 8352 2932 8358 2984
rect 9508 2981 9536 3012
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 9033 2975 9091 2981
rect 9033 2941 9045 2975
rect 9079 2972 9091 2975
rect 9401 2975 9459 2981
rect 9401 2972 9413 2975
rect 9079 2944 9413 2972
rect 9079 2941 9091 2944
rect 9033 2935 9091 2941
rect 9401 2941 9413 2944
rect 9447 2941 9459 2975
rect 9401 2935 9459 2941
rect 9493 2975 9551 2981
rect 9493 2941 9505 2975
rect 9539 2941 9551 2975
rect 9493 2935 9551 2941
rect 9582 2932 9588 2984
rect 9640 2932 9646 2984
rect 9674 2932 9680 2984
rect 9732 2972 9738 2984
rect 9769 2975 9827 2981
rect 9769 2972 9781 2975
rect 9732 2944 9781 2972
rect 9732 2932 9738 2944
rect 9769 2941 9781 2944
rect 9815 2941 9827 2975
rect 9968 2972 9996 3080
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3040 10287 3043
rect 10318 3040 10324 3052
rect 10275 3012 10324 3040
rect 10275 3009 10287 3012
rect 10229 3003 10287 3009
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10888 2981 10916 3148
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 12434 3136 12440 3188
rect 12492 3136 12498 3188
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 13541 3179 13599 3185
rect 13541 3176 13553 3179
rect 13136 3148 13553 3176
rect 13136 3136 13142 3148
rect 13541 3145 13553 3148
rect 13587 3145 13599 3179
rect 13541 3139 13599 3145
rect 16206 3136 16212 3188
rect 16264 3176 16270 3188
rect 16758 3176 16764 3188
rect 16264 3148 16764 3176
rect 16264 3136 16270 3148
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 20165 3179 20223 3185
rect 20165 3176 20177 3179
rect 17000 3148 20177 3176
rect 17000 3136 17006 3148
rect 20165 3145 20177 3148
rect 20211 3176 20223 3179
rect 20346 3176 20352 3188
rect 20211 3148 20352 3176
rect 20211 3145 20223 3148
rect 20165 3139 20223 3145
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 20438 3136 20444 3188
rect 20496 3136 20502 3188
rect 11422 3068 11428 3120
rect 11480 3108 11486 3120
rect 13170 3108 13176 3120
rect 11480 3080 13176 3108
rect 11480 3068 11486 3080
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 13722 3068 13728 3120
rect 13780 3108 13786 3120
rect 13780 3080 15976 3108
rect 13780 3068 13786 3080
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 14185 3043 14243 3049
rect 14185 3040 14197 3043
rect 14056 3012 14197 3040
rect 14056 3000 14062 3012
rect 14185 3009 14197 3012
rect 14231 3040 14243 3043
rect 14458 3040 14464 3052
rect 14231 3012 14464 3040
rect 14231 3009 14243 3012
rect 14185 3003 14243 3009
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 10045 2975 10103 2981
rect 10045 2972 10057 2975
rect 9968 2944 10057 2972
rect 9769 2935 9827 2941
rect 10045 2941 10057 2944
rect 10091 2941 10103 2975
rect 10045 2935 10103 2941
rect 10873 2975 10931 2981
rect 10873 2941 10885 2975
rect 10919 2941 10931 2975
rect 10873 2935 10931 2941
rect 10962 2932 10968 2984
rect 11020 2932 11026 2984
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11514 2972 11520 2984
rect 11287 2944 11520 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 11606 2932 11612 2984
rect 11664 2972 11670 2984
rect 11885 2975 11943 2981
rect 11885 2972 11897 2975
rect 11664 2944 11897 2972
rect 11664 2932 11670 2944
rect 11885 2941 11897 2944
rect 11931 2941 11943 2975
rect 11885 2935 11943 2941
rect 12158 2932 12164 2984
rect 12216 2932 12222 2984
rect 12250 2932 12256 2984
rect 12308 2981 12314 2984
rect 12308 2975 12335 2981
rect 12323 2972 12335 2975
rect 13722 2972 13728 2984
rect 12323 2944 13728 2972
rect 12323 2941 12335 2944
rect 12308 2935 12335 2941
rect 12308 2932 12314 2935
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 13906 2932 13912 2984
rect 13964 2932 13970 2984
rect 3504 2907 3562 2913
rect 3504 2873 3516 2907
rect 3550 2904 3562 2907
rect 3694 2904 3700 2916
rect 3550 2876 3700 2904
rect 3550 2873 3562 2876
rect 3504 2867 3562 2873
rect 3694 2864 3700 2876
rect 3752 2864 3758 2916
rect 5534 2864 5540 2916
rect 5592 2904 5598 2916
rect 6638 2904 6644 2916
rect 5592 2876 6644 2904
rect 5592 2864 5598 2876
rect 6638 2864 6644 2876
rect 6696 2904 6702 2916
rect 8021 2907 8079 2913
rect 8021 2904 8033 2907
rect 6696 2876 8033 2904
rect 6696 2864 6702 2876
rect 8021 2873 8033 2876
rect 8067 2904 8079 2907
rect 11057 2907 11115 2913
rect 11057 2904 11069 2907
rect 8067 2876 11069 2904
rect 8067 2873 8079 2876
rect 8021 2867 8079 2873
rect 11057 2873 11069 2876
rect 11103 2904 11115 2907
rect 12069 2907 12127 2913
rect 12069 2904 12081 2907
rect 11103 2876 12081 2904
rect 11103 2873 11115 2876
rect 11057 2867 11115 2873
rect 12069 2873 12081 2876
rect 12115 2904 12127 2907
rect 12802 2904 12808 2916
rect 12115 2876 12808 2904
rect 12115 2873 12127 2876
rect 12069 2867 12127 2873
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 14001 2907 14059 2913
rect 14001 2904 14013 2907
rect 13556 2876 14013 2904
rect 5166 2796 5172 2848
rect 5224 2796 5230 2848
rect 8110 2796 8116 2848
rect 8168 2836 8174 2848
rect 9674 2836 9680 2848
rect 8168 2808 9680 2836
rect 8168 2796 8174 2808
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 9858 2796 9864 2848
rect 9916 2796 9922 2848
rect 10502 2796 10508 2848
rect 10560 2836 10566 2848
rect 10689 2839 10747 2845
rect 10689 2836 10701 2839
rect 10560 2808 10701 2836
rect 10560 2796 10566 2808
rect 10689 2805 10701 2808
rect 10735 2805 10747 2839
rect 10689 2799 10747 2805
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 13556 2836 13584 2876
rect 14001 2873 14013 2876
rect 14047 2904 14059 2907
rect 14182 2904 14188 2916
rect 14047 2876 14188 2904
rect 14047 2873 14059 2876
rect 14001 2867 14059 2873
rect 14182 2864 14188 2876
rect 14240 2864 14246 2916
rect 14476 2904 14504 3000
rect 15838 2932 15844 2984
rect 15896 2932 15902 2984
rect 15948 2972 15976 3080
rect 16592 3080 16887 3108
rect 16592 3052 16620 3080
rect 16574 3040 16580 3052
rect 16224 3012 16580 3040
rect 16224 2981 16252 3012
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 16209 2975 16267 2981
rect 16209 2972 16221 2975
rect 15948 2944 16221 2972
rect 16209 2941 16221 2944
rect 16255 2941 16267 2975
rect 16209 2935 16267 2941
rect 16482 2932 16488 2984
rect 16540 2932 16546 2984
rect 16758 2932 16764 2984
rect 16816 2932 16822 2984
rect 16859 2981 16887 3080
rect 18138 3000 18144 3052
rect 18196 3040 18202 3052
rect 18785 3043 18843 3049
rect 18785 3040 18797 3043
rect 18196 3012 18797 3040
rect 18196 3000 18202 3012
rect 18785 3009 18797 3012
rect 18831 3009 18843 3043
rect 18785 3003 18843 3009
rect 16853 2975 16911 2981
rect 16853 2941 16865 2975
rect 16899 2941 16911 2975
rect 16853 2935 16911 2941
rect 18322 2932 18328 2984
rect 18380 2932 18386 2984
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 20257 2975 20315 2981
rect 20257 2972 20269 2975
rect 19484 2944 20269 2972
rect 19484 2932 19490 2944
rect 20257 2941 20269 2944
rect 20303 2941 20315 2975
rect 20257 2935 20315 2941
rect 14737 2907 14795 2913
rect 14737 2904 14749 2907
rect 14476 2876 14749 2904
rect 14737 2873 14749 2876
rect 14783 2873 14795 2907
rect 14737 2867 14795 2873
rect 16022 2864 16028 2916
rect 16080 2864 16086 2916
rect 16114 2864 16120 2916
rect 16172 2864 16178 2916
rect 16666 2864 16672 2916
rect 16724 2864 16730 2916
rect 19030 2907 19088 2913
rect 19030 2904 19042 2907
rect 18524 2876 19042 2904
rect 11664 2808 13584 2836
rect 11664 2796 11670 2808
rect 14458 2796 14464 2848
rect 14516 2796 14522 2848
rect 16393 2839 16451 2845
rect 16393 2805 16405 2839
rect 16439 2836 16451 2839
rect 16482 2836 16488 2848
rect 16439 2808 16488 2836
rect 16439 2805 16451 2808
rect 16393 2799 16451 2805
rect 16482 2796 16488 2808
rect 16540 2796 16546 2848
rect 16942 2796 16948 2848
rect 17000 2836 17006 2848
rect 18524 2845 18552 2876
rect 19030 2873 19042 2876
rect 19076 2873 19088 2907
rect 19030 2867 19088 2873
rect 17037 2839 17095 2845
rect 17037 2836 17049 2839
rect 17000 2808 17049 2836
rect 17000 2796 17006 2808
rect 17037 2805 17049 2808
rect 17083 2805 17095 2839
rect 17037 2799 17095 2805
rect 18509 2839 18567 2845
rect 18509 2805 18521 2839
rect 18555 2805 18567 2839
rect 18509 2799 18567 2805
rect 552 2746 27576 2768
rect 552 2694 7114 2746
rect 7166 2694 7178 2746
rect 7230 2694 7242 2746
rect 7294 2694 7306 2746
rect 7358 2694 7370 2746
rect 7422 2694 13830 2746
rect 13882 2694 13894 2746
rect 13946 2694 13958 2746
rect 14010 2694 14022 2746
rect 14074 2694 14086 2746
rect 14138 2694 20546 2746
rect 20598 2694 20610 2746
rect 20662 2694 20674 2746
rect 20726 2694 20738 2746
rect 20790 2694 20802 2746
rect 20854 2694 27262 2746
rect 27314 2694 27326 2746
rect 27378 2694 27390 2746
rect 27442 2694 27454 2746
rect 27506 2694 27518 2746
rect 27570 2694 27576 2746
rect 552 2672 27576 2694
rect 3694 2592 3700 2644
rect 3752 2592 3758 2644
rect 7650 2632 7656 2644
rect 6472 2604 7656 2632
rect 6472 2573 6500 2604
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 7742 2592 7748 2644
rect 7800 2632 7806 2644
rect 7800 2604 8524 2632
rect 7800 2592 7806 2604
rect 6457 2567 6515 2573
rect 6457 2533 6469 2567
rect 6503 2533 6515 2567
rect 6457 2527 6515 2533
rect 6549 2567 6607 2573
rect 6549 2533 6561 2567
rect 6595 2564 6607 2567
rect 6638 2564 6644 2576
rect 6595 2536 6644 2564
rect 6595 2533 6607 2536
rect 6549 2527 6607 2533
rect 6638 2524 6644 2536
rect 6696 2524 6702 2576
rect 8386 2564 8392 2576
rect 7484 2536 8392 2564
rect 3602 2456 3608 2508
rect 3660 2496 3666 2508
rect 3881 2499 3939 2505
rect 3881 2496 3893 2499
rect 3660 2468 3893 2496
rect 3660 2456 3666 2468
rect 3881 2465 3893 2468
rect 3927 2465 3939 2499
rect 3881 2459 3939 2465
rect 5166 2456 5172 2508
rect 5224 2456 5230 2508
rect 5350 2456 5356 2508
rect 5408 2456 5414 2508
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 5868 2468 6377 2496
rect 5868 2456 5874 2468
rect 6365 2465 6377 2468
rect 6411 2465 6423 2499
rect 6365 2459 6423 2465
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7374 2496 7380 2508
rect 6779 2468 7380 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7374 2456 7380 2468
rect 7432 2456 7438 2508
rect 7484 2505 7512 2536
rect 8386 2524 8392 2536
rect 8444 2524 8450 2576
rect 8496 2564 8524 2604
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 14185 2635 14243 2641
rect 14185 2632 14197 2635
rect 9640 2604 14197 2632
rect 9640 2592 9646 2604
rect 14185 2601 14197 2604
rect 14231 2601 14243 2635
rect 14185 2595 14243 2601
rect 14274 2592 14280 2644
rect 14332 2632 14338 2644
rect 14645 2635 14703 2641
rect 14645 2632 14657 2635
rect 14332 2604 14657 2632
rect 14332 2592 14338 2604
rect 14645 2601 14657 2604
rect 14691 2601 14703 2635
rect 14645 2595 14703 2601
rect 16206 2592 16212 2644
rect 16264 2632 16270 2644
rect 20070 2632 20076 2644
rect 16264 2604 20076 2632
rect 16264 2592 16270 2604
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 11422 2564 11428 2576
rect 8496 2536 11428 2564
rect 11422 2524 11428 2536
rect 11480 2524 11486 2576
rect 12526 2564 12532 2576
rect 11633 2536 12532 2564
rect 7469 2499 7527 2505
rect 7469 2465 7481 2499
rect 7515 2465 7527 2499
rect 7469 2459 7527 2465
rect 7834 2456 7840 2508
rect 7892 2456 7898 2508
rect 8021 2499 8079 2505
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 8110 2496 8116 2508
rect 8067 2468 8116 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 8110 2456 8116 2468
rect 8168 2456 8174 2508
rect 8665 2499 8723 2505
rect 8665 2465 8677 2499
rect 8711 2496 8723 2499
rect 9858 2496 9864 2508
rect 8711 2468 9864 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 10502 2456 10508 2508
rect 10560 2456 10566 2508
rect 11633 2505 11661 2536
rect 12526 2524 12532 2536
rect 12584 2524 12590 2576
rect 15286 2524 15292 2576
rect 15344 2564 15350 2576
rect 15657 2567 15715 2573
rect 15657 2564 15669 2567
rect 15344 2536 15669 2564
rect 15344 2524 15350 2536
rect 15657 2533 15669 2536
rect 15703 2533 15715 2567
rect 15657 2527 15715 2533
rect 16669 2567 16727 2573
rect 16669 2533 16681 2567
rect 16715 2564 16727 2567
rect 16715 2536 17540 2564
rect 16715 2533 16727 2536
rect 16669 2527 16727 2533
rect 11609 2499 11667 2505
rect 11609 2465 11621 2499
rect 11655 2465 11667 2499
rect 11609 2459 11667 2465
rect 12434 2456 12440 2508
rect 12492 2456 12498 2508
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2496 14335 2499
rect 14366 2496 14372 2508
rect 14323 2468 14372 2496
rect 14323 2465 14335 2468
rect 14277 2459 14335 2465
rect 14366 2456 14372 2468
rect 14424 2456 14430 2508
rect 14458 2456 14464 2508
rect 14516 2456 14522 2508
rect 16393 2499 16451 2505
rect 16393 2496 16405 2499
rect 14568 2468 16405 2496
rect 6086 2388 6092 2440
rect 6144 2428 6150 2440
rect 6825 2431 6883 2437
rect 6825 2428 6837 2431
rect 6144 2400 6837 2428
rect 6144 2388 6150 2400
rect 6825 2397 6837 2400
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 7742 2428 7748 2440
rect 7607 2400 7748 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 10689 2431 10747 2437
rect 10689 2428 10701 2431
rect 9140 2400 10701 2428
rect 5350 2320 5356 2372
rect 5408 2360 5414 2372
rect 9140 2360 9168 2400
rect 10689 2397 10701 2400
rect 10735 2428 10747 2431
rect 11793 2431 11851 2437
rect 11793 2428 11805 2431
rect 10735 2400 11805 2428
rect 10735 2397 10747 2400
rect 10689 2391 10747 2397
rect 11793 2397 11805 2400
rect 11839 2428 11851 2431
rect 12253 2431 12311 2437
rect 12253 2428 12265 2431
rect 11839 2400 12265 2428
rect 11839 2397 11851 2400
rect 11793 2391 11851 2397
rect 12253 2397 12265 2400
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2428 12679 2431
rect 12710 2428 12716 2440
rect 12667 2400 12716 2428
rect 12667 2397 12679 2400
rect 12621 2391 12679 2397
rect 5408 2332 9168 2360
rect 5408 2320 5414 2332
rect 9950 2320 9956 2372
rect 10008 2360 10014 2372
rect 12268 2360 12296 2391
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2428 14151 2431
rect 14476 2428 14504 2456
rect 14139 2400 14504 2428
rect 14139 2397 14151 2400
rect 14093 2391 14151 2397
rect 14458 2360 14464 2372
rect 10008 2332 11652 2360
rect 12268 2332 14464 2360
rect 10008 2320 10014 2332
rect 4985 2295 5043 2301
rect 4985 2261 4997 2295
rect 5031 2292 5043 2295
rect 5074 2292 5080 2304
rect 5031 2264 5080 2292
rect 5031 2261 5043 2264
rect 4985 2255 5043 2261
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 6181 2295 6239 2301
rect 6181 2261 6193 2295
rect 6227 2292 6239 2295
rect 6362 2292 6368 2304
rect 6227 2264 6368 2292
rect 6227 2261 6239 2264
rect 6181 2255 6239 2261
rect 6362 2252 6368 2264
rect 6420 2252 6426 2304
rect 8478 2252 8484 2304
rect 8536 2252 8542 2304
rect 10318 2252 10324 2304
rect 10376 2252 10382 2304
rect 11425 2295 11483 2301
rect 11425 2261 11437 2295
rect 11471 2292 11483 2295
rect 11514 2292 11520 2304
rect 11471 2264 11520 2292
rect 11471 2261 11483 2264
rect 11425 2255 11483 2261
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 11624 2292 11652 2332
rect 14458 2320 14464 2332
rect 14516 2360 14522 2372
rect 14568 2360 14596 2468
rect 16393 2465 16405 2468
rect 16439 2465 16451 2499
rect 16393 2459 16451 2465
rect 16408 2428 16436 2459
rect 16482 2456 16488 2508
rect 16540 2456 16546 2508
rect 16942 2456 16948 2508
rect 17000 2456 17006 2508
rect 17512 2505 17540 2536
rect 17129 2499 17187 2505
rect 17129 2465 17141 2499
rect 17175 2496 17187 2499
rect 17221 2499 17279 2505
rect 17221 2496 17233 2499
rect 17175 2468 17233 2496
rect 17175 2465 17187 2468
rect 17129 2459 17187 2465
rect 17221 2465 17233 2468
rect 17267 2465 17279 2499
rect 17221 2459 17279 2465
rect 17497 2499 17555 2505
rect 17497 2465 17509 2499
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 19794 2456 19800 2508
rect 19852 2456 19858 2508
rect 19978 2456 19984 2508
rect 20036 2456 20042 2508
rect 20070 2456 20076 2508
rect 20128 2496 20134 2508
rect 20349 2499 20407 2505
rect 20349 2496 20361 2499
rect 20128 2468 20361 2496
rect 20128 2456 20134 2468
rect 20349 2465 20361 2468
rect 20395 2465 20407 2499
rect 20349 2459 20407 2465
rect 16761 2431 16819 2437
rect 16761 2428 16773 2431
rect 16408 2400 16773 2428
rect 16761 2397 16773 2400
rect 16807 2397 16819 2431
rect 16761 2391 16819 2397
rect 20530 2388 20536 2440
rect 20588 2388 20594 2440
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2428 21051 2431
rect 21818 2428 21824 2440
rect 21039 2400 21824 2428
rect 21039 2397 21051 2400
rect 20993 2391 21051 2397
rect 21818 2388 21824 2400
rect 21876 2388 21882 2440
rect 21450 2360 21456 2372
rect 14516 2332 14596 2360
rect 14660 2332 21456 2360
rect 14516 2320 14522 2332
rect 14660 2292 14688 2332
rect 21450 2320 21456 2332
rect 21508 2320 21514 2372
rect 11624 2264 14688 2292
rect 14734 2252 14740 2304
rect 14792 2292 14798 2304
rect 15565 2295 15623 2301
rect 15565 2292 15577 2295
rect 14792 2264 15577 2292
rect 14792 2252 14798 2264
rect 15565 2261 15577 2264
rect 15611 2292 15623 2295
rect 16114 2292 16120 2304
rect 15611 2264 16120 2292
rect 15611 2261 15623 2264
rect 15565 2255 15623 2261
rect 16114 2252 16120 2264
rect 16172 2252 16178 2304
rect 17405 2295 17463 2301
rect 17405 2261 17417 2295
rect 17451 2292 17463 2295
rect 17586 2292 17592 2304
rect 17451 2264 17592 2292
rect 17451 2261 17463 2264
rect 17405 2255 17463 2261
rect 17586 2252 17592 2264
rect 17644 2252 17650 2304
rect 17681 2295 17739 2301
rect 17681 2261 17693 2295
rect 17727 2292 17739 2295
rect 17770 2292 17776 2304
rect 17727 2264 17776 2292
rect 17727 2261 17739 2264
rect 17681 2255 17739 2261
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 552 2202 27416 2224
rect 552 2150 3756 2202
rect 3808 2150 3820 2202
rect 3872 2150 3884 2202
rect 3936 2150 3948 2202
rect 4000 2150 4012 2202
rect 4064 2150 10472 2202
rect 10524 2150 10536 2202
rect 10588 2150 10600 2202
rect 10652 2150 10664 2202
rect 10716 2150 10728 2202
rect 10780 2150 17188 2202
rect 17240 2150 17252 2202
rect 17304 2150 17316 2202
rect 17368 2150 17380 2202
rect 17432 2150 17444 2202
rect 17496 2150 23904 2202
rect 23956 2150 23968 2202
rect 24020 2150 24032 2202
rect 24084 2150 24096 2202
rect 24148 2150 24160 2202
rect 24212 2150 27416 2202
rect 552 2128 27416 2150
rect 6546 2048 6552 2100
rect 6604 2088 6610 2100
rect 7650 2088 7656 2100
rect 6604 2060 7656 2088
rect 6604 2048 6610 2060
rect 7650 2048 7656 2060
rect 7708 2048 7714 2100
rect 8294 2048 8300 2100
rect 8352 2088 8358 2100
rect 9030 2088 9036 2100
rect 8352 2060 9036 2088
rect 8352 2048 8358 2060
rect 9030 2048 9036 2060
rect 9088 2088 9094 2100
rect 9582 2088 9588 2100
rect 9088 2060 9588 2088
rect 9088 2048 9094 2060
rect 9582 2048 9588 2060
rect 9640 2088 9646 2100
rect 9769 2091 9827 2097
rect 9769 2088 9781 2091
rect 9640 2060 9781 2088
rect 9640 2048 9646 2060
rect 9769 2057 9781 2060
rect 9815 2057 9827 2091
rect 15654 2088 15660 2100
rect 9769 2051 9827 2057
rect 12406 2060 15660 2088
rect 5718 1980 5724 2032
rect 5776 2020 5782 2032
rect 5905 2023 5963 2029
rect 5905 2020 5917 2023
rect 5776 1992 5917 2020
rect 5776 1980 5782 1992
rect 5905 1989 5917 1992
rect 5951 2020 5963 2023
rect 5951 1992 7972 2020
rect 5951 1989 5963 1992
rect 5905 1983 5963 1989
rect 6730 1912 6736 1964
rect 6788 1952 6794 1964
rect 7653 1955 7711 1961
rect 6788 1924 7604 1952
rect 6788 1912 6794 1924
rect 7576 1896 7604 1924
rect 7653 1921 7665 1955
rect 7699 1952 7711 1955
rect 7742 1952 7748 1964
rect 7699 1924 7748 1952
rect 7699 1921 7711 1924
rect 7653 1915 7711 1921
rect 7742 1912 7748 1924
rect 7800 1912 7806 1964
rect 4522 1844 4528 1896
rect 4580 1844 4586 1896
rect 5350 1844 5356 1896
rect 5408 1884 5414 1896
rect 6181 1887 6239 1893
rect 6181 1884 6193 1887
rect 5408 1856 6193 1884
rect 5408 1844 5414 1856
rect 6181 1853 6193 1856
rect 6227 1853 6239 1887
rect 6181 1847 6239 1853
rect 6362 1844 6368 1896
rect 6420 1844 6426 1896
rect 6549 1887 6607 1893
rect 6549 1853 6561 1887
rect 6595 1884 6607 1887
rect 6825 1887 6883 1893
rect 6825 1884 6837 1887
rect 6595 1856 6837 1884
rect 6595 1853 6607 1856
rect 6549 1847 6607 1853
rect 6825 1853 6837 1856
rect 6871 1853 6883 1887
rect 6825 1847 6883 1853
rect 7558 1844 7564 1896
rect 7616 1844 7622 1896
rect 7944 1893 7972 1992
rect 12406 1952 12434 2060
rect 15654 2048 15660 2060
rect 15712 2048 15718 2100
rect 13722 1980 13728 2032
rect 13780 2020 13786 2032
rect 14369 2023 14427 2029
rect 13780 1992 14136 2020
rect 13780 1980 13786 1992
rect 9508 1924 12434 1952
rect 7929 1887 7987 1893
rect 7929 1853 7941 1887
rect 7975 1853 7987 1887
rect 7929 1847 7987 1853
rect 4792 1819 4850 1825
rect 4792 1785 4804 1819
rect 4838 1816 4850 1819
rect 4890 1816 4896 1828
rect 4838 1788 4896 1816
rect 4838 1785 4850 1788
rect 4792 1779 4850 1785
rect 4890 1776 4896 1788
rect 4948 1776 4954 1828
rect 6917 1819 6975 1825
rect 6917 1816 6929 1819
rect 5000 1788 6929 1816
rect 4338 1708 4344 1760
rect 4396 1748 4402 1760
rect 5000 1748 5028 1788
rect 6917 1785 6929 1788
rect 6963 1785 6975 1819
rect 6917 1779 6975 1785
rect 4396 1720 5028 1748
rect 4396 1708 4402 1720
rect 6638 1708 6644 1760
rect 6696 1708 6702 1760
rect 7944 1748 7972 1847
rect 8110 1844 8116 1896
rect 8168 1844 8174 1896
rect 8389 1887 8447 1893
rect 8389 1853 8401 1887
rect 8435 1884 8447 1887
rect 9398 1884 9404 1896
rect 8435 1856 9404 1884
rect 8435 1853 8447 1856
rect 8389 1847 8447 1853
rect 9398 1844 9404 1856
rect 9456 1844 9462 1896
rect 8478 1776 8484 1828
rect 8536 1816 8542 1828
rect 8634 1819 8692 1825
rect 8634 1816 8646 1819
rect 8536 1788 8646 1816
rect 8536 1776 8542 1788
rect 8634 1785 8646 1788
rect 8680 1785 8692 1819
rect 8634 1779 8692 1785
rect 9508 1748 9536 1924
rect 12802 1912 12808 1964
rect 12860 1952 12866 1964
rect 12860 1924 14044 1952
rect 12860 1912 12866 1924
rect 10318 1844 10324 1896
rect 10376 1884 10382 1896
rect 10413 1887 10471 1893
rect 10413 1884 10425 1887
rect 10376 1856 10425 1884
rect 10376 1844 10382 1856
rect 10413 1853 10425 1856
rect 10459 1853 10471 1887
rect 10413 1847 10471 1853
rect 11514 1844 11520 1896
rect 11572 1844 11578 1896
rect 12621 1887 12679 1893
rect 12621 1853 12633 1887
rect 12667 1884 12679 1887
rect 12710 1884 12716 1896
rect 12667 1856 12716 1884
rect 12667 1853 12679 1856
rect 12621 1847 12679 1853
rect 12710 1844 12716 1856
rect 12768 1844 12774 1896
rect 14016 1893 14044 1924
rect 13817 1887 13875 1893
rect 13817 1853 13829 1887
rect 13863 1853 13875 1887
rect 13817 1847 13875 1853
rect 14001 1887 14059 1893
rect 14001 1853 14013 1887
rect 14047 1853 14059 1887
rect 14108 1884 14136 1992
rect 14369 1989 14381 2023
rect 14415 1989 14427 2023
rect 14369 1983 14427 1989
rect 16301 2023 16359 2029
rect 16301 1989 16313 2023
rect 16347 2020 16359 2023
rect 16574 2020 16580 2032
rect 16347 1992 16580 2020
rect 16347 1989 16359 1992
rect 16301 1983 16359 1989
rect 14384 1952 14412 1983
rect 16574 1980 16580 1992
rect 16632 1980 16638 2032
rect 14384 1924 14688 1952
rect 14185 1887 14243 1893
rect 14185 1884 14197 1887
rect 14108 1856 14197 1884
rect 14001 1847 14059 1853
rect 14185 1853 14197 1856
rect 14231 1853 14243 1887
rect 14185 1847 14243 1853
rect 9674 1776 9680 1828
rect 9732 1816 9738 1828
rect 12894 1816 12900 1828
rect 9732 1788 12900 1816
rect 9732 1776 9738 1788
rect 12894 1776 12900 1788
rect 12952 1776 12958 1828
rect 7944 1720 9536 1748
rect 10226 1708 10232 1760
rect 10284 1708 10290 1760
rect 11330 1708 11336 1760
rect 11388 1708 11394 1760
rect 12802 1708 12808 1760
rect 12860 1708 12866 1760
rect 13832 1748 13860 1847
rect 14458 1844 14464 1896
rect 14516 1844 14522 1896
rect 14660 1893 14688 1924
rect 19058 1912 19064 1964
rect 19116 1952 19122 1964
rect 19429 1955 19487 1961
rect 19429 1952 19441 1955
rect 19116 1924 19441 1952
rect 19116 1912 19122 1924
rect 19429 1921 19441 1924
rect 19475 1952 19487 1955
rect 20530 1952 20536 1964
rect 19475 1924 20536 1952
rect 19475 1921 19487 1924
rect 19429 1915 19487 1921
rect 20530 1912 20536 1924
rect 20588 1952 20594 1964
rect 20717 1955 20775 1961
rect 20717 1952 20729 1955
rect 20588 1924 20729 1952
rect 20588 1912 20594 1924
rect 20717 1921 20729 1924
rect 20763 1921 20775 1955
rect 20717 1915 20775 1921
rect 14645 1887 14703 1893
rect 14645 1853 14657 1887
rect 14691 1853 14703 1887
rect 14645 1847 14703 1853
rect 14829 1887 14887 1893
rect 14829 1853 14841 1887
rect 14875 1884 14887 1887
rect 14921 1887 14979 1893
rect 14921 1884 14933 1887
rect 14875 1856 14933 1884
rect 14875 1853 14887 1856
rect 14829 1847 14887 1853
rect 14921 1853 14933 1856
rect 14967 1853 14979 1887
rect 14921 1847 14979 1853
rect 15562 1844 15568 1896
rect 15620 1884 15626 1896
rect 15749 1887 15807 1893
rect 15749 1884 15761 1887
rect 15620 1856 15761 1884
rect 15620 1844 15626 1856
rect 15749 1853 15761 1856
rect 15795 1853 15807 1887
rect 15749 1847 15807 1853
rect 15930 1844 15936 1896
rect 15988 1844 15994 1896
rect 16114 1844 16120 1896
rect 16172 1893 16178 1896
rect 16172 1884 16180 1893
rect 16172 1856 16217 1884
rect 16172 1847 16180 1856
rect 16172 1844 16178 1847
rect 17770 1844 17776 1896
rect 17828 1893 17834 1896
rect 17828 1884 17840 1893
rect 17828 1856 17873 1884
rect 17828 1847 17840 1856
rect 17828 1844 17834 1847
rect 18046 1844 18052 1896
rect 18104 1844 18110 1896
rect 18138 1844 18144 1896
rect 18196 1884 18202 1896
rect 18969 1887 19027 1893
rect 18969 1884 18981 1887
rect 18196 1856 18981 1884
rect 18196 1844 18202 1856
rect 18969 1853 18981 1856
rect 19015 1853 19027 1887
rect 18969 1847 19027 1853
rect 13906 1776 13912 1828
rect 13964 1816 13970 1828
rect 14093 1819 14151 1825
rect 14093 1816 14105 1819
rect 13964 1788 14105 1816
rect 13964 1776 13970 1788
rect 14093 1785 14105 1788
rect 14139 1785 14151 1819
rect 14093 1779 14151 1785
rect 16025 1819 16083 1825
rect 16025 1785 16037 1819
rect 16071 1816 16083 1819
rect 16390 1816 16396 1828
rect 16071 1788 16396 1816
rect 16071 1785 16083 1788
rect 16025 1779 16083 1785
rect 16390 1776 16396 1788
rect 16448 1776 16454 1828
rect 18984 1816 19012 1847
rect 19150 1844 19156 1896
rect 19208 1844 19214 1896
rect 19521 1887 19579 1893
rect 19521 1853 19533 1887
rect 19567 1884 19579 1887
rect 19702 1884 19708 1896
rect 19567 1856 19708 1884
rect 19567 1853 19579 1856
rect 19521 1847 19579 1853
rect 19702 1844 19708 1856
rect 19760 1844 19766 1896
rect 20257 1887 20315 1893
rect 20257 1884 20269 1887
rect 19812 1856 20269 1884
rect 19812 1828 19840 1856
rect 20257 1853 20269 1856
rect 20303 1853 20315 1887
rect 20257 1847 20315 1853
rect 20438 1844 20444 1896
rect 20496 1844 20502 1896
rect 20622 1844 20628 1896
rect 20680 1884 20686 1896
rect 20809 1887 20867 1893
rect 20809 1884 20821 1887
rect 20680 1856 20821 1884
rect 20680 1844 20686 1856
rect 20809 1853 20821 1856
rect 20855 1853 20867 1887
rect 20809 1847 20867 1853
rect 19794 1816 19800 1828
rect 18984 1788 19800 1816
rect 19794 1776 19800 1788
rect 19852 1776 19858 1828
rect 20165 1819 20223 1825
rect 20165 1785 20177 1819
rect 20211 1816 20223 1819
rect 27062 1816 27068 1828
rect 20211 1788 27068 1816
rect 20211 1785 20223 1788
rect 20165 1779 20223 1785
rect 27062 1776 27068 1788
rect 27120 1776 27126 1828
rect 14366 1748 14372 1760
rect 13832 1720 14372 1748
rect 14366 1708 14372 1720
rect 14424 1708 14430 1760
rect 15102 1708 15108 1760
rect 15160 1708 15166 1760
rect 15838 1708 15844 1760
rect 15896 1748 15902 1760
rect 16669 1751 16727 1757
rect 16669 1748 16681 1751
rect 15896 1720 16681 1748
rect 15896 1708 15902 1720
rect 16669 1717 16681 1720
rect 16715 1748 16727 1751
rect 17862 1748 17868 1760
rect 16715 1720 17868 1748
rect 16715 1717 16727 1720
rect 16669 1711 16727 1717
rect 17862 1708 17868 1720
rect 17920 1708 17926 1760
rect 21361 1751 21419 1757
rect 21361 1717 21373 1751
rect 21407 1748 21419 1751
rect 25314 1748 25320 1760
rect 21407 1720 25320 1748
rect 21407 1717 21419 1720
rect 21361 1711 21419 1717
rect 25314 1708 25320 1720
rect 25372 1708 25378 1760
rect 552 1658 27576 1680
rect 552 1606 7114 1658
rect 7166 1606 7178 1658
rect 7230 1606 7242 1658
rect 7294 1606 7306 1658
rect 7358 1606 7370 1658
rect 7422 1606 13830 1658
rect 13882 1606 13894 1658
rect 13946 1606 13958 1658
rect 14010 1606 14022 1658
rect 14074 1606 14086 1658
rect 14138 1606 20546 1658
rect 20598 1606 20610 1658
rect 20662 1606 20674 1658
rect 20726 1606 20738 1658
rect 20790 1606 20802 1658
rect 20854 1606 27262 1658
rect 27314 1606 27326 1658
rect 27378 1606 27390 1658
rect 27442 1606 27454 1658
rect 27506 1606 27518 1658
rect 27570 1606 27576 1658
rect 552 1584 27576 1606
rect 4890 1504 4896 1556
rect 4948 1504 4954 1556
rect 7193 1547 7251 1553
rect 7193 1513 7205 1547
rect 7239 1544 7251 1547
rect 7466 1544 7472 1556
rect 7239 1516 7472 1544
rect 7239 1513 7251 1516
rect 7193 1507 7251 1513
rect 7466 1504 7472 1516
rect 7524 1504 7530 1556
rect 9214 1504 9220 1556
rect 9272 1544 9278 1556
rect 9490 1544 9496 1556
rect 9272 1516 9496 1544
rect 9272 1504 9278 1516
rect 9490 1504 9496 1516
rect 9548 1504 9554 1556
rect 9766 1544 9772 1556
rect 9600 1516 9772 1544
rect 842 1436 848 1488
rect 900 1476 906 1488
rect 6080 1479 6138 1485
rect 900 1448 5396 1476
rect 900 1436 906 1448
rect 5074 1368 5080 1420
rect 5132 1368 5138 1420
rect 5368 1408 5396 1448
rect 6080 1445 6092 1479
rect 6126 1476 6138 1479
rect 6638 1476 6644 1488
rect 6126 1448 6644 1476
rect 6126 1445 6138 1448
rect 6080 1439 6138 1445
rect 6638 1436 6644 1448
rect 6696 1436 6702 1488
rect 8588 1448 9076 1476
rect 8588 1417 8616 1448
rect 7929 1411 7987 1417
rect 7929 1408 7941 1411
rect 5368 1380 7941 1408
rect 7929 1377 7941 1380
rect 7975 1377 7987 1411
rect 7929 1371 7987 1377
rect 8573 1411 8631 1417
rect 8573 1377 8585 1411
rect 8619 1377 8631 1411
rect 8573 1371 8631 1377
rect 8938 1368 8944 1420
rect 8996 1368 9002 1420
rect 9048 1408 9076 1448
rect 9600 1408 9628 1516
rect 9766 1504 9772 1516
rect 9824 1504 9830 1556
rect 10318 1504 10324 1556
rect 10376 1544 10382 1556
rect 10781 1547 10839 1553
rect 10781 1544 10793 1547
rect 10376 1516 10793 1544
rect 10376 1504 10382 1516
rect 10781 1513 10793 1516
rect 10827 1544 10839 1547
rect 11422 1544 11428 1556
rect 10827 1516 11428 1544
rect 10827 1513 10839 1516
rect 10781 1507 10839 1513
rect 11422 1504 11428 1516
rect 11480 1504 11486 1556
rect 12345 1547 12403 1553
rect 12345 1513 12357 1547
rect 12391 1544 12403 1547
rect 12986 1544 12992 1556
rect 12391 1516 12992 1544
rect 12391 1513 12403 1516
rect 12345 1507 12403 1513
rect 12986 1504 12992 1516
rect 13044 1504 13050 1556
rect 13909 1547 13967 1553
rect 13909 1513 13921 1547
rect 13955 1544 13967 1547
rect 14182 1544 14188 1556
rect 13955 1516 14188 1544
rect 13955 1513 13967 1516
rect 13909 1507 13967 1513
rect 14182 1504 14188 1516
rect 14240 1504 14246 1556
rect 16206 1544 16212 1556
rect 14292 1516 16212 1544
rect 9668 1479 9726 1485
rect 9668 1445 9680 1479
rect 9714 1476 9726 1479
rect 10226 1476 10232 1488
rect 9714 1448 10232 1476
rect 9714 1445 9726 1448
rect 9668 1439 9726 1445
rect 10226 1436 10232 1448
rect 10284 1436 10290 1488
rect 11232 1479 11290 1485
rect 11232 1445 11244 1479
rect 11278 1476 11290 1479
rect 11330 1476 11336 1488
rect 11278 1448 11336 1476
rect 11278 1445 11290 1448
rect 11232 1439 11290 1445
rect 11330 1436 11336 1448
rect 11388 1436 11394 1488
rect 12802 1485 12808 1488
rect 12796 1476 12808 1485
rect 12763 1448 12808 1476
rect 12796 1439 12808 1448
rect 12802 1436 12808 1439
rect 12860 1436 12866 1488
rect 12894 1436 12900 1488
rect 12952 1476 12958 1488
rect 14292 1476 14320 1516
rect 16206 1504 16212 1516
rect 16264 1504 16270 1556
rect 16301 1547 16359 1553
rect 16301 1513 16313 1547
rect 16347 1544 16359 1547
rect 16390 1544 16396 1556
rect 16347 1516 16396 1544
rect 16347 1513 16359 1516
rect 16301 1507 16359 1513
rect 16390 1504 16396 1516
rect 16448 1504 16454 1556
rect 17954 1504 17960 1556
rect 18012 1544 18018 1556
rect 18506 1544 18512 1556
rect 18012 1516 18512 1544
rect 18012 1504 18018 1516
rect 18506 1504 18512 1516
rect 18564 1504 18570 1556
rect 19058 1504 19064 1556
rect 19116 1504 19122 1556
rect 12952 1448 14320 1476
rect 12952 1436 12958 1448
rect 15102 1436 15108 1488
rect 15160 1485 15166 1488
rect 15160 1476 15172 1485
rect 17436 1479 17494 1485
rect 15160 1448 15205 1476
rect 15160 1439 15172 1448
rect 17436 1445 17448 1479
rect 17482 1476 17494 1479
rect 17586 1476 17592 1488
rect 17482 1448 17592 1476
rect 17482 1445 17494 1448
rect 17436 1439 17494 1445
rect 15160 1436 15166 1439
rect 17586 1436 17592 1448
rect 17644 1436 17650 1488
rect 19076 1476 19104 1504
rect 21450 1476 21456 1488
rect 17788 1448 20576 1476
rect 14550 1408 14556 1420
rect 9048 1380 13768 1408
rect 4522 1300 4528 1352
rect 4580 1340 4586 1352
rect 5442 1340 5448 1352
rect 4580 1312 5448 1340
rect 4580 1300 4586 1312
rect 5442 1300 5448 1312
rect 5500 1340 5506 1352
rect 5813 1343 5871 1349
rect 5813 1340 5825 1343
rect 5500 1312 5825 1340
rect 5500 1300 5506 1312
rect 5813 1309 5825 1312
rect 5859 1309 5871 1343
rect 5813 1303 5871 1309
rect 8665 1343 8723 1349
rect 8665 1309 8677 1343
rect 8711 1309 8723 1343
rect 8665 1303 8723 1309
rect 8680 1272 8708 1303
rect 8846 1300 8852 1352
rect 8904 1300 8910 1352
rect 9398 1300 9404 1352
rect 9456 1300 9462 1352
rect 10965 1343 11023 1349
rect 10965 1309 10977 1343
rect 11011 1309 11023 1343
rect 10965 1303 11023 1309
rect 12529 1343 12587 1349
rect 12529 1309 12541 1343
rect 12575 1309 12587 1343
rect 13740 1340 13768 1380
rect 14016 1380 14556 1408
rect 13906 1340 13912 1352
rect 13740 1312 13912 1340
rect 12529 1303 12587 1309
rect 9030 1272 9036 1284
rect 8680 1244 9036 1272
rect 9030 1232 9036 1244
rect 9088 1232 9094 1284
rect 9416 1204 9444 1300
rect 10980 1272 11008 1303
rect 10336 1244 11008 1272
rect 10336 1204 10364 1244
rect 9416 1176 10364 1204
rect 10980 1204 11008 1244
rect 12544 1204 12572 1303
rect 13906 1300 13912 1312
rect 13964 1300 13970 1352
rect 14016 1272 14044 1380
rect 14550 1368 14556 1380
rect 14608 1408 14614 1420
rect 15473 1411 15531 1417
rect 15473 1408 15485 1411
rect 14608 1380 15485 1408
rect 14608 1368 14614 1380
rect 15473 1377 15485 1380
rect 15519 1377 15531 1411
rect 15473 1371 15531 1377
rect 15562 1368 15568 1420
rect 15620 1408 15626 1420
rect 17788 1417 17816 1448
rect 17773 1411 17831 1417
rect 17773 1408 17785 1411
rect 15620 1380 17785 1408
rect 15620 1368 15626 1380
rect 17773 1377 17785 1380
rect 17819 1377 17831 1411
rect 17773 1371 17831 1377
rect 17954 1368 17960 1420
rect 18012 1368 18018 1420
rect 18049 1411 18107 1417
rect 18049 1377 18061 1411
rect 18095 1377 18107 1411
rect 18049 1371 18107 1377
rect 15381 1343 15439 1349
rect 15381 1309 15393 1343
rect 15427 1340 15439 1343
rect 17681 1343 17739 1349
rect 15427 1312 16574 1340
rect 15427 1309 15439 1312
rect 15381 1303 15439 1309
rect 13464 1244 14044 1272
rect 10980 1176 12572 1204
rect 12710 1164 12716 1216
rect 12768 1204 12774 1216
rect 13464 1204 13492 1244
rect 12768 1176 13492 1204
rect 14001 1207 14059 1213
rect 12768 1164 12774 1176
rect 14001 1173 14013 1207
rect 14047 1204 14059 1207
rect 14366 1204 14372 1216
rect 14047 1176 14372 1204
rect 14047 1173 14059 1176
rect 14001 1167 14059 1173
rect 14366 1164 14372 1176
rect 14424 1164 14430 1216
rect 15562 1164 15568 1216
rect 15620 1164 15626 1216
rect 16546 1204 16574 1312
rect 17681 1309 17693 1343
rect 17727 1309 17739 1343
rect 17681 1303 17739 1309
rect 17696 1272 17724 1303
rect 17862 1300 17868 1352
rect 17920 1340 17926 1352
rect 18064 1340 18092 1371
rect 18138 1368 18144 1420
rect 18196 1417 18202 1420
rect 19045 1417 19073 1448
rect 18196 1408 18204 1417
rect 19045 1411 19119 1417
rect 18196 1380 18241 1408
rect 18196 1371 18204 1380
rect 19045 1378 19073 1411
rect 19061 1377 19073 1378
rect 19107 1377 19119 1411
rect 19061 1371 19119 1377
rect 18196 1368 18202 1371
rect 19242 1368 19248 1420
rect 19300 1368 19306 1420
rect 19334 1368 19340 1420
rect 19392 1368 19398 1420
rect 19481 1411 19539 1417
rect 19481 1377 19493 1411
rect 19527 1408 19539 1411
rect 19794 1408 19800 1420
rect 19527 1380 19800 1408
rect 19527 1377 19539 1380
rect 19481 1371 19539 1377
rect 19794 1368 19800 1380
rect 19852 1368 19858 1420
rect 19886 1368 19892 1420
rect 19944 1408 19950 1420
rect 20548 1417 20576 1448
rect 20640 1448 21456 1476
rect 19981 1411 20039 1417
rect 19981 1408 19993 1411
rect 19944 1380 19993 1408
rect 19944 1368 19950 1380
rect 19981 1377 19993 1380
rect 20027 1377 20039 1411
rect 19981 1371 20039 1377
rect 20349 1411 20407 1417
rect 20349 1377 20361 1411
rect 20395 1408 20407 1411
rect 20533 1411 20591 1417
rect 20395 1380 20484 1408
rect 20395 1377 20407 1380
rect 20349 1371 20407 1377
rect 17920 1312 18092 1340
rect 20456 1340 20484 1380
rect 20533 1377 20545 1411
rect 20579 1377 20591 1411
rect 20533 1371 20591 1377
rect 20640 1340 20668 1448
rect 21450 1436 21456 1448
rect 21508 1436 21514 1488
rect 20993 1411 21051 1417
rect 20993 1377 21005 1411
rect 21039 1408 21051 1411
rect 23566 1408 23572 1420
rect 21039 1380 23572 1408
rect 21039 1377 21051 1380
rect 20993 1371 21051 1377
rect 23566 1368 23572 1380
rect 23624 1368 23630 1420
rect 20456 1312 20668 1340
rect 17920 1300 17926 1312
rect 18046 1272 18052 1284
rect 17696 1244 18052 1272
rect 17696 1204 17724 1244
rect 18046 1232 18052 1244
rect 18104 1232 18110 1284
rect 16546 1176 17724 1204
rect 18322 1164 18328 1216
rect 18380 1164 18386 1216
rect 19613 1207 19671 1213
rect 19613 1173 19625 1207
rect 19659 1204 19671 1207
rect 20070 1204 20076 1216
rect 19659 1176 20076 1204
rect 19659 1173 19671 1176
rect 19613 1167 19671 1173
rect 20070 1164 20076 1176
rect 20128 1164 20134 1216
rect 552 1114 27416 1136
rect 552 1062 3756 1114
rect 3808 1062 3820 1114
rect 3872 1062 3884 1114
rect 3936 1062 3948 1114
rect 4000 1062 4012 1114
rect 4064 1062 10472 1114
rect 10524 1062 10536 1114
rect 10588 1062 10600 1114
rect 10652 1062 10664 1114
rect 10716 1062 10728 1114
rect 10780 1062 17188 1114
rect 17240 1062 17252 1114
rect 17304 1062 17316 1114
rect 17368 1062 17380 1114
rect 17432 1062 17444 1114
rect 17496 1062 23904 1114
rect 23956 1062 23968 1114
rect 24020 1062 24032 1114
rect 24084 1062 24096 1114
rect 24148 1062 24160 1114
rect 24212 1062 27416 1114
rect 552 1040 27416 1062
rect 12406 972 13216 1000
rect 7834 892 7840 944
rect 7892 932 7898 944
rect 8481 935 8539 941
rect 8481 932 8493 935
rect 7892 904 8493 932
rect 7892 892 7898 904
rect 8481 901 8493 904
rect 8527 901 8539 935
rect 9030 932 9036 944
rect 8481 895 8539 901
rect 8588 904 9036 932
rect 7742 824 7748 876
rect 7800 864 7806 876
rect 8588 864 8616 904
rect 9030 892 9036 904
rect 9088 892 9094 944
rect 9582 892 9588 944
rect 9640 932 9646 944
rect 9953 935 10011 941
rect 9953 932 9965 935
rect 9640 904 9965 932
rect 9640 892 9646 904
rect 9953 901 9965 904
rect 9999 901 10011 935
rect 9953 895 10011 901
rect 10152 904 11008 932
rect 8846 864 8852 876
rect 7800 836 8616 864
rect 8680 836 8852 864
rect 7800 824 7806 836
rect 7650 756 7656 808
rect 7708 756 7714 808
rect 8021 799 8079 805
rect 8021 765 8033 799
rect 8067 765 8079 799
rect 8021 759 8079 765
rect 2590 688 2596 740
rect 2648 728 2654 740
rect 7009 731 7067 737
rect 7009 728 7021 731
rect 2648 700 7021 728
rect 2648 688 2654 700
rect 7009 697 7021 700
rect 7055 697 7067 731
rect 7009 691 7067 697
rect 7466 688 7472 740
rect 7524 728 7530 740
rect 8036 728 8064 759
rect 8110 756 8116 808
rect 8168 796 8174 808
rect 8680 805 8708 836
rect 8846 824 8852 836
rect 8904 864 8910 876
rect 10152 864 10180 904
rect 10318 864 10324 876
rect 8904 836 10180 864
rect 8904 824 8910 836
rect 8205 799 8263 805
rect 8205 796 8217 799
rect 8168 768 8217 796
rect 8168 756 8174 768
rect 8205 765 8217 768
rect 8251 796 8263 799
rect 8660 799 8718 805
rect 8660 796 8672 799
rect 8251 768 8672 796
rect 8251 765 8263 768
rect 8205 759 8263 765
rect 8660 765 8672 768
rect 8706 765 8718 799
rect 8660 759 8718 765
rect 8754 756 8760 808
rect 8812 756 8818 808
rect 9030 756 9036 808
rect 9088 796 9094 808
rect 10152 805 10180 836
rect 10244 836 10324 864
rect 10244 805 10272 836
rect 10318 824 10324 836
rect 10376 824 10382 876
rect 10980 864 11008 904
rect 11330 892 11336 944
rect 11388 892 11394 944
rect 12406 864 12434 972
rect 12710 892 12716 944
rect 12768 892 12774 944
rect 12986 892 12992 944
rect 13044 892 13050 944
rect 13078 892 13084 944
rect 13136 892 13142 944
rect 13188 932 13216 972
rect 14734 932 14740 944
rect 13188 904 14740 932
rect 12728 864 12756 892
rect 13004 864 13032 892
rect 10980 836 12434 864
rect 12544 836 12756 864
rect 12820 836 13032 864
rect 11532 805 11560 836
rect 10132 799 10190 805
rect 9088 768 9352 796
rect 9088 756 9094 768
rect 7524 700 8064 728
rect 8849 731 8907 737
rect 7524 688 7530 700
rect 8849 697 8861 731
rect 8895 728 8907 731
rect 9214 728 9220 740
rect 8895 700 9220 728
rect 8895 697 8907 700
rect 8849 691 8907 697
rect 9214 688 9220 700
rect 9272 688 9278 740
rect 9324 660 9352 768
rect 10132 765 10144 799
rect 10178 765 10190 799
rect 10132 759 10190 765
rect 10229 799 10287 805
rect 10229 765 10241 799
rect 10275 765 10287 799
rect 10229 759 10287 765
rect 10505 799 10563 805
rect 10505 765 10517 799
rect 10551 796 10563 799
rect 11512 799 11570 805
rect 10551 768 10640 796
rect 10551 765 10563 768
rect 10505 759 10563 765
rect 9950 688 9956 740
rect 10008 728 10014 740
rect 10321 731 10379 737
rect 10321 728 10333 731
rect 10008 700 10333 728
rect 10008 688 10014 700
rect 10321 697 10333 700
rect 10367 697 10379 731
rect 10321 691 10379 697
rect 10612 660 10640 768
rect 11512 765 11524 799
rect 11558 765 11570 799
rect 11512 759 11570 765
rect 11606 756 11612 808
rect 11664 756 11670 808
rect 12544 805 12572 836
rect 12820 805 12848 836
rect 11885 799 11943 805
rect 11885 765 11897 799
rect 11931 796 11943 799
rect 12529 799 12587 805
rect 12529 796 12541 799
rect 11931 768 12541 796
rect 11931 765 11943 768
rect 11885 759 11943 765
rect 12529 765 12541 768
rect 12575 765 12587 799
rect 12713 799 12771 805
rect 12713 796 12725 799
rect 12529 759 12587 765
rect 12636 768 12725 796
rect 11146 688 11152 740
rect 11204 728 11210 740
rect 11701 731 11759 737
rect 11701 728 11713 731
rect 11204 700 11713 728
rect 11204 688 11210 700
rect 11701 697 11713 700
rect 11747 697 11759 731
rect 11701 691 11759 697
rect 11900 660 11928 759
rect 9324 632 11928 660
rect 12636 660 12664 768
rect 12713 765 12725 768
rect 12759 765 12771 799
rect 12713 759 12771 765
rect 12805 799 12863 805
rect 12805 765 12817 799
rect 12851 765 12863 799
rect 12805 759 12863 765
rect 12949 799 13007 805
rect 12949 765 12961 799
rect 12995 796 13007 799
rect 13188 796 13216 904
rect 14734 892 14740 904
rect 14792 892 14798 944
rect 14826 892 14832 944
rect 14884 892 14890 944
rect 15562 864 15568 876
rect 14292 836 15568 864
rect 14292 805 14320 836
rect 15562 824 15568 836
rect 15620 824 15626 876
rect 12995 768 13216 796
rect 14277 799 14335 805
rect 12995 765 13007 768
rect 12949 759 13007 765
rect 14277 765 14289 799
rect 14323 765 14335 799
rect 14277 759 14335 765
rect 14366 756 14372 808
rect 14424 796 14430 808
rect 14734 805 14740 808
rect 14553 799 14611 805
rect 14553 796 14565 799
rect 14424 768 14565 796
rect 14424 756 14430 768
rect 14553 765 14565 768
rect 14599 765 14611 799
rect 14553 759 14611 765
rect 14697 799 14740 805
rect 14697 765 14709 799
rect 14697 759 14740 765
rect 14734 756 14740 759
rect 14792 756 14798 808
rect 13906 688 13912 740
rect 13964 728 13970 740
rect 14461 731 14519 737
rect 14461 728 14473 731
rect 13964 700 14473 728
rect 13964 688 13970 700
rect 14461 697 14473 700
rect 14507 697 14519 731
rect 14461 691 14519 697
rect 19702 660 19708 672
rect 12636 632 19708 660
rect 19702 620 19708 632
rect 19760 620 19766 672
rect 552 570 27576 592
rect 552 518 7114 570
rect 7166 518 7178 570
rect 7230 518 7242 570
rect 7294 518 7306 570
rect 7358 518 7370 570
rect 7422 518 13830 570
rect 13882 518 13894 570
rect 13946 518 13958 570
rect 14010 518 14022 570
rect 14074 518 14086 570
rect 14138 518 20546 570
rect 20598 518 20610 570
rect 20662 518 20674 570
rect 20726 518 20738 570
rect 20790 518 20802 570
rect 20854 518 27262 570
rect 27314 518 27326 570
rect 27378 518 27390 570
rect 27442 518 27454 570
rect 27506 518 27518 570
rect 27570 518 27576 570
rect 552 496 27576 518
<< via1 >>
rect 17500 17484 17552 17536
rect 17776 17484 17828 17536
rect 3756 17382 3808 17434
rect 3820 17382 3872 17434
rect 3884 17382 3936 17434
rect 3948 17382 4000 17434
rect 4012 17382 4064 17434
rect 10472 17382 10524 17434
rect 10536 17382 10588 17434
rect 10600 17382 10652 17434
rect 10664 17382 10716 17434
rect 10728 17382 10780 17434
rect 17188 17382 17240 17434
rect 17252 17382 17304 17434
rect 17316 17382 17368 17434
rect 17380 17382 17432 17434
rect 17444 17382 17496 17434
rect 23904 17382 23956 17434
rect 23968 17382 24020 17434
rect 24032 17382 24084 17434
rect 24096 17382 24148 17434
rect 24160 17382 24212 17434
rect 848 17323 900 17332
rect 848 17289 857 17323
rect 857 17289 891 17323
rect 891 17289 900 17323
rect 848 17280 900 17289
rect 1492 17323 1544 17332
rect 1492 17289 1501 17323
rect 1501 17289 1535 17323
rect 1535 17289 1544 17323
rect 1492 17280 1544 17289
rect 3608 17280 3660 17332
rect 5908 17280 5960 17332
rect 6552 17280 6604 17332
rect 9128 17280 9180 17332
rect 12992 17280 13044 17332
rect 14280 17280 14332 17332
rect 15568 17280 15620 17332
rect 7196 17212 7248 17264
rect 13636 17212 13688 17264
rect 14924 17212 14976 17264
rect 16580 17212 16632 17264
rect 2688 17144 2740 17196
rect 3424 17187 3476 17196
rect 3424 17153 3433 17187
rect 3433 17153 3467 17187
rect 3467 17153 3476 17187
rect 3424 17144 3476 17153
rect 4712 17187 4764 17196
rect 4712 17153 4721 17187
rect 4721 17153 4755 17187
rect 4755 17153 4764 17187
rect 4712 17144 4764 17153
rect 5264 17144 5316 17196
rect 8484 17144 8536 17196
rect 9864 17144 9916 17196
rect 5908 17076 5960 17128
rect 6000 17051 6052 17060
rect 6000 17017 6009 17051
rect 6009 17017 6043 17051
rect 6043 17017 6052 17051
rect 6000 17008 6052 17017
rect 10140 17119 10192 17128
rect 10140 17085 10149 17119
rect 10149 17085 10183 17119
rect 10183 17085 10192 17119
rect 10140 17076 10192 17085
rect 10232 17119 10284 17128
rect 10232 17085 10241 17119
rect 10241 17085 10275 17119
rect 10275 17085 10284 17119
rect 10232 17076 10284 17085
rect 25228 17144 25280 17196
rect 10692 17076 10744 17128
rect 12900 17076 12952 17128
rect 13084 17076 13136 17128
rect 13544 17076 13596 17128
rect 14372 17119 14424 17128
rect 14372 17085 14381 17119
rect 14381 17085 14415 17119
rect 14415 17085 14424 17119
rect 14372 17076 14424 17085
rect 14556 17076 14608 17128
rect 15844 17076 15896 17128
rect 15568 17008 15620 17060
rect 16212 17076 16264 17128
rect 16856 17076 16908 17128
rect 17776 17119 17828 17128
rect 17776 17085 17785 17119
rect 17785 17085 17819 17119
rect 17819 17085 17828 17119
rect 17776 17076 17828 17085
rect 19432 17076 19484 17128
rect 21640 17119 21692 17128
rect 21640 17085 21649 17119
rect 21649 17085 21683 17119
rect 21683 17085 21692 17119
rect 21640 17076 21692 17085
rect 22008 17076 22060 17128
rect 22652 17076 22704 17128
rect 23296 17076 23348 17128
rect 23756 17076 23808 17128
rect 24584 17076 24636 17128
rect 25780 17119 25832 17128
rect 25780 17085 25789 17119
rect 25789 17085 25823 17119
rect 25823 17085 25832 17119
rect 25780 17076 25832 17085
rect 26516 17076 26568 17128
rect 19524 17008 19576 17060
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 12532 16940 12584 16992
rect 14740 16983 14792 16992
rect 14740 16949 14749 16983
rect 14749 16949 14783 16983
rect 14783 16949 14792 16983
rect 14740 16940 14792 16949
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 17040 16940 17092 16992
rect 19800 16940 19852 16992
rect 20352 16940 20404 16992
rect 21456 16983 21508 16992
rect 21456 16949 21465 16983
rect 21465 16949 21499 16983
rect 21499 16949 21508 16983
rect 21456 16940 21508 16949
rect 21732 16940 21784 16992
rect 22744 16983 22796 16992
rect 22744 16949 22753 16983
rect 22753 16949 22787 16983
rect 22787 16949 22796 16983
rect 22744 16940 22796 16949
rect 24032 16983 24084 16992
rect 24032 16949 24041 16983
rect 24041 16949 24075 16983
rect 24075 16949 24084 16983
rect 24032 16940 24084 16949
rect 24676 16983 24728 16992
rect 24676 16949 24685 16983
rect 24685 16949 24719 16983
rect 24719 16949 24728 16983
rect 24676 16940 24728 16949
rect 24860 16940 24912 16992
rect 25964 16983 26016 16992
rect 25964 16949 25973 16983
rect 25973 16949 26007 16983
rect 26007 16949 26016 16983
rect 25964 16940 26016 16949
rect 26792 16983 26844 16992
rect 26792 16949 26801 16983
rect 26801 16949 26835 16983
rect 26835 16949 26844 16983
rect 26792 16940 26844 16949
rect 7114 16838 7166 16890
rect 7178 16838 7230 16890
rect 7242 16838 7294 16890
rect 7306 16838 7358 16890
rect 7370 16838 7422 16890
rect 13830 16838 13882 16890
rect 13894 16838 13946 16890
rect 13958 16838 14010 16890
rect 14022 16838 14074 16890
rect 14086 16838 14138 16890
rect 20546 16838 20598 16890
rect 20610 16838 20662 16890
rect 20674 16838 20726 16890
rect 20738 16838 20790 16890
rect 20802 16838 20854 16890
rect 27262 16838 27314 16890
rect 27326 16838 27378 16890
rect 27390 16838 27442 16890
rect 27454 16838 27506 16890
rect 27518 16838 27570 16890
rect 10140 16736 10192 16788
rect 11704 16736 11756 16788
rect 12348 16736 12400 16788
rect 14372 16736 14424 16788
rect 15384 16736 15436 16788
rect 17132 16779 17184 16788
rect 17132 16745 17141 16779
rect 17141 16745 17175 16779
rect 17175 16745 17184 16779
rect 17132 16736 17184 16745
rect 18512 16736 18564 16788
rect 19156 16736 19208 16788
rect 19984 16736 20036 16788
rect 4620 16600 4672 16652
rect 5264 16600 5316 16652
rect 9772 16668 9824 16720
rect 11152 16668 11204 16720
rect 14556 16668 14608 16720
rect 15292 16668 15344 16720
rect 6368 16643 6420 16652
rect 6368 16609 6402 16643
rect 6402 16609 6420 16643
rect 6368 16600 6420 16609
rect 7748 16643 7800 16652
rect 7748 16609 7757 16643
rect 7757 16609 7791 16643
rect 7791 16609 7800 16643
rect 7748 16600 7800 16609
rect 8484 16600 8536 16652
rect 8576 16600 8628 16652
rect 10876 16600 10928 16652
rect 11060 16600 11112 16652
rect 2044 16464 2096 16516
rect 5908 16464 5960 16516
rect 10692 16507 10744 16516
rect 10692 16473 10701 16507
rect 10701 16473 10735 16507
rect 10735 16473 10744 16507
rect 10692 16464 10744 16473
rect 10968 16464 11020 16516
rect 11244 16464 11296 16516
rect 11888 16600 11940 16652
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 12440 16643 12492 16652
rect 12440 16609 12449 16643
rect 12449 16609 12483 16643
rect 12483 16609 12492 16643
rect 12440 16600 12492 16609
rect 12624 16600 12676 16652
rect 12808 16575 12860 16584
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 12808 16532 12860 16541
rect 15200 16600 15252 16652
rect 16028 16668 16080 16720
rect 16672 16668 16724 16720
rect 19616 16668 19668 16720
rect 21548 16736 21600 16788
rect 25780 16736 25832 16788
rect 16856 16600 16908 16652
rect 19524 16643 19576 16652
rect 19524 16609 19533 16643
rect 19533 16609 19567 16643
rect 19567 16609 19576 16643
rect 19524 16600 19576 16609
rect 17684 16464 17736 16516
rect 18144 16507 18196 16516
rect 18144 16473 18153 16507
rect 18153 16473 18187 16507
rect 18187 16473 18196 16507
rect 18144 16464 18196 16473
rect 21732 16532 21784 16584
rect 24768 16643 24820 16652
rect 24768 16609 24777 16643
rect 24777 16609 24811 16643
rect 24811 16609 24820 16643
rect 24768 16600 24820 16609
rect 24860 16643 24912 16652
rect 24860 16609 24869 16643
rect 24869 16609 24903 16643
rect 24903 16609 24912 16643
rect 24860 16600 24912 16609
rect 25320 16532 25372 16584
rect 25872 16600 25924 16652
rect 26424 16643 26476 16652
rect 26424 16609 26433 16643
rect 26433 16609 26467 16643
rect 26467 16609 26476 16643
rect 26424 16600 26476 16609
rect 27068 16668 27120 16720
rect 26700 16643 26752 16652
rect 26700 16609 26709 16643
rect 26709 16609 26743 16643
rect 26743 16609 26752 16643
rect 26700 16600 26752 16609
rect 26884 16643 26936 16652
rect 26884 16609 26898 16643
rect 26898 16609 26932 16643
rect 26932 16609 26936 16643
rect 26884 16600 26936 16609
rect 26240 16532 26292 16584
rect 8024 16396 8076 16448
rect 9496 16396 9548 16448
rect 13728 16396 13780 16448
rect 21456 16464 21508 16516
rect 22744 16464 22796 16516
rect 24032 16396 24084 16448
rect 25228 16439 25280 16448
rect 25228 16405 25237 16439
rect 25237 16405 25271 16439
rect 25271 16405 25280 16439
rect 25228 16396 25280 16405
rect 25412 16396 25464 16448
rect 26976 16396 27028 16448
rect 3756 16294 3808 16346
rect 3820 16294 3872 16346
rect 3884 16294 3936 16346
rect 3948 16294 4000 16346
rect 4012 16294 4064 16346
rect 10472 16294 10524 16346
rect 10536 16294 10588 16346
rect 10600 16294 10652 16346
rect 10664 16294 10716 16346
rect 10728 16294 10780 16346
rect 17188 16294 17240 16346
rect 17252 16294 17304 16346
rect 17316 16294 17368 16346
rect 17380 16294 17432 16346
rect 17444 16294 17496 16346
rect 23904 16294 23956 16346
rect 23968 16294 24020 16346
rect 24032 16294 24084 16346
rect 24096 16294 24148 16346
rect 24160 16294 24212 16346
rect 5908 16192 5960 16244
rect 6368 16235 6420 16244
rect 6368 16201 6377 16235
rect 6377 16201 6411 16235
rect 6411 16201 6420 16235
rect 6368 16192 6420 16201
rect 8484 16192 8536 16244
rect 8024 16099 8076 16108
rect 8024 16065 8033 16099
rect 8033 16065 8067 16099
rect 8067 16065 8076 16099
rect 8024 16056 8076 16065
rect 9680 16124 9732 16176
rect 10232 16192 10284 16244
rect 10876 16192 10928 16244
rect 10968 16124 11020 16176
rect 11152 16235 11204 16244
rect 11152 16201 11161 16235
rect 11161 16201 11195 16235
rect 11195 16201 11204 16235
rect 11152 16192 11204 16201
rect 12624 16192 12676 16244
rect 9772 16056 9824 16108
rect 6644 16031 6696 16040
rect 6644 15997 6653 16031
rect 6653 15997 6687 16031
rect 6687 15997 6696 16031
rect 6644 15988 6696 15997
rect 5908 15963 5960 15972
rect 5908 15929 5917 15963
rect 5917 15929 5951 15963
rect 5951 15929 5960 15963
rect 5908 15920 5960 15929
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 7012 16031 7064 16040
rect 7012 15997 7021 16031
rect 7021 15997 7055 16031
rect 7055 15997 7064 16031
rect 7012 15988 7064 15997
rect 8852 15988 8904 16040
rect 9496 16031 9548 16040
rect 9496 15997 9505 16031
rect 9505 15997 9539 16031
rect 9539 15997 9548 16031
rect 9496 15988 9548 15997
rect 10140 16031 10192 16040
rect 10140 15997 10182 16031
rect 10182 15997 10192 16031
rect 10140 15988 10192 15997
rect 10692 16099 10744 16108
rect 10692 16065 10701 16099
rect 10701 16065 10735 16099
rect 10735 16065 10744 16099
rect 10692 16056 10744 16065
rect 10600 16031 10652 16040
rect 10600 15997 10609 16031
rect 10609 15997 10643 16031
rect 10643 15997 10652 16031
rect 10600 15988 10652 15997
rect 10876 15988 10928 16040
rect 10968 16031 11020 16040
rect 10968 15997 10977 16031
rect 10977 15997 11011 16031
rect 11011 15997 11020 16031
rect 10968 15988 11020 15997
rect 7472 15895 7524 15904
rect 7472 15861 7481 15895
rect 7481 15861 7515 15895
rect 7515 15861 7524 15895
rect 7472 15852 7524 15861
rect 11060 15920 11112 15972
rect 11244 15988 11296 16040
rect 12164 16167 12216 16176
rect 12164 16133 12173 16167
rect 12173 16133 12207 16167
rect 12207 16133 12216 16167
rect 12164 16124 12216 16133
rect 11980 16031 12032 16040
rect 11980 15997 11989 16031
rect 11989 15997 12023 16031
rect 12023 15997 12032 16031
rect 11980 15988 12032 15997
rect 12532 16031 12584 16040
rect 12532 15997 12541 16031
rect 12541 15997 12575 16031
rect 12575 15997 12584 16031
rect 12532 15988 12584 15997
rect 12716 15988 12768 16040
rect 10508 15852 10560 15904
rect 12164 15920 12216 15972
rect 13176 16235 13228 16244
rect 13176 16201 13185 16235
rect 13185 16201 13219 16235
rect 13219 16201 13228 16235
rect 13176 16192 13228 16201
rect 15200 16192 15252 16244
rect 18144 16192 18196 16244
rect 24676 16192 24728 16244
rect 12992 16099 13044 16108
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 13452 16124 13504 16176
rect 17684 16124 17736 16176
rect 25964 16124 26016 16176
rect 13728 15988 13780 16040
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 14372 16031 14424 16040
rect 14372 15997 14381 16031
rect 14381 15997 14415 16031
rect 14415 15997 14424 16031
rect 14372 15988 14424 15997
rect 23940 16056 23992 16108
rect 26792 16056 26844 16108
rect 14648 16031 14700 16040
rect 14648 15997 14657 16031
rect 14657 15997 14691 16031
rect 14691 15997 14700 16031
rect 14648 15988 14700 15997
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 15384 15988 15436 16040
rect 18788 16031 18840 16040
rect 18788 15997 18797 16031
rect 18797 15997 18831 16031
rect 18831 15997 18840 16031
rect 18788 15988 18840 15997
rect 20076 16031 20128 16040
rect 20076 15997 20085 16031
rect 20085 15997 20119 16031
rect 20119 15997 20128 16031
rect 20076 15988 20128 15997
rect 20260 16031 20312 16040
rect 20260 15997 20269 16031
rect 20269 15997 20303 16031
rect 20303 15997 20312 16031
rect 20260 15988 20312 15997
rect 21732 16031 21784 16040
rect 21732 15997 21741 16031
rect 21741 15997 21775 16031
rect 21775 15997 21784 16031
rect 21732 15988 21784 15997
rect 24492 15988 24544 16040
rect 25320 16031 25372 16040
rect 25320 15997 25329 16031
rect 25329 15997 25363 16031
rect 25363 15997 25372 16031
rect 25320 15988 25372 15997
rect 25504 16031 25556 16040
rect 25504 15997 25513 16031
rect 25513 15997 25547 16031
rect 25547 15997 25556 16031
rect 25504 15988 25556 15997
rect 26608 15988 26660 16040
rect 13176 15852 13228 15904
rect 13636 15895 13688 15904
rect 13636 15861 13645 15895
rect 13645 15861 13679 15895
rect 13679 15861 13688 15895
rect 13636 15852 13688 15861
rect 14188 15852 14240 15904
rect 19340 15895 19392 15904
rect 19340 15861 19349 15895
rect 19349 15861 19383 15895
rect 19383 15861 19392 15895
rect 19340 15852 19392 15861
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 20904 15852 20956 15904
rect 21088 15895 21140 15904
rect 21088 15861 21097 15895
rect 21097 15861 21131 15895
rect 21131 15861 21140 15895
rect 21088 15852 21140 15861
rect 24400 15895 24452 15904
rect 24400 15861 24409 15895
rect 24409 15861 24443 15895
rect 24443 15861 24452 15895
rect 24400 15852 24452 15861
rect 24952 15852 25004 15904
rect 26056 15852 26108 15904
rect 7114 15750 7166 15802
rect 7178 15750 7230 15802
rect 7242 15750 7294 15802
rect 7306 15750 7358 15802
rect 7370 15750 7422 15802
rect 13830 15750 13882 15802
rect 13894 15750 13946 15802
rect 13958 15750 14010 15802
rect 14022 15750 14074 15802
rect 14086 15750 14138 15802
rect 20546 15750 20598 15802
rect 20610 15750 20662 15802
rect 20674 15750 20726 15802
rect 20738 15750 20790 15802
rect 20802 15750 20854 15802
rect 27262 15750 27314 15802
rect 27326 15750 27378 15802
rect 27390 15750 27442 15802
rect 27454 15750 27506 15802
rect 27518 15750 27570 15802
rect 6644 15691 6696 15700
rect 6644 15657 6653 15691
rect 6653 15657 6687 15691
rect 6687 15657 6696 15691
rect 6644 15648 6696 15657
rect 6828 15648 6880 15700
rect 8852 15691 8904 15700
rect 8852 15657 8861 15691
rect 8861 15657 8895 15691
rect 8895 15657 8904 15691
rect 8852 15648 8904 15657
rect 10508 15691 10560 15700
rect 6000 15580 6052 15632
rect 8300 15580 8352 15632
rect 3424 15555 3476 15564
rect 3424 15521 3458 15555
rect 3458 15521 3476 15555
rect 3424 15512 3476 15521
rect 1400 15444 1452 15496
rect 6644 15555 6696 15564
rect 6644 15521 6653 15555
rect 6653 15521 6687 15555
rect 6687 15521 6696 15555
rect 6644 15512 6696 15521
rect 7380 15512 7432 15564
rect 6828 15444 6880 15496
rect 8484 15555 8536 15564
rect 8484 15521 8493 15555
rect 8493 15521 8527 15555
rect 8527 15521 8536 15555
rect 8484 15512 8536 15521
rect 9312 15555 9364 15564
rect 9312 15521 9321 15555
rect 9321 15521 9355 15555
rect 9355 15521 9364 15555
rect 10508 15657 10517 15691
rect 10517 15657 10551 15691
rect 10551 15657 10560 15691
rect 10508 15648 10560 15657
rect 11980 15648 12032 15700
rect 9312 15512 9364 15521
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 9772 15555 9824 15564
rect 9772 15521 9781 15555
rect 9781 15521 9815 15555
rect 9815 15521 9824 15555
rect 9772 15512 9824 15521
rect 9496 15444 9548 15496
rect 9680 15376 9732 15428
rect 9864 15376 9916 15428
rect 10508 15512 10560 15564
rect 10692 15512 10744 15564
rect 12256 15555 12308 15564
rect 12256 15521 12265 15555
rect 12265 15521 12299 15555
rect 12299 15521 12308 15555
rect 12256 15512 12308 15521
rect 14188 15648 14240 15700
rect 18788 15691 18840 15700
rect 18788 15657 18797 15691
rect 18797 15657 18831 15691
rect 18831 15657 18840 15691
rect 18788 15648 18840 15657
rect 20260 15691 20312 15700
rect 20260 15657 20269 15691
rect 20269 15657 20303 15691
rect 20303 15657 20312 15691
rect 20260 15648 20312 15657
rect 14372 15580 14424 15632
rect 18880 15580 18932 15632
rect 19432 15580 19484 15632
rect 22836 15648 22888 15700
rect 24492 15648 24544 15700
rect 25780 15648 25832 15700
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 13636 15512 13688 15564
rect 16212 15512 16264 15564
rect 16396 15555 16448 15564
rect 16396 15521 16405 15555
rect 16405 15521 16439 15555
rect 16439 15521 16448 15555
rect 16396 15512 16448 15521
rect 16672 15555 16724 15564
rect 12808 15444 12860 15496
rect 16672 15521 16680 15555
rect 16680 15521 16714 15555
rect 16714 15521 16724 15555
rect 16672 15512 16724 15521
rect 16764 15555 16816 15564
rect 16764 15521 16773 15555
rect 16773 15521 16807 15555
rect 16807 15521 16816 15555
rect 16764 15512 16816 15521
rect 18696 15512 18748 15564
rect 19892 15512 19944 15564
rect 20168 15512 20220 15564
rect 16948 15444 17000 15496
rect 4252 15308 4304 15360
rect 6644 15308 6696 15360
rect 8944 15308 8996 15360
rect 9772 15308 9824 15360
rect 15200 15308 15252 15360
rect 20444 15444 20496 15496
rect 21088 15512 21140 15564
rect 22652 15580 22704 15632
rect 22560 15512 22612 15564
rect 22928 15555 22980 15564
rect 22928 15521 22932 15555
rect 22932 15521 22966 15555
rect 22966 15521 22980 15555
rect 22928 15512 22980 15521
rect 23112 15555 23164 15564
rect 23112 15521 23121 15555
rect 23121 15521 23155 15555
rect 23155 15521 23164 15555
rect 23112 15512 23164 15521
rect 25228 15580 25280 15632
rect 23388 15555 23440 15564
rect 23388 15521 23397 15555
rect 23397 15521 23431 15555
rect 23431 15521 23440 15555
rect 23388 15512 23440 15521
rect 23572 15512 23624 15564
rect 23940 15555 23992 15564
rect 23940 15521 23949 15555
rect 23949 15521 23983 15555
rect 23983 15521 23992 15555
rect 23940 15512 23992 15521
rect 24860 15512 24912 15564
rect 23480 15444 23532 15496
rect 17776 15308 17828 15360
rect 21732 15308 21784 15360
rect 22744 15351 22796 15360
rect 22744 15317 22753 15351
rect 22753 15317 22787 15351
rect 22787 15317 22796 15351
rect 22744 15308 22796 15317
rect 24676 15308 24728 15360
rect 25780 15308 25832 15360
rect 3756 15206 3808 15258
rect 3820 15206 3872 15258
rect 3884 15206 3936 15258
rect 3948 15206 4000 15258
rect 4012 15206 4064 15258
rect 10472 15206 10524 15258
rect 10536 15206 10588 15258
rect 10600 15206 10652 15258
rect 10664 15206 10716 15258
rect 10728 15206 10780 15258
rect 17188 15206 17240 15258
rect 17252 15206 17304 15258
rect 17316 15206 17368 15258
rect 17380 15206 17432 15258
rect 17444 15206 17496 15258
rect 23904 15206 23956 15258
rect 23968 15206 24020 15258
rect 24032 15206 24084 15258
rect 24096 15206 24148 15258
rect 24160 15206 24212 15258
rect 4804 15104 4856 15156
rect 5264 15104 5316 15156
rect 1400 14900 1452 14952
rect 4252 14900 4304 14952
rect 4344 14832 4396 14884
rect 3792 14764 3844 14816
rect 6000 15147 6052 15156
rect 6000 15113 6009 15147
rect 6009 15113 6043 15147
rect 6043 15113 6052 15147
rect 6000 15104 6052 15113
rect 9312 15104 9364 15156
rect 9680 15104 9732 15156
rect 10324 15036 10376 15088
rect 5356 14943 5408 14952
rect 5356 14909 5365 14943
rect 5365 14909 5399 14943
rect 5399 14909 5408 14943
rect 5356 14900 5408 14909
rect 5540 14943 5592 14952
rect 5540 14909 5549 14943
rect 5549 14909 5583 14943
rect 5583 14909 5592 14943
rect 5540 14900 5592 14909
rect 5080 14875 5132 14884
rect 5080 14841 5089 14875
rect 5089 14841 5123 14875
rect 5123 14841 5132 14875
rect 5080 14832 5132 14841
rect 6644 14943 6696 14952
rect 6644 14909 6653 14943
rect 6653 14909 6687 14943
rect 6687 14909 6696 14943
rect 6644 14900 6696 14909
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 8208 14832 8260 14884
rect 8300 14832 8352 14884
rect 9496 14900 9548 14952
rect 9956 14943 10008 14952
rect 9956 14909 9965 14943
rect 9965 14909 9999 14943
rect 9999 14909 10008 14943
rect 9956 14900 10008 14909
rect 10876 15104 10928 15156
rect 12532 15104 12584 15156
rect 12256 15036 12308 15088
rect 16764 15104 16816 15156
rect 18604 15104 18656 15156
rect 18696 15147 18748 15156
rect 18696 15113 18705 15147
rect 18705 15113 18739 15147
rect 18739 15113 18748 15147
rect 18696 15104 18748 15113
rect 16212 14968 16264 15020
rect 12440 14900 12492 14952
rect 12992 14900 13044 14952
rect 14188 14900 14240 14952
rect 15936 14900 15988 14952
rect 18052 14900 18104 14952
rect 10324 14832 10376 14884
rect 5816 14764 5868 14816
rect 6460 14807 6512 14816
rect 6460 14773 6469 14807
rect 6469 14773 6503 14807
rect 6503 14773 6512 14807
rect 6460 14764 6512 14773
rect 6736 14807 6788 14816
rect 6736 14773 6745 14807
rect 6745 14773 6779 14807
rect 6779 14773 6788 14807
rect 6736 14764 6788 14773
rect 8576 14764 8628 14816
rect 9128 14764 9180 14816
rect 9220 14807 9272 14816
rect 9220 14773 9229 14807
rect 9229 14773 9263 14807
rect 9263 14773 9272 14807
rect 9220 14764 9272 14773
rect 9588 14764 9640 14816
rect 15292 14832 15344 14884
rect 17684 14832 17736 14884
rect 15660 14764 15712 14816
rect 16672 14764 16724 14816
rect 17224 14764 17276 14816
rect 18144 14875 18196 14884
rect 18144 14841 18153 14875
rect 18153 14841 18187 14875
rect 18187 14841 18196 14875
rect 18144 14832 18196 14841
rect 19340 15036 19392 15088
rect 18788 14968 18840 15020
rect 18604 14900 18656 14952
rect 19524 15011 19576 15020
rect 19524 14977 19533 15011
rect 19533 14977 19567 15011
rect 19567 14977 19576 15011
rect 19524 14968 19576 14977
rect 19064 14943 19116 14952
rect 19064 14909 19073 14943
rect 19073 14909 19107 14943
rect 19107 14909 19116 14943
rect 19064 14900 19116 14909
rect 19892 14900 19944 14952
rect 20260 14900 20312 14952
rect 24492 15147 24544 15156
rect 24492 15113 24501 15147
rect 24501 15113 24535 15147
rect 24535 15113 24544 15147
rect 24492 15104 24544 15113
rect 24032 15036 24084 15088
rect 26976 15104 27028 15156
rect 20904 14968 20956 15020
rect 20812 14943 20864 14952
rect 20812 14909 20821 14943
rect 20821 14909 20855 14943
rect 20855 14909 20864 14943
rect 20812 14900 20864 14909
rect 23480 14968 23532 15020
rect 19340 14764 19392 14816
rect 21180 14832 21232 14884
rect 22008 14832 22060 14884
rect 24676 14900 24728 14952
rect 25964 14900 26016 14952
rect 25780 14832 25832 14884
rect 23204 14807 23256 14816
rect 23204 14773 23213 14807
rect 23213 14773 23247 14807
rect 23247 14773 23256 14807
rect 23204 14764 23256 14773
rect 25136 14764 25188 14816
rect 25872 14764 25924 14816
rect 7114 14662 7166 14714
rect 7178 14662 7230 14714
rect 7242 14662 7294 14714
rect 7306 14662 7358 14714
rect 7370 14662 7422 14714
rect 13830 14662 13882 14714
rect 13894 14662 13946 14714
rect 13958 14662 14010 14714
rect 14022 14662 14074 14714
rect 14086 14662 14138 14714
rect 20546 14662 20598 14714
rect 20610 14662 20662 14714
rect 20674 14662 20726 14714
rect 20738 14662 20790 14714
rect 20802 14662 20854 14714
rect 27262 14662 27314 14714
rect 27326 14662 27378 14714
rect 27390 14662 27442 14714
rect 27454 14662 27506 14714
rect 27518 14662 27570 14714
rect 3424 14560 3476 14612
rect 4344 14560 4396 14612
rect 3240 14424 3292 14476
rect 3792 14467 3844 14476
rect 3792 14433 3801 14467
rect 3801 14433 3835 14467
rect 3835 14433 3844 14467
rect 3792 14424 3844 14433
rect 4160 14467 4212 14476
rect 4160 14433 4169 14467
rect 4169 14433 4203 14467
rect 4203 14433 4212 14467
rect 4160 14424 4212 14433
rect 5264 14560 5316 14612
rect 5356 14603 5408 14612
rect 5356 14569 5365 14603
rect 5365 14569 5399 14603
rect 5399 14569 5408 14603
rect 5356 14560 5408 14569
rect 6460 14560 6512 14612
rect 9864 14560 9916 14612
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 11060 14560 11112 14612
rect 4804 14467 4856 14476
rect 4804 14433 4813 14467
rect 4813 14433 4847 14467
rect 4847 14433 4856 14467
rect 4804 14424 4856 14433
rect 5540 14492 5592 14544
rect 6000 14492 6052 14544
rect 6828 14492 6880 14544
rect 7564 14492 7616 14544
rect 8484 14492 8536 14544
rect 8852 14535 8904 14544
rect 8852 14501 8886 14535
rect 8886 14501 8904 14535
rect 8852 14492 8904 14501
rect 1400 14356 1452 14408
rect 6276 14424 6328 14476
rect 8576 14467 8628 14476
rect 8576 14433 8585 14467
rect 8585 14433 8619 14467
rect 8619 14433 8628 14467
rect 8576 14424 8628 14433
rect 5356 14356 5408 14408
rect 7012 14356 7064 14408
rect 7472 14356 7524 14408
rect 9864 14424 9916 14476
rect 10048 14492 10100 14544
rect 13268 14492 13320 14544
rect 12164 14424 12216 14476
rect 15200 14492 15252 14544
rect 3056 14263 3108 14272
rect 3056 14229 3065 14263
rect 3065 14229 3099 14263
rect 3099 14229 3108 14263
rect 3056 14220 3108 14229
rect 3424 14220 3476 14272
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 8392 14263 8444 14272
rect 8392 14229 8401 14263
rect 8401 14229 8435 14263
rect 8435 14229 8444 14263
rect 8392 14220 8444 14229
rect 8760 14220 8812 14272
rect 8944 14220 8996 14272
rect 11336 14356 11388 14408
rect 11888 14356 11940 14408
rect 14464 14467 14516 14476
rect 14464 14433 14473 14467
rect 14473 14433 14507 14467
rect 14507 14433 14516 14467
rect 14464 14424 14516 14433
rect 15108 14399 15160 14408
rect 15108 14365 15117 14399
rect 15117 14365 15151 14399
rect 15151 14365 15160 14399
rect 15108 14356 15160 14365
rect 10232 14220 10284 14272
rect 12256 14263 12308 14272
rect 12256 14229 12265 14263
rect 12265 14229 12299 14263
rect 12299 14229 12308 14263
rect 12256 14220 12308 14229
rect 13820 14263 13872 14272
rect 13820 14229 13829 14263
rect 13829 14229 13863 14263
rect 13863 14229 13872 14263
rect 13820 14220 13872 14229
rect 15660 14467 15712 14476
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 15936 14603 15988 14612
rect 15936 14569 15945 14603
rect 15945 14569 15979 14603
rect 15979 14569 15988 14603
rect 15936 14560 15988 14569
rect 16396 14560 16448 14612
rect 19524 14560 19576 14612
rect 20076 14603 20128 14612
rect 20076 14569 20085 14603
rect 20085 14569 20119 14603
rect 20119 14569 20128 14603
rect 20076 14560 20128 14569
rect 20168 14560 20220 14612
rect 20720 14560 20772 14612
rect 18052 14492 18104 14544
rect 17224 14424 17276 14476
rect 20168 14424 20220 14476
rect 20904 14492 20956 14544
rect 21180 14492 21232 14544
rect 22560 14560 22612 14612
rect 24860 14560 24912 14612
rect 25504 14560 25556 14612
rect 23112 14535 23164 14544
rect 20444 14467 20496 14476
rect 20444 14433 20453 14467
rect 20453 14433 20487 14467
rect 20487 14433 20496 14467
rect 20444 14424 20496 14433
rect 16488 14356 16540 14408
rect 17868 14399 17920 14408
rect 17868 14365 17877 14399
rect 17877 14365 17911 14399
rect 17911 14365 17920 14399
rect 17868 14356 17920 14365
rect 19892 14399 19944 14408
rect 19892 14365 19901 14399
rect 19901 14365 19935 14399
rect 19935 14365 19944 14399
rect 19892 14356 19944 14365
rect 20720 14467 20772 14476
rect 20720 14433 20729 14467
rect 20729 14433 20763 14467
rect 20763 14433 20772 14467
rect 20720 14424 20772 14433
rect 20996 14424 21048 14476
rect 21548 14467 21600 14476
rect 21548 14433 21557 14467
rect 21557 14433 21591 14467
rect 21591 14433 21600 14467
rect 21548 14424 21600 14433
rect 21640 14356 21692 14408
rect 21824 14467 21876 14476
rect 21824 14433 21832 14467
rect 21832 14433 21866 14467
rect 21866 14433 21876 14467
rect 21824 14424 21876 14433
rect 21916 14467 21968 14476
rect 21916 14433 21925 14467
rect 21925 14433 21959 14467
rect 21959 14433 21968 14467
rect 21916 14424 21968 14433
rect 23112 14501 23121 14535
rect 23121 14501 23155 14535
rect 23155 14501 23164 14535
rect 23112 14492 23164 14501
rect 23664 14492 23716 14544
rect 22928 14467 22980 14476
rect 22928 14433 22932 14467
rect 22932 14433 22966 14467
rect 22966 14433 22980 14467
rect 22928 14424 22980 14433
rect 23020 14467 23072 14476
rect 23020 14433 23029 14467
rect 23029 14433 23063 14467
rect 23063 14433 23072 14467
rect 23020 14424 23072 14433
rect 23204 14467 23256 14476
rect 23204 14433 23249 14467
rect 23249 14433 23256 14467
rect 23204 14424 23256 14433
rect 23388 14467 23440 14476
rect 23388 14433 23397 14467
rect 23397 14433 23431 14467
rect 23431 14433 23440 14467
rect 23388 14424 23440 14433
rect 23756 14424 23808 14476
rect 24032 14467 24084 14476
rect 24032 14433 24041 14467
rect 24041 14433 24075 14467
rect 24075 14433 24084 14467
rect 24032 14424 24084 14433
rect 19064 14220 19116 14272
rect 22008 14399 22060 14408
rect 22008 14365 22017 14399
rect 22017 14365 22051 14399
rect 22051 14365 22060 14399
rect 22008 14356 22060 14365
rect 22284 14356 22336 14408
rect 24400 14424 24452 14476
rect 22836 14220 22888 14272
rect 24768 14356 24820 14408
rect 24952 14467 25004 14476
rect 24952 14433 24961 14467
rect 24961 14433 24995 14467
rect 24995 14433 25004 14467
rect 24952 14424 25004 14433
rect 25044 14467 25096 14476
rect 25044 14433 25053 14467
rect 25053 14433 25087 14467
rect 25087 14433 25096 14467
rect 25044 14424 25096 14433
rect 26240 14560 26292 14612
rect 26332 14492 26384 14544
rect 25320 14424 25372 14476
rect 25504 14467 25556 14476
rect 25504 14433 25508 14467
rect 25508 14433 25542 14467
rect 25542 14433 25556 14467
rect 25504 14424 25556 14433
rect 25136 14356 25188 14408
rect 23664 14288 23716 14340
rect 26424 14467 26476 14476
rect 26424 14433 26433 14467
rect 26433 14433 26467 14467
rect 26467 14433 26476 14467
rect 26424 14424 26476 14433
rect 26608 14467 26660 14476
rect 26608 14433 26615 14467
rect 26615 14433 26660 14467
rect 26608 14424 26660 14433
rect 26700 14467 26752 14476
rect 26700 14433 26709 14467
rect 26709 14433 26743 14467
rect 26743 14433 26752 14467
rect 26700 14424 26752 14433
rect 26792 14467 26844 14476
rect 26792 14433 26801 14467
rect 26801 14433 26835 14467
rect 26835 14433 26844 14467
rect 26792 14424 26844 14433
rect 26884 14467 26936 14476
rect 26884 14433 26898 14467
rect 26898 14433 26932 14467
rect 26932 14433 26936 14467
rect 26884 14424 26936 14433
rect 24584 14263 24636 14272
rect 24584 14229 24593 14263
rect 24593 14229 24627 14263
rect 24627 14229 24636 14263
rect 24584 14220 24636 14229
rect 25872 14288 25924 14340
rect 26516 14220 26568 14272
rect 3756 14118 3808 14170
rect 3820 14118 3872 14170
rect 3884 14118 3936 14170
rect 3948 14118 4000 14170
rect 4012 14118 4064 14170
rect 10472 14118 10524 14170
rect 10536 14118 10588 14170
rect 10600 14118 10652 14170
rect 10664 14118 10716 14170
rect 10728 14118 10780 14170
rect 17188 14118 17240 14170
rect 17252 14118 17304 14170
rect 17316 14118 17368 14170
rect 17380 14118 17432 14170
rect 17444 14118 17496 14170
rect 23904 14118 23956 14170
rect 23968 14118 24020 14170
rect 24032 14118 24084 14170
rect 24096 14118 24148 14170
rect 24160 14118 24212 14170
rect 3240 14059 3292 14068
rect 3240 14025 3249 14059
rect 3249 14025 3283 14059
rect 3283 14025 3292 14059
rect 3240 14016 3292 14025
rect 4436 14016 4488 14068
rect 5816 14016 5868 14068
rect 8208 14016 8260 14068
rect 11336 14016 11388 14068
rect 3332 13948 3384 14000
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 4344 13991 4396 14000
rect 4344 13957 4353 13991
rect 4353 13957 4387 13991
rect 4387 13957 4396 13991
rect 4344 13948 4396 13957
rect 4528 13880 4580 13932
rect 5080 13923 5132 13932
rect 5080 13889 5089 13923
rect 5089 13889 5123 13923
rect 5123 13889 5132 13923
rect 5080 13880 5132 13889
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 4252 13812 4304 13864
rect 3056 13744 3108 13796
rect 4528 13787 4580 13796
rect 4068 13719 4120 13728
rect 4068 13685 4093 13719
rect 4093 13685 4120 13719
rect 4528 13753 4539 13787
rect 4539 13753 4580 13787
rect 4528 13744 4580 13753
rect 5264 13855 5316 13864
rect 5264 13821 5273 13855
rect 5273 13821 5307 13855
rect 5307 13821 5316 13855
rect 5264 13812 5316 13821
rect 5632 13855 5684 13864
rect 5632 13821 5641 13855
rect 5641 13821 5675 13855
rect 5675 13821 5684 13855
rect 5632 13812 5684 13821
rect 6000 13812 6052 13864
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 7748 13880 7800 13932
rect 9404 13880 9456 13932
rect 12808 14016 12860 14068
rect 15108 14016 15160 14068
rect 16488 14059 16540 14068
rect 16488 14025 16497 14059
rect 16497 14025 16531 14059
rect 16531 14025 16540 14059
rect 16488 14016 16540 14025
rect 17500 14016 17552 14068
rect 18788 14016 18840 14068
rect 21640 14016 21692 14068
rect 22284 14059 22336 14068
rect 22284 14025 22293 14059
rect 22293 14025 22327 14059
rect 22327 14025 22336 14059
rect 22284 14016 22336 14025
rect 18144 13948 18196 14000
rect 12808 13880 12860 13932
rect 6276 13855 6328 13864
rect 6276 13821 6285 13855
rect 6285 13821 6319 13855
rect 6319 13821 6328 13855
rect 6276 13812 6328 13821
rect 8668 13855 8720 13864
rect 8668 13821 8702 13855
rect 8702 13821 8720 13855
rect 8668 13812 8720 13821
rect 9588 13812 9640 13864
rect 8208 13744 8260 13796
rect 10324 13812 10376 13864
rect 12256 13812 12308 13864
rect 13820 13855 13872 13864
rect 13820 13821 13854 13855
rect 13854 13821 13872 13855
rect 13820 13812 13872 13821
rect 15200 13812 15252 13864
rect 17868 13812 17920 13864
rect 4068 13676 4120 13685
rect 6644 13676 6696 13728
rect 8760 13676 8812 13728
rect 9404 13676 9456 13728
rect 9496 13676 9548 13728
rect 14372 13744 14424 13796
rect 16120 13744 16172 13796
rect 21548 13948 21600 14000
rect 19708 13812 19760 13864
rect 20168 13855 20220 13864
rect 20168 13821 20177 13855
rect 20177 13821 20211 13855
rect 20211 13821 20220 13855
rect 20168 13812 20220 13821
rect 21088 13812 21140 13864
rect 23204 14016 23256 14068
rect 23388 14016 23440 14068
rect 26424 14016 26476 14068
rect 26608 14016 26660 14068
rect 22836 13880 22888 13932
rect 24584 13948 24636 14000
rect 24860 13880 24912 13932
rect 22744 13855 22796 13864
rect 22744 13821 22753 13855
rect 22753 13821 22787 13855
rect 22787 13821 22796 13855
rect 22744 13812 22796 13821
rect 18236 13744 18288 13796
rect 19432 13744 19484 13796
rect 20996 13744 21048 13796
rect 23756 13812 23808 13864
rect 24584 13855 24636 13864
rect 24584 13821 24593 13855
rect 24593 13821 24627 13855
rect 24627 13821 24636 13855
rect 24584 13812 24636 13821
rect 24676 13812 24728 13864
rect 26056 13812 26108 13864
rect 25872 13744 25924 13796
rect 13176 13676 13228 13728
rect 14280 13676 14332 13728
rect 16212 13676 16264 13728
rect 18788 13676 18840 13728
rect 19708 13676 19760 13728
rect 20904 13676 20956 13728
rect 22192 13719 22244 13728
rect 22192 13685 22201 13719
rect 22201 13685 22235 13719
rect 22235 13685 22244 13719
rect 22192 13676 22244 13685
rect 23848 13719 23900 13728
rect 23848 13685 23857 13719
rect 23857 13685 23891 13719
rect 23891 13685 23900 13719
rect 23848 13676 23900 13685
rect 25688 13676 25740 13728
rect 7114 13574 7166 13626
rect 7178 13574 7230 13626
rect 7242 13574 7294 13626
rect 7306 13574 7358 13626
rect 7370 13574 7422 13626
rect 13830 13574 13882 13626
rect 13894 13574 13946 13626
rect 13958 13574 14010 13626
rect 14022 13574 14074 13626
rect 14086 13574 14138 13626
rect 20546 13574 20598 13626
rect 20610 13574 20662 13626
rect 20674 13574 20726 13626
rect 20738 13574 20790 13626
rect 20802 13574 20854 13626
rect 27262 13574 27314 13626
rect 27326 13574 27378 13626
rect 27390 13574 27442 13626
rect 27454 13574 27506 13626
rect 27518 13574 27570 13626
rect 4160 13472 4212 13524
rect 4252 13515 4304 13524
rect 4252 13481 4261 13515
rect 4261 13481 4295 13515
rect 4295 13481 4304 13515
rect 4252 13472 4304 13481
rect 3516 13404 3568 13456
rect 4712 13472 4764 13524
rect 5264 13472 5316 13524
rect 6276 13515 6328 13524
rect 6276 13481 6285 13515
rect 6285 13481 6319 13515
rect 6319 13481 6328 13515
rect 6276 13472 6328 13481
rect 8484 13472 8536 13524
rect 8668 13472 8720 13524
rect 8852 13472 8904 13524
rect 3792 13379 3844 13388
rect 3792 13345 3801 13379
rect 3801 13345 3835 13379
rect 3835 13345 3844 13379
rect 3792 13336 3844 13345
rect 3240 13311 3292 13320
rect 3240 13277 3249 13311
rect 3249 13277 3283 13311
rect 3283 13277 3292 13311
rect 3240 13268 3292 13277
rect 4344 13336 4396 13388
rect 4804 13447 4856 13456
rect 4804 13413 4813 13447
rect 4813 13413 4847 13447
rect 4847 13413 4856 13447
rect 4804 13404 4856 13413
rect 5632 13404 5684 13456
rect 6552 13404 6604 13456
rect 8392 13404 8444 13456
rect 4068 13268 4120 13320
rect 6276 13379 6328 13388
rect 6276 13345 6285 13379
rect 6285 13345 6319 13379
rect 6319 13345 6328 13379
rect 6276 13336 6328 13345
rect 6736 13336 6788 13388
rect 7012 13268 7064 13320
rect 4160 13200 4212 13252
rect 4344 13200 4396 13252
rect 2044 13132 2096 13184
rect 4988 13132 5040 13184
rect 5816 13200 5868 13252
rect 7564 13336 7616 13388
rect 8576 13336 8628 13388
rect 8852 13379 8904 13388
rect 8852 13345 8861 13379
rect 8861 13345 8895 13379
rect 8895 13345 8904 13379
rect 8852 13336 8904 13345
rect 9588 13404 9640 13456
rect 11888 13515 11940 13524
rect 11888 13481 11897 13515
rect 11897 13481 11931 13515
rect 11931 13481 11940 13515
rect 11888 13472 11940 13481
rect 9220 13379 9272 13388
rect 9220 13345 9229 13379
rect 9229 13345 9263 13379
rect 9263 13345 9272 13379
rect 9220 13336 9272 13345
rect 9404 13379 9456 13388
rect 9404 13345 9413 13379
rect 9413 13345 9447 13379
rect 9447 13345 9456 13379
rect 9404 13336 9456 13345
rect 7932 13268 7984 13320
rect 8300 13311 8352 13320
rect 8300 13277 8309 13311
rect 8309 13277 8343 13311
rect 8343 13277 8352 13311
rect 8300 13268 8352 13277
rect 8760 13268 8812 13320
rect 11980 13404 12032 13456
rect 9864 13336 9916 13388
rect 10232 13336 10284 13388
rect 12164 13379 12216 13388
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 9404 13200 9456 13252
rect 13176 13379 13228 13388
rect 13176 13345 13185 13379
rect 13185 13345 13219 13379
rect 13219 13345 13228 13379
rect 13176 13336 13228 13345
rect 14280 13472 14332 13524
rect 14372 13447 14424 13456
rect 14372 13413 14381 13447
rect 14381 13413 14415 13447
rect 14415 13413 14424 13447
rect 14372 13404 14424 13413
rect 14280 13379 14332 13388
rect 14280 13345 14289 13379
rect 14289 13345 14323 13379
rect 14323 13345 14332 13379
rect 14280 13336 14332 13345
rect 15108 13404 15160 13456
rect 16120 13515 16172 13524
rect 16120 13481 16129 13515
rect 16129 13481 16163 13515
rect 16163 13481 16172 13515
rect 16120 13472 16172 13481
rect 16948 13472 17000 13524
rect 17684 13472 17736 13524
rect 17776 13472 17828 13524
rect 12716 13268 12768 13320
rect 14464 13268 14516 13320
rect 6276 13132 6328 13184
rect 8024 13132 8076 13184
rect 8208 13132 8260 13184
rect 9772 13132 9824 13184
rect 16396 13379 16448 13388
rect 16396 13345 16405 13379
rect 16405 13345 16439 13379
rect 16439 13345 16448 13379
rect 16396 13336 16448 13345
rect 14740 13311 14792 13320
rect 14740 13277 14749 13311
rect 14749 13277 14783 13311
rect 14783 13277 14792 13311
rect 14740 13268 14792 13277
rect 14924 13268 14976 13320
rect 16580 13379 16632 13388
rect 16580 13345 16589 13379
rect 16589 13345 16623 13379
rect 16623 13345 16632 13379
rect 16580 13336 16632 13345
rect 16764 13379 16816 13388
rect 16764 13345 16773 13379
rect 16773 13345 16807 13379
rect 16807 13345 16816 13379
rect 16764 13336 16816 13345
rect 19892 13472 19944 13524
rect 21088 13472 21140 13524
rect 21548 13472 21600 13524
rect 22928 13472 22980 13524
rect 23572 13472 23624 13524
rect 24584 13472 24636 13524
rect 25964 13515 26016 13524
rect 25964 13481 25973 13515
rect 25973 13481 26007 13515
rect 26007 13481 26016 13515
rect 25964 13472 26016 13481
rect 16948 13268 17000 13320
rect 16672 13200 16724 13252
rect 16764 13200 16816 13252
rect 17684 13379 17736 13388
rect 17684 13345 17693 13379
rect 17693 13345 17727 13379
rect 17727 13345 17736 13379
rect 17684 13336 17736 13345
rect 18788 13404 18840 13456
rect 18236 13379 18288 13391
rect 18236 13345 18268 13379
rect 18268 13345 18288 13379
rect 18236 13339 18288 13345
rect 18420 13379 18472 13388
rect 18420 13345 18427 13379
rect 18427 13345 18472 13379
rect 17592 13268 17644 13320
rect 18420 13336 18472 13345
rect 17960 13268 18012 13320
rect 18604 13379 18656 13388
rect 18604 13345 18613 13379
rect 18613 13345 18647 13379
rect 18647 13345 18656 13379
rect 18604 13336 18656 13345
rect 18696 13379 18748 13388
rect 18696 13345 18710 13379
rect 18710 13345 18744 13379
rect 18744 13345 18748 13379
rect 18696 13336 18748 13345
rect 19248 13379 19300 13388
rect 19248 13345 19257 13379
rect 19257 13345 19291 13379
rect 19291 13345 19300 13379
rect 19248 13336 19300 13345
rect 19340 13379 19392 13388
rect 19340 13345 19349 13379
rect 19349 13345 19383 13379
rect 19383 13345 19392 13379
rect 19340 13336 19392 13345
rect 19432 13268 19484 13320
rect 20076 13379 20128 13388
rect 20076 13345 20085 13379
rect 20085 13345 20119 13379
rect 20119 13345 20128 13379
rect 20076 13336 20128 13345
rect 20168 13379 20220 13388
rect 20168 13345 20177 13379
rect 20177 13345 20211 13379
rect 20211 13345 20220 13379
rect 20168 13336 20220 13345
rect 20904 13404 20956 13456
rect 22192 13404 22244 13456
rect 24860 13447 24912 13456
rect 20628 13379 20680 13388
rect 20628 13345 20637 13379
rect 20637 13345 20671 13379
rect 20671 13345 20680 13379
rect 20628 13336 20680 13345
rect 22928 13379 22980 13388
rect 22928 13345 22937 13379
rect 22937 13345 22971 13379
rect 22971 13345 22980 13379
rect 22928 13336 22980 13345
rect 23848 13336 23900 13388
rect 24860 13413 24894 13447
rect 24894 13413 24912 13447
rect 24860 13404 24912 13413
rect 24676 13336 24728 13388
rect 27068 13379 27120 13388
rect 27068 13345 27077 13379
rect 27077 13345 27111 13379
rect 27111 13345 27120 13379
rect 27068 13336 27120 13345
rect 21180 13268 21232 13320
rect 15108 13132 15160 13184
rect 20996 13200 21048 13252
rect 18144 13132 18196 13184
rect 18696 13132 18748 13184
rect 19984 13132 20036 13184
rect 22468 13132 22520 13184
rect 24952 13132 25004 13184
rect 3756 13030 3808 13082
rect 3820 13030 3872 13082
rect 3884 13030 3936 13082
rect 3948 13030 4000 13082
rect 4012 13030 4064 13082
rect 10472 13030 10524 13082
rect 10536 13030 10588 13082
rect 10600 13030 10652 13082
rect 10664 13030 10716 13082
rect 10728 13030 10780 13082
rect 17188 13030 17240 13082
rect 17252 13030 17304 13082
rect 17316 13030 17368 13082
rect 17380 13030 17432 13082
rect 17444 13030 17496 13082
rect 23904 13030 23956 13082
rect 23968 13030 24020 13082
rect 24032 13030 24084 13082
rect 24096 13030 24148 13082
rect 24160 13030 24212 13082
rect 4160 12928 4212 12980
rect 7472 12928 7524 12980
rect 9404 12928 9456 12980
rect 14188 12928 14240 12980
rect 3792 12792 3844 12844
rect 4252 12792 4304 12844
rect 4620 12835 4672 12844
rect 4620 12801 4629 12835
rect 4629 12801 4663 12835
rect 4663 12801 4672 12835
rect 4620 12792 4672 12801
rect 6736 12860 6788 12912
rect 7012 12792 7064 12844
rect 12440 12860 12492 12912
rect 12532 12860 12584 12912
rect 15292 12928 15344 12980
rect 16304 12928 16356 12980
rect 18236 12928 18288 12980
rect 18604 12928 18656 12980
rect 20352 12928 20404 12980
rect 23020 12928 23072 12980
rect 25044 12928 25096 12980
rect 17868 12860 17920 12912
rect 19248 12860 19300 12912
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 3056 12767 3108 12776
rect 3056 12733 3065 12767
rect 3065 12733 3099 12767
rect 3099 12733 3108 12767
rect 3056 12724 3108 12733
rect 3148 12724 3200 12776
rect 4804 12767 4856 12776
rect 4804 12733 4813 12767
rect 4813 12733 4847 12767
rect 4847 12733 4856 12767
rect 4804 12724 4856 12733
rect 6552 12767 6604 12776
rect 6552 12733 6561 12767
rect 6561 12733 6595 12767
rect 6595 12733 6604 12767
rect 6552 12724 6604 12733
rect 7472 12767 7524 12776
rect 7472 12733 7481 12767
rect 7481 12733 7515 12767
rect 7515 12733 7524 12767
rect 7472 12724 7524 12733
rect 7564 12767 7616 12776
rect 7564 12733 7573 12767
rect 7573 12733 7607 12767
rect 7607 12733 7616 12767
rect 7564 12724 7616 12733
rect 8208 12724 8260 12776
rect 8668 12767 8720 12776
rect 8668 12733 8677 12767
rect 8677 12733 8711 12767
rect 8711 12733 8720 12767
rect 8668 12724 8720 12733
rect 8760 12767 8812 12776
rect 8760 12733 8769 12767
rect 8769 12733 8803 12767
rect 8803 12733 8812 12767
rect 8760 12724 8812 12733
rect 9496 12767 9548 12776
rect 9496 12733 9505 12767
rect 9505 12733 9539 12767
rect 9539 12733 9548 12767
rect 9496 12724 9548 12733
rect 9864 12724 9916 12776
rect 10140 12767 10192 12776
rect 10140 12733 10147 12767
rect 10147 12733 10192 12767
rect 10140 12724 10192 12733
rect 10232 12767 10284 12776
rect 10232 12733 10241 12767
rect 10241 12733 10275 12767
rect 10275 12733 10284 12767
rect 10232 12724 10284 12733
rect 10324 12767 10376 12776
rect 10324 12733 10333 12767
rect 10333 12733 10367 12767
rect 10367 12733 10376 12767
rect 10324 12724 10376 12733
rect 4068 12656 4120 12708
rect 4896 12656 4948 12708
rect 3332 12631 3384 12640
rect 3332 12597 3341 12631
rect 3341 12597 3375 12631
rect 3375 12597 3384 12631
rect 3332 12588 3384 12597
rect 3424 12588 3476 12640
rect 7472 12588 7524 12640
rect 9220 12656 9272 12708
rect 10692 12767 10744 12776
rect 10692 12733 10701 12767
rect 10701 12733 10735 12767
rect 10735 12733 10744 12767
rect 10692 12724 10744 12733
rect 10968 12656 11020 12708
rect 7932 12588 7984 12640
rect 8852 12588 8904 12640
rect 8944 12631 8996 12640
rect 8944 12597 8953 12631
rect 8953 12597 8987 12631
rect 8987 12597 8996 12631
rect 8944 12588 8996 12597
rect 9036 12588 9088 12640
rect 11612 12767 11664 12776
rect 11612 12733 11621 12767
rect 11621 12733 11655 12767
rect 11655 12733 11664 12767
rect 11612 12724 11664 12733
rect 15200 12835 15252 12844
rect 15200 12801 15209 12835
rect 15209 12801 15243 12835
rect 15243 12801 15252 12835
rect 15200 12792 15252 12801
rect 11796 12767 11848 12776
rect 11796 12733 11805 12767
rect 11805 12733 11839 12767
rect 11839 12733 11848 12767
rect 11796 12724 11848 12733
rect 11980 12724 12032 12776
rect 13268 12767 13320 12776
rect 12532 12656 12584 12708
rect 11336 12631 11388 12640
rect 11336 12597 11345 12631
rect 11345 12597 11379 12631
rect 11379 12597 11388 12631
rect 11336 12588 11388 12597
rect 12072 12631 12124 12640
rect 12072 12597 12081 12631
rect 12081 12597 12115 12631
rect 12115 12597 12124 12631
rect 12072 12588 12124 12597
rect 12256 12588 12308 12640
rect 13268 12733 13276 12767
rect 13276 12733 13310 12767
rect 13310 12733 13320 12767
rect 13268 12724 13320 12733
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 15108 12724 15160 12776
rect 15292 12767 15344 12776
rect 15292 12733 15301 12767
rect 15301 12733 15335 12767
rect 15335 12733 15344 12767
rect 15292 12724 15344 12733
rect 12992 12699 13044 12708
rect 12992 12665 13001 12699
rect 13001 12665 13035 12699
rect 13035 12665 13044 12699
rect 12992 12656 13044 12665
rect 13176 12656 13228 12708
rect 13452 12588 13504 12640
rect 14280 12656 14332 12708
rect 16672 12792 16724 12844
rect 15476 12767 15528 12776
rect 15476 12733 15485 12767
rect 15485 12733 15519 12767
rect 15519 12733 15528 12767
rect 15476 12724 15528 12733
rect 16488 12724 16540 12776
rect 16948 12767 17000 12776
rect 16948 12733 16957 12767
rect 16957 12733 16991 12767
rect 16991 12733 17000 12767
rect 16948 12724 17000 12733
rect 18328 12767 18380 12776
rect 18328 12733 18337 12767
rect 18337 12733 18371 12767
rect 18371 12733 18380 12767
rect 18328 12724 18380 12733
rect 22100 12767 22152 12776
rect 22100 12733 22109 12767
rect 22109 12733 22143 12767
rect 22143 12733 22152 12767
rect 22100 12724 22152 12733
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 23664 12792 23716 12844
rect 24860 12860 24912 12912
rect 23020 12724 23072 12776
rect 23388 12724 23440 12776
rect 15752 12656 15804 12708
rect 16672 12656 16724 12708
rect 14832 12588 14884 12640
rect 18236 12656 18288 12708
rect 20260 12656 20312 12708
rect 20444 12699 20496 12708
rect 20444 12665 20453 12699
rect 20453 12665 20487 12699
rect 20487 12665 20496 12699
rect 20444 12656 20496 12665
rect 24308 12767 24360 12776
rect 24308 12733 24322 12767
rect 24322 12733 24356 12767
rect 24356 12733 24360 12767
rect 24308 12724 24360 12733
rect 24492 12724 24544 12776
rect 24676 12724 24728 12776
rect 24860 12767 24912 12776
rect 24860 12733 24869 12767
rect 24869 12733 24903 12767
rect 24903 12733 24912 12767
rect 24860 12724 24912 12733
rect 24952 12767 25004 12776
rect 24952 12733 24961 12767
rect 24961 12733 24995 12767
rect 24995 12733 25004 12767
rect 24952 12724 25004 12733
rect 25320 12767 25372 12776
rect 25320 12733 25329 12767
rect 25329 12733 25363 12767
rect 25363 12733 25372 12767
rect 25320 12724 25372 12733
rect 25872 12860 25924 12912
rect 25688 12767 25740 12776
rect 25688 12733 25697 12767
rect 25697 12733 25731 12767
rect 25731 12733 25740 12767
rect 25688 12724 25740 12733
rect 25780 12724 25832 12776
rect 26424 12792 26476 12844
rect 17684 12631 17736 12640
rect 17684 12597 17693 12631
rect 17693 12597 17727 12631
rect 17727 12597 17736 12631
rect 17684 12588 17736 12597
rect 21180 12588 21232 12640
rect 21824 12588 21876 12640
rect 21916 12588 21968 12640
rect 26332 12699 26384 12708
rect 26332 12665 26341 12699
rect 26341 12665 26375 12699
rect 26375 12665 26384 12699
rect 26332 12656 26384 12665
rect 26424 12699 26476 12708
rect 26424 12665 26433 12699
rect 26433 12665 26467 12699
rect 26467 12665 26476 12699
rect 26424 12656 26476 12665
rect 24400 12588 24452 12640
rect 25228 12631 25280 12640
rect 25228 12597 25237 12631
rect 25237 12597 25271 12631
rect 25271 12597 25280 12631
rect 25228 12588 25280 12597
rect 7114 12486 7166 12538
rect 7178 12486 7230 12538
rect 7242 12486 7294 12538
rect 7306 12486 7358 12538
rect 7370 12486 7422 12538
rect 13830 12486 13882 12538
rect 13894 12486 13946 12538
rect 13958 12486 14010 12538
rect 14022 12486 14074 12538
rect 14086 12486 14138 12538
rect 20546 12486 20598 12538
rect 20610 12486 20662 12538
rect 20674 12486 20726 12538
rect 20738 12486 20790 12538
rect 20802 12486 20854 12538
rect 27262 12486 27314 12538
rect 27326 12486 27378 12538
rect 27390 12486 27442 12538
rect 27454 12486 27506 12538
rect 27518 12486 27570 12538
rect 2688 12384 2740 12436
rect 4804 12384 4856 12436
rect 6920 12384 6972 12436
rect 7748 12384 7800 12436
rect 8024 12384 8076 12436
rect 10876 12384 10928 12436
rect 14740 12384 14792 12436
rect 14924 12384 14976 12436
rect 16488 12384 16540 12436
rect 18328 12384 18380 12436
rect 27068 12384 27120 12436
rect 1400 12316 1452 12368
rect 3608 12316 3660 12368
rect 4160 12316 4212 12368
rect 4344 12316 4396 12368
rect 5172 12316 5224 12368
rect 8852 12316 8904 12368
rect 2044 12291 2096 12300
rect 2044 12257 2078 12291
rect 2078 12257 2096 12291
rect 2044 12248 2096 12257
rect 3332 12248 3384 12300
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 3792 12180 3844 12232
rect 3148 12087 3200 12096
rect 3148 12053 3157 12087
rect 3157 12053 3191 12087
rect 3191 12053 3200 12087
rect 3148 12044 3200 12053
rect 3608 12044 3660 12096
rect 4528 12291 4580 12300
rect 4528 12257 4537 12291
rect 4537 12257 4571 12291
rect 4571 12257 4580 12291
rect 4528 12248 4580 12257
rect 4804 12248 4856 12300
rect 6644 12291 6696 12300
rect 6644 12257 6653 12291
rect 6653 12257 6687 12291
rect 6687 12257 6696 12291
rect 6644 12248 6696 12257
rect 8576 12248 8628 12300
rect 8944 12291 8996 12300
rect 8944 12257 8953 12291
rect 8953 12257 8987 12291
rect 8987 12257 8996 12291
rect 8944 12248 8996 12257
rect 9036 12291 9088 12300
rect 9036 12257 9045 12291
rect 9045 12257 9079 12291
rect 9079 12257 9088 12291
rect 9036 12248 9088 12257
rect 9220 12291 9272 12300
rect 9220 12257 9229 12291
rect 9229 12257 9263 12291
rect 9263 12257 9272 12291
rect 9220 12248 9272 12257
rect 9496 12248 9548 12300
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 9864 12291 9916 12300
rect 9864 12257 9873 12291
rect 9873 12257 9907 12291
rect 9907 12257 9916 12291
rect 9864 12248 9916 12257
rect 11612 12316 11664 12368
rect 12808 12316 12860 12368
rect 14188 12316 14240 12368
rect 5448 12180 5500 12232
rect 4068 12155 4120 12164
rect 4068 12121 4077 12155
rect 4077 12121 4111 12155
rect 4111 12121 4120 12155
rect 4068 12112 4120 12121
rect 4436 12112 4488 12164
rect 4804 12112 4856 12164
rect 5356 12112 5408 12164
rect 9956 12180 10008 12232
rect 10232 12180 10284 12232
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 10968 12291 11020 12300
rect 10968 12257 10977 12291
rect 10977 12257 11011 12291
rect 11011 12257 11020 12291
rect 10968 12248 11020 12257
rect 11060 12248 11112 12300
rect 11244 12180 11296 12232
rect 11796 12180 11848 12232
rect 13084 12180 13136 12232
rect 5632 12044 5684 12096
rect 6644 12044 6696 12096
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 8576 12044 8628 12096
rect 9036 12044 9088 12096
rect 9404 12087 9456 12096
rect 9404 12053 9413 12087
rect 9413 12053 9447 12087
rect 9447 12053 9456 12087
rect 9404 12044 9456 12053
rect 12716 12112 12768 12164
rect 12808 12112 12860 12164
rect 13728 12044 13780 12096
rect 13820 12087 13872 12096
rect 13820 12053 13829 12087
rect 13829 12053 13863 12087
rect 13863 12053 13872 12087
rect 13820 12044 13872 12053
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 14832 12248 14884 12300
rect 15108 12294 15160 12300
rect 15108 12260 15117 12294
rect 15117 12260 15151 12294
rect 15151 12260 15160 12294
rect 15108 12248 15160 12260
rect 16764 12316 16816 12368
rect 16672 12291 16724 12300
rect 16672 12257 16681 12291
rect 16681 12257 16715 12291
rect 16715 12257 16724 12291
rect 16672 12248 16724 12257
rect 16304 12180 16356 12232
rect 17592 12291 17644 12300
rect 17592 12257 17601 12291
rect 17601 12257 17635 12291
rect 17635 12257 17644 12291
rect 17592 12248 17644 12257
rect 16948 12180 17000 12232
rect 17868 12291 17920 12300
rect 17868 12257 17877 12291
rect 17877 12257 17911 12291
rect 17911 12257 17920 12291
rect 17868 12248 17920 12257
rect 17960 12291 18012 12300
rect 17960 12257 17969 12291
rect 17969 12257 18003 12291
rect 18003 12257 18012 12291
rect 17960 12248 18012 12257
rect 18144 12248 18196 12300
rect 18420 12316 18472 12368
rect 18604 12291 18656 12300
rect 18604 12257 18613 12291
rect 18613 12257 18647 12291
rect 18647 12257 18656 12291
rect 18604 12248 18656 12257
rect 19800 12316 19852 12368
rect 25228 12316 25280 12368
rect 19524 12291 19576 12300
rect 19524 12257 19558 12291
rect 19558 12257 19576 12291
rect 19524 12248 19576 12257
rect 20444 12248 20496 12300
rect 26240 12248 26292 12300
rect 26884 12248 26936 12300
rect 19248 12223 19300 12232
rect 19248 12189 19257 12223
rect 19257 12189 19291 12223
rect 19291 12189 19300 12223
rect 19248 12180 19300 12189
rect 16120 12087 16172 12096
rect 16120 12053 16129 12087
rect 16129 12053 16163 12087
rect 16163 12053 16172 12087
rect 16120 12044 16172 12053
rect 21916 12180 21968 12232
rect 23756 12223 23808 12232
rect 23756 12189 23765 12223
rect 23765 12189 23799 12223
rect 23799 12189 23808 12223
rect 23756 12180 23808 12189
rect 24400 12223 24452 12232
rect 24400 12189 24409 12223
rect 24409 12189 24443 12223
rect 24443 12189 24452 12223
rect 24400 12180 24452 12189
rect 24768 12180 24820 12232
rect 26424 12223 26476 12232
rect 26424 12189 26433 12223
rect 26433 12189 26467 12223
rect 26467 12189 26476 12223
rect 26424 12180 26476 12189
rect 23020 12044 23072 12096
rect 23480 12044 23532 12096
rect 3756 11942 3808 11994
rect 3820 11942 3872 11994
rect 3884 11942 3936 11994
rect 3948 11942 4000 11994
rect 4012 11942 4064 11994
rect 10472 11942 10524 11994
rect 10536 11942 10588 11994
rect 10600 11942 10652 11994
rect 10664 11942 10716 11994
rect 10728 11942 10780 11994
rect 17188 11942 17240 11994
rect 17252 11942 17304 11994
rect 17316 11942 17368 11994
rect 17380 11942 17432 11994
rect 17444 11942 17496 11994
rect 23904 11942 23956 11994
rect 23968 11942 24020 11994
rect 24032 11942 24084 11994
rect 24096 11942 24148 11994
rect 24160 11942 24212 11994
rect 3608 11840 3660 11892
rect 4896 11840 4948 11892
rect 5908 11840 5960 11892
rect 9956 11840 10008 11892
rect 10232 11840 10284 11892
rect 9588 11772 9640 11824
rect 13176 11840 13228 11892
rect 13452 11840 13504 11892
rect 13728 11840 13780 11892
rect 12716 11772 12768 11824
rect 14556 11840 14608 11892
rect 16396 11840 16448 11892
rect 16948 11840 17000 11892
rect 18420 11840 18472 11892
rect 20352 11840 20404 11892
rect 21088 11840 21140 11892
rect 24400 11840 24452 11892
rect 26424 11883 26476 11892
rect 26424 11849 26433 11883
rect 26433 11849 26467 11883
rect 26467 11849 26476 11883
rect 26424 11840 26476 11849
rect 4804 11704 4856 11756
rect 3056 11636 3108 11688
rect 4712 11679 4764 11688
rect 4712 11645 4721 11679
rect 4721 11645 4755 11679
rect 4755 11645 4764 11679
rect 4712 11636 4764 11645
rect 5356 11636 5408 11688
rect 6000 11636 6052 11688
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 7012 11704 7064 11756
rect 9128 11636 9180 11688
rect 9312 11636 9364 11688
rect 8392 11568 8444 11620
rect 8484 11568 8536 11620
rect 9864 11568 9916 11620
rect 10140 11568 10192 11620
rect 10968 11568 11020 11620
rect 11060 11568 11112 11620
rect 11612 11568 11664 11620
rect 12072 11568 12124 11620
rect 13820 11679 13872 11688
rect 13820 11645 13854 11679
rect 13854 11645 13872 11679
rect 13176 11568 13228 11620
rect 13820 11636 13872 11645
rect 15200 11679 15252 11688
rect 15200 11645 15209 11679
rect 15209 11645 15243 11679
rect 15243 11645 15252 11679
rect 15200 11636 15252 11645
rect 17684 11636 17736 11688
rect 21272 11747 21324 11756
rect 21272 11713 21281 11747
rect 21281 11713 21315 11747
rect 21315 11713 21324 11747
rect 21272 11704 21324 11713
rect 23756 11704 23808 11756
rect 24768 11704 24820 11756
rect 24400 11679 24452 11688
rect 24400 11645 24409 11679
rect 24409 11645 24443 11679
rect 24443 11645 24452 11679
rect 24400 11636 24452 11645
rect 16120 11568 16172 11620
rect 16488 11568 16540 11620
rect 18052 11568 18104 11620
rect 21640 11568 21692 11620
rect 25596 11568 25648 11620
rect 9036 11500 9088 11552
rect 9588 11500 9640 11552
rect 10324 11500 10376 11552
rect 16028 11500 16080 11552
rect 7114 11398 7166 11450
rect 7178 11398 7230 11450
rect 7242 11398 7294 11450
rect 7306 11398 7358 11450
rect 7370 11398 7422 11450
rect 13830 11398 13882 11450
rect 13894 11398 13946 11450
rect 13958 11398 14010 11450
rect 14022 11398 14074 11450
rect 14086 11398 14138 11450
rect 20546 11398 20598 11450
rect 20610 11398 20662 11450
rect 20674 11398 20726 11450
rect 20738 11398 20790 11450
rect 20802 11398 20854 11450
rect 27262 11398 27314 11450
rect 27326 11398 27378 11450
rect 27390 11398 27442 11450
rect 27454 11398 27506 11450
rect 27518 11398 27570 11450
rect 4436 11296 4488 11348
rect 4988 11296 5040 11348
rect 8392 11296 8444 11348
rect 10232 11296 10284 11348
rect 2688 11160 2740 11212
rect 4436 11203 4488 11212
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 4988 11203 5040 11212
rect 4988 11169 4997 11203
rect 4997 11169 5031 11203
rect 5031 11169 5040 11203
rect 4988 11160 5040 11169
rect 5172 11203 5224 11212
rect 5172 11169 5181 11203
rect 5181 11169 5215 11203
rect 5215 11169 5224 11203
rect 5172 11160 5224 11169
rect 5356 11160 5408 11212
rect 5540 11160 5592 11212
rect 5724 11160 5776 11212
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 10048 11228 10100 11280
rect 11612 11339 11664 11348
rect 11612 11305 11621 11339
rect 11621 11305 11655 11339
rect 11655 11305 11664 11339
rect 11612 11296 11664 11305
rect 10876 11228 10928 11280
rect 12624 11296 12676 11348
rect 13084 11339 13136 11348
rect 13084 11305 13093 11339
rect 13093 11305 13127 11339
rect 13127 11305 13136 11339
rect 13084 11296 13136 11305
rect 13452 11296 13504 11348
rect 14832 11296 14884 11348
rect 15476 11296 15528 11348
rect 17960 11296 18012 11348
rect 6920 11203 6972 11212
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 7564 11160 7616 11212
rect 8300 11160 8352 11212
rect 8668 11160 8720 11212
rect 9772 11160 9824 11212
rect 12256 11228 12308 11280
rect 5172 10956 5224 11008
rect 5540 10999 5592 11008
rect 5540 10965 5549 10999
rect 5549 10965 5583 10999
rect 5583 10965 5592 10999
rect 5540 10956 5592 10965
rect 7656 10956 7708 11008
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 12440 11203 12492 11212
rect 12440 11169 12449 11203
rect 12449 11169 12483 11203
rect 12483 11169 12492 11203
rect 12440 11160 12492 11169
rect 17868 11228 17920 11280
rect 12808 11203 12860 11212
rect 12808 11169 12817 11203
rect 12817 11169 12851 11203
rect 12851 11169 12860 11203
rect 12808 11160 12860 11169
rect 13176 11203 13228 11212
rect 13176 11169 13185 11203
rect 13185 11169 13219 11203
rect 13219 11169 13228 11203
rect 13176 11160 13228 11169
rect 13452 11203 13504 11212
rect 13452 11169 13486 11203
rect 13486 11169 13504 11203
rect 13452 11160 13504 11169
rect 12716 11024 12768 11076
rect 13084 11024 13136 11076
rect 13176 11024 13228 11076
rect 14556 11092 14608 11144
rect 14832 11160 14884 11212
rect 15108 11203 15160 11212
rect 15108 11169 15122 11203
rect 15122 11169 15156 11203
rect 15156 11169 15160 11203
rect 15108 11160 15160 11169
rect 15476 11160 15528 11212
rect 15752 11160 15804 11212
rect 18604 11160 18656 11212
rect 19248 11160 19300 11212
rect 19524 11339 19576 11348
rect 19524 11305 19533 11339
rect 19533 11305 19567 11339
rect 19567 11305 19576 11339
rect 19524 11296 19576 11305
rect 19800 11203 19852 11212
rect 19800 11169 19809 11203
rect 19809 11169 19843 11203
rect 19843 11169 19852 11203
rect 19800 11160 19852 11169
rect 18788 11092 18840 11144
rect 19984 11203 20036 11212
rect 19984 11169 19993 11203
rect 19993 11169 20027 11203
rect 20027 11169 20036 11203
rect 19984 11160 20036 11169
rect 20996 11296 21048 11348
rect 22652 11339 22704 11348
rect 22652 11305 22661 11339
rect 22661 11305 22695 11339
rect 22695 11305 22704 11339
rect 22652 11296 22704 11305
rect 26240 11296 26292 11348
rect 22192 11228 22244 11280
rect 20536 11203 20588 11212
rect 20536 11169 20545 11203
rect 20545 11169 20579 11203
rect 20579 11169 20588 11203
rect 20536 11160 20588 11169
rect 21088 11160 21140 11212
rect 21272 11203 21324 11212
rect 21272 11169 21281 11203
rect 21281 11169 21315 11203
rect 21315 11169 21324 11203
rect 21272 11160 21324 11169
rect 21548 11203 21600 11212
rect 21548 11169 21582 11203
rect 21582 11169 21600 11203
rect 21548 11160 21600 11169
rect 24952 11160 25004 11212
rect 26240 11203 26292 11212
rect 26240 11169 26249 11203
rect 26249 11169 26283 11203
rect 26283 11169 26292 11203
rect 26240 11160 26292 11169
rect 12164 10956 12216 11008
rect 13360 10956 13412 11008
rect 17592 11024 17644 11076
rect 20812 11092 20864 11144
rect 23756 11092 23808 11144
rect 25320 11092 25372 11144
rect 20352 11024 20404 11076
rect 20536 11024 20588 11076
rect 25136 11024 25188 11076
rect 26884 11160 26936 11212
rect 18052 10956 18104 11008
rect 20168 10956 20220 11008
rect 22376 10956 22428 11008
rect 24492 10956 24544 11008
rect 24768 10956 24820 11008
rect 25780 10956 25832 11008
rect 27068 10999 27120 11008
rect 27068 10965 27077 10999
rect 27077 10965 27111 10999
rect 27111 10965 27120 10999
rect 27068 10956 27120 10965
rect 3756 10854 3808 10906
rect 3820 10854 3872 10906
rect 3884 10854 3936 10906
rect 3948 10854 4000 10906
rect 4012 10854 4064 10906
rect 10472 10854 10524 10906
rect 10536 10854 10588 10906
rect 10600 10854 10652 10906
rect 10664 10854 10716 10906
rect 10728 10854 10780 10906
rect 17188 10854 17240 10906
rect 17252 10854 17304 10906
rect 17316 10854 17368 10906
rect 17380 10854 17432 10906
rect 17444 10854 17496 10906
rect 23904 10854 23956 10906
rect 23968 10854 24020 10906
rect 24032 10854 24084 10906
rect 24096 10854 24148 10906
rect 24160 10854 24212 10906
rect 7840 10752 7892 10804
rect 4988 10616 5040 10668
rect 3148 10548 3200 10600
rect 4160 10480 4212 10532
rect 4344 10412 4396 10464
rect 4620 10591 4672 10600
rect 4620 10557 4629 10591
rect 4629 10557 4663 10591
rect 4663 10557 4672 10591
rect 4620 10548 4672 10557
rect 6000 10591 6052 10600
rect 6000 10557 6009 10591
rect 6009 10557 6043 10591
rect 6043 10557 6052 10591
rect 6000 10548 6052 10557
rect 8024 10684 8076 10736
rect 6828 10548 6880 10600
rect 7012 10548 7064 10600
rect 7472 10616 7524 10668
rect 8300 10548 8352 10600
rect 4804 10480 4856 10532
rect 5080 10523 5132 10532
rect 5080 10489 5089 10523
rect 5089 10489 5123 10523
rect 5123 10489 5132 10523
rect 5080 10480 5132 10489
rect 10048 10727 10100 10736
rect 10048 10693 10057 10727
rect 10057 10693 10091 10727
rect 10091 10693 10100 10727
rect 10048 10684 10100 10693
rect 16580 10795 16632 10804
rect 16580 10761 16589 10795
rect 16589 10761 16623 10795
rect 16623 10761 16632 10795
rect 16580 10752 16632 10761
rect 18144 10752 18196 10804
rect 18604 10752 18656 10804
rect 20812 10795 20864 10804
rect 20812 10761 20821 10795
rect 20821 10761 20855 10795
rect 20855 10761 20864 10795
rect 20812 10752 20864 10761
rect 21548 10795 21600 10804
rect 21548 10761 21557 10795
rect 21557 10761 21591 10795
rect 21591 10761 21600 10795
rect 21548 10752 21600 10761
rect 21640 10795 21692 10804
rect 21640 10761 21649 10795
rect 21649 10761 21683 10795
rect 21683 10761 21692 10795
rect 21640 10752 21692 10761
rect 24400 10752 24452 10804
rect 24952 10752 25004 10804
rect 8576 10616 8628 10668
rect 9404 10616 9456 10668
rect 8668 10548 8720 10600
rect 8760 10548 8812 10600
rect 10324 10659 10376 10668
rect 10324 10625 10333 10659
rect 10333 10625 10367 10659
rect 10367 10625 10376 10659
rect 10324 10616 10376 10625
rect 11060 10616 11112 10668
rect 12992 10616 13044 10668
rect 14740 10659 14792 10668
rect 14740 10625 14749 10659
rect 14749 10625 14783 10659
rect 14783 10625 14792 10659
rect 14740 10616 14792 10625
rect 14832 10616 14884 10668
rect 20168 10684 20220 10736
rect 9588 10548 9640 10600
rect 11244 10548 11296 10600
rect 15660 10548 15712 10600
rect 5356 10455 5408 10464
rect 5356 10421 5365 10455
rect 5365 10421 5399 10455
rect 5399 10421 5408 10455
rect 5356 10412 5408 10421
rect 5448 10412 5500 10464
rect 7564 10455 7616 10464
rect 7564 10421 7573 10455
rect 7573 10421 7607 10455
rect 7607 10421 7616 10455
rect 7564 10412 7616 10421
rect 8300 10412 8352 10464
rect 11980 10480 12032 10532
rect 12256 10480 12308 10532
rect 17868 10591 17920 10600
rect 17868 10557 17877 10591
rect 17877 10557 17911 10591
rect 17911 10557 17920 10591
rect 17868 10548 17920 10557
rect 18236 10616 18288 10668
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 18144 10548 18196 10600
rect 19984 10616 20036 10668
rect 20536 10616 20588 10668
rect 20168 10548 20220 10600
rect 20352 10591 20404 10600
rect 20352 10557 20361 10591
rect 20361 10557 20395 10591
rect 20395 10557 20404 10591
rect 20352 10548 20404 10557
rect 9220 10412 9272 10464
rect 9772 10412 9824 10464
rect 13728 10412 13780 10464
rect 15384 10412 15436 10464
rect 17592 10480 17644 10532
rect 19064 10480 19116 10532
rect 20996 10548 21048 10600
rect 21088 10591 21140 10600
rect 21088 10557 21097 10591
rect 21097 10557 21131 10591
rect 21131 10557 21140 10591
rect 21088 10548 21140 10557
rect 22100 10616 22152 10668
rect 22192 10659 22244 10668
rect 22192 10625 22201 10659
rect 22201 10625 22235 10659
rect 22235 10625 22244 10659
rect 22192 10616 22244 10625
rect 22376 10548 22428 10600
rect 22928 10591 22980 10600
rect 22928 10557 22937 10591
rect 22937 10557 22971 10591
rect 22971 10557 22980 10591
rect 22928 10548 22980 10557
rect 22836 10480 22888 10532
rect 23480 10548 23532 10600
rect 24768 10616 24820 10668
rect 26792 10659 26844 10668
rect 26792 10625 26801 10659
rect 26801 10625 26835 10659
rect 26835 10625 26844 10659
rect 26792 10616 26844 10625
rect 24492 10591 24544 10600
rect 24492 10557 24501 10591
rect 24501 10557 24535 10591
rect 24535 10557 24544 10591
rect 24492 10548 24544 10557
rect 25136 10548 25188 10600
rect 17684 10412 17736 10464
rect 18880 10412 18932 10464
rect 19800 10412 19852 10464
rect 20260 10412 20312 10464
rect 22100 10412 22152 10464
rect 24860 10480 24912 10532
rect 25780 10480 25832 10532
rect 25136 10412 25188 10464
rect 25228 10412 25280 10464
rect 7114 10310 7166 10362
rect 7178 10310 7230 10362
rect 7242 10310 7294 10362
rect 7306 10310 7358 10362
rect 7370 10310 7422 10362
rect 13830 10310 13882 10362
rect 13894 10310 13946 10362
rect 13958 10310 14010 10362
rect 14022 10310 14074 10362
rect 14086 10310 14138 10362
rect 20546 10310 20598 10362
rect 20610 10310 20662 10362
rect 20674 10310 20726 10362
rect 20738 10310 20790 10362
rect 20802 10310 20854 10362
rect 27262 10310 27314 10362
rect 27326 10310 27378 10362
rect 27390 10310 27442 10362
rect 27454 10310 27506 10362
rect 27518 10310 27570 10362
rect 4620 10208 4672 10260
rect 5264 10208 5316 10260
rect 5448 10208 5500 10260
rect 8668 10251 8720 10260
rect 8668 10217 8677 10251
rect 8677 10217 8711 10251
rect 8711 10217 8720 10251
rect 8668 10208 8720 10217
rect 11980 10251 12032 10260
rect 11980 10217 11989 10251
rect 11989 10217 12023 10251
rect 12023 10217 12032 10251
rect 11980 10208 12032 10217
rect 12532 10208 12584 10260
rect 2688 10072 2740 10124
rect 2872 10115 2924 10124
rect 2872 10081 2906 10115
rect 2906 10081 2924 10115
rect 2872 10072 2924 10081
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 4988 10072 5040 10124
rect 5264 10115 5316 10124
rect 5264 10081 5273 10115
rect 5273 10081 5307 10115
rect 5307 10081 5316 10115
rect 10324 10140 10376 10192
rect 11520 10140 11572 10192
rect 12164 10140 12216 10192
rect 13452 10208 13504 10260
rect 15200 10251 15252 10260
rect 15200 10217 15209 10251
rect 15209 10217 15243 10251
rect 15243 10217 15252 10251
rect 15200 10208 15252 10217
rect 5264 10072 5316 10081
rect 7564 10115 7616 10124
rect 7564 10081 7598 10115
rect 7598 10081 7616 10115
rect 7564 10072 7616 10081
rect 9128 10115 9180 10124
rect 9128 10081 9137 10115
rect 9137 10081 9171 10115
rect 9171 10081 9180 10115
rect 9128 10072 9180 10081
rect 9404 10115 9456 10124
rect 9404 10081 9438 10115
rect 9438 10081 9456 10115
rect 9404 10072 9456 10081
rect 12256 10115 12308 10124
rect 12256 10081 12265 10115
rect 12265 10081 12299 10115
rect 12299 10081 12308 10115
rect 12256 10072 12308 10081
rect 12532 10072 12584 10124
rect 12808 10072 12860 10124
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 4804 10004 4856 10056
rect 4252 9911 4304 9920
rect 4252 9877 4261 9911
rect 4261 9877 4295 9911
rect 4295 9877 4304 9911
rect 4252 9868 4304 9877
rect 4344 9868 4396 9920
rect 5816 9911 5868 9920
rect 5816 9877 5825 9911
rect 5825 9877 5859 9911
rect 5859 9877 5868 9911
rect 5816 9868 5868 9877
rect 6920 10004 6972 10056
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 11244 10004 11296 10013
rect 12164 9936 12216 9988
rect 13360 10115 13412 10124
rect 13360 10081 13369 10115
rect 13369 10081 13403 10115
rect 13403 10081 13412 10115
rect 13360 10072 13412 10081
rect 13452 10004 13504 10056
rect 13820 10115 13872 10124
rect 13820 10081 13843 10115
rect 13843 10081 13872 10115
rect 13820 10072 13872 10081
rect 16304 10140 16356 10192
rect 16672 10208 16724 10260
rect 17040 10208 17092 10260
rect 17684 10251 17736 10260
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 17684 10208 17736 10217
rect 17868 10208 17920 10260
rect 19064 10208 19116 10260
rect 14188 10115 14240 10124
rect 14188 10081 14197 10115
rect 14197 10081 14231 10115
rect 14231 10081 14240 10115
rect 14188 10072 14240 10081
rect 14832 10072 14884 10124
rect 15384 10115 15436 10124
rect 15384 10081 15393 10115
rect 15393 10081 15427 10115
rect 15427 10081 15436 10115
rect 15384 10072 15436 10081
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 15752 10115 15804 10124
rect 15752 10081 15761 10115
rect 15761 10081 15795 10115
rect 15795 10081 15804 10115
rect 15752 10072 15804 10081
rect 17040 10072 17092 10124
rect 18604 10115 18656 10124
rect 18604 10081 18613 10115
rect 18613 10081 18647 10115
rect 18647 10081 18656 10115
rect 18604 10072 18656 10081
rect 13360 9936 13412 9988
rect 14188 9936 14240 9988
rect 15016 10004 15068 10056
rect 16304 10004 16356 10056
rect 18236 10047 18288 10056
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 18880 10115 18932 10124
rect 18880 10081 18889 10115
rect 18889 10081 18923 10115
rect 18923 10081 18932 10115
rect 18880 10072 18932 10081
rect 19064 10072 19116 10124
rect 19340 10115 19392 10124
rect 19340 10081 19349 10115
rect 19349 10081 19383 10115
rect 19383 10081 19392 10115
rect 19340 10072 19392 10081
rect 20996 10208 21048 10260
rect 21088 10208 21140 10260
rect 21364 10140 21416 10192
rect 22284 10208 22336 10260
rect 22928 10208 22980 10260
rect 24400 10208 24452 10260
rect 24492 10208 24544 10260
rect 25596 10251 25648 10260
rect 25596 10217 25605 10251
rect 25605 10217 25639 10251
rect 25639 10217 25648 10251
rect 25596 10208 25648 10217
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 20168 10115 20220 10124
rect 20168 10081 20177 10115
rect 20177 10081 20211 10115
rect 20211 10081 20220 10115
rect 20168 10072 20220 10081
rect 20352 10072 20404 10124
rect 20812 10072 20864 10124
rect 21640 10115 21692 10124
rect 21640 10081 21649 10115
rect 21649 10081 21683 10115
rect 21683 10081 21692 10115
rect 21640 10072 21692 10081
rect 21732 10115 21784 10124
rect 21732 10081 21741 10115
rect 21741 10081 21775 10115
rect 21775 10081 21784 10115
rect 21732 10072 21784 10081
rect 22836 10072 22888 10124
rect 23664 10140 23716 10192
rect 25320 10140 25372 10192
rect 24308 10115 24360 10124
rect 24308 10081 24317 10115
rect 24317 10081 24351 10115
rect 24351 10081 24360 10115
rect 24308 10072 24360 10081
rect 24492 10072 24544 10124
rect 24768 10072 24820 10124
rect 25136 10115 25188 10124
rect 25136 10081 25145 10115
rect 25145 10081 25179 10115
rect 25179 10081 25188 10115
rect 25136 10072 25188 10081
rect 25228 10115 25280 10124
rect 25228 10081 25237 10115
rect 25237 10081 25271 10115
rect 25271 10081 25280 10115
rect 25228 10072 25280 10081
rect 27068 10072 27120 10124
rect 6920 9868 6972 9920
rect 10324 9868 10376 9920
rect 11980 9868 12032 9920
rect 12716 9911 12768 9920
rect 12716 9877 12725 9911
rect 12725 9877 12759 9911
rect 12759 9877 12768 9911
rect 12716 9868 12768 9877
rect 12808 9868 12860 9920
rect 16856 9911 16908 9920
rect 16856 9877 16865 9911
rect 16865 9877 16899 9911
rect 16899 9877 16908 9911
rect 16856 9868 16908 9877
rect 17684 9868 17736 9920
rect 17868 9868 17920 9920
rect 18880 9868 18932 9920
rect 21732 9936 21784 9988
rect 26884 10004 26936 10056
rect 24860 9936 24912 9988
rect 19616 9868 19668 9920
rect 19800 9868 19852 9920
rect 23480 9868 23532 9920
rect 24492 9868 24544 9920
rect 25136 9868 25188 9920
rect 25780 9868 25832 9920
rect 3756 9766 3808 9818
rect 3820 9766 3872 9818
rect 3884 9766 3936 9818
rect 3948 9766 4000 9818
rect 4012 9766 4064 9818
rect 10472 9766 10524 9818
rect 10536 9766 10588 9818
rect 10600 9766 10652 9818
rect 10664 9766 10716 9818
rect 10728 9766 10780 9818
rect 17188 9766 17240 9818
rect 17252 9766 17304 9818
rect 17316 9766 17368 9818
rect 17380 9766 17432 9818
rect 17444 9766 17496 9818
rect 23904 9766 23956 9818
rect 23968 9766 24020 9818
rect 24032 9766 24084 9818
rect 24096 9766 24148 9818
rect 24160 9766 24212 9818
rect 2872 9664 2924 9716
rect 7012 9664 7064 9716
rect 7564 9707 7616 9716
rect 7564 9673 7573 9707
rect 7573 9673 7607 9707
rect 7607 9673 7616 9707
rect 7564 9664 7616 9673
rect 9404 9664 9456 9716
rect 4160 9596 4212 9648
rect 5540 9596 5592 9648
rect 5724 9596 5776 9648
rect 11244 9664 11296 9716
rect 13176 9664 13228 9716
rect 15476 9664 15528 9716
rect 16304 9664 16356 9716
rect 13268 9596 13320 9648
rect 20444 9664 20496 9716
rect 23664 9664 23716 9716
rect 25228 9664 25280 9716
rect 26792 9664 26844 9716
rect 17592 9596 17644 9648
rect 17776 9596 17828 9648
rect 19432 9639 19484 9648
rect 19432 9605 19441 9639
rect 19441 9605 19475 9639
rect 19475 9605 19484 9639
rect 19432 9596 19484 9605
rect 20076 9596 20128 9648
rect 24676 9639 24728 9648
rect 24676 9605 24685 9639
rect 24685 9605 24719 9639
rect 24719 9605 24728 9639
rect 24676 9596 24728 9605
rect 3332 9503 3384 9512
rect 3332 9469 3341 9503
rect 3341 9469 3375 9503
rect 3375 9469 3384 9503
rect 3332 9460 3384 9469
rect 4252 9460 4304 9512
rect 5816 9528 5868 9580
rect 4804 9503 4856 9512
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 5356 9460 5408 9512
rect 6368 9503 6420 9512
rect 6368 9469 6377 9503
rect 6377 9469 6411 9503
rect 6411 9469 6420 9503
rect 6368 9460 6420 9469
rect 3240 9392 3292 9444
rect 4436 9392 4488 9444
rect 4988 9392 5040 9444
rect 6644 9503 6696 9512
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 6644 9460 6696 9469
rect 6552 9392 6604 9444
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 2964 9324 3016 9376
rect 6276 9324 6328 9376
rect 7012 9503 7064 9512
rect 7012 9469 7021 9503
rect 7021 9469 7055 9503
rect 7055 9469 7064 9503
rect 7012 9460 7064 9469
rect 7380 9528 7432 9580
rect 8300 9460 8352 9512
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 8760 9460 8812 9512
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 9680 9528 9732 9580
rect 14280 9571 14332 9580
rect 14280 9537 14289 9571
rect 14289 9537 14323 9571
rect 14323 9537 14332 9571
rect 14280 9528 14332 9537
rect 9312 9503 9364 9512
rect 9312 9469 9321 9503
rect 9321 9469 9355 9503
rect 9355 9469 9364 9503
rect 9312 9460 9364 9469
rect 10324 9460 10376 9512
rect 11060 9460 11112 9512
rect 13452 9460 13504 9512
rect 16856 9460 16908 9512
rect 17592 9460 17644 9512
rect 18236 9571 18288 9580
rect 18236 9537 18245 9571
rect 18245 9537 18279 9571
rect 18279 9537 18288 9571
rect 18236 9528 18288 9537
rect 7564 9324 7616 9376
rect 11152 9392 11204 9444
rect 12072 9392 12124 9444
rect 9404 9324 9456 9376
rect 15384 9392 15436 9444
rect 16028 9435 16080 9444
rect 16028 9401 16037 9435
rect 16037 9401 16071 9435
rect 16071 9401 16080 9435
rect 16028 9392 16080 9401
rect 12532 9324 12584 9376
rect 12808 9324 12860 9376
rect 17868 9392 17920 9444
rect 18972 9460 19024 9512
rect 16764 9324 16816 9376
rect 19064 9367 19116 9376
rect 19064 9333 19073 9367
rect 19073 9333 19107 9367
rect 19107 9333 19116 9367
rect 19064 9324 19116 9333
rect 20352 9324 20404 9376
rect 21364 9460 21416 9512
rect 23756 9528 23808 9580
rect 23848 9503 23900 9512
rect 20812 9324 20864 9376
rect 20904 9324 20956 9376
rect 21456 9367 21508 9376
rect 21456 9333 21465 9367
rect 21465 9333 21499 9367
rect 21499 9333 21508 9367
rect 21456 9324 21508 9333
rect 23848 9469 23857 9503
rect 23857 9469 23891 9503
rect 23891 9469 23900 9503
rect 23848 9460 23900 9469
rect 24860 9503 24912 9512
rect 24860 9469 24869 9503
rect 24869 9469 24903 9503
rect 24903 9469 24912 9503
rect 24860 9460 24912 9469
rect 21732 9392 21784 9444
rect 23204 9392 23256 9444
rect 22928 9324 22980 9376
rect 24124 9392 24176 9444
rect 24308 9392 24360 9444
rect 25412 9460 25464 9512
rect 25780 9503 25832 9512
rect 25780 9469 25814 9503
rect 25814 9469 25832 9503
rect 25780 9460 25832 9469
rect 23756 9324 23808 9376
rect 24584 9324 24636 9376
rect 7114 9222 7166 9274
rect 7178 9222 7230 9274
rect 7242 9222 7294 9274
rect 7306 9222 7358 9274
rect 7370 9222 7422 9274
rect 13830 9222 13882 9274
rect 13894 9222 13946 9274
rect 13958 9222 14010 9274
rect 14022 9222 14074 9274
rect 14086 9222 14138 9274
rect 20546 9222 20598 9274
rect 20610 9222 20662 9274
rect 20674 9222 20726 9274
rect 20738 9222 20790 9274
rect 20802 9222 20854 9274
rect 27262 9222 27314 9274
rect 27326 9222 27378 9274
rect 27390 9222 27442 9274
rect 27454 9222 27506 9274
rect 27518 9222 27570 9274
rect 7012 9120 7064 9172
rect 6368 9052 6420 9104
rect 3608 8984 3660 9036
rect 6920 9052 6972 9104
rect 1584 8916 1636 8968
rect 4896 8916 4948 8968
rect 6644 8984 6696 9036
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 7288 9027 7340 9036
rect 7288 8993 7297 9027
rect 7297 8993 7331 9027
rect 7331 8993 7340 9027
rect 7288 8984 7340 8993
rect 11152 9120 11204 9172
rect 12072 9163 12124 9172
rect 12072 9129 12081 9163
rect 12081 9129 12115 9163
rect 12115 9129 12124 9163
rect 12072 9120 12124 9129
rect 7564 9027 7616 9036
rect 7564 8993 7573 9027
rect 7573 8993 7607 9027
rect 7607 8993 7616 9027
rect 7564 8984 7616 8993
rect 8208 9027 8260 9036
rect 8208 8993 8217 9027
rect 8217 8993 8251 9027
rect 8251 8993 8260 9027
rect 8208 8984 8260 8993
rect 8300 9027 8352 9036
rect 8300 8993 8310 9027
rect 8310 8993 8344 9027
rect 8344 8993 8352 9027
rect 8300 8984 8352 8993
rect 8484 9027 8536 9036
rect 8484 8993 8493 9027
rect 8493 8993 8527 9027
rect 8527 8993 8536 9027
rect 8484 8984 8536 8993
rect 7656 8916 7708 8968
rect 8668 9027 8720 9036
rect 8668 8993 8682 9027
rect 8682 8993 8716 9027
rect 8716 8993 8720 9027
rect 8668 8984 8720 8993
rect 9128 9027 9180 9036
rect 9128 8993 9137 9027
rect 9137 8993 9171 9027
rect 9171 8993 9180 9027
rect 9128 8984 9180 8993
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 9496 9027 9548 9036
rect 9496 8993 9505 9027
rect 9505 8993 9539 9027
rect 9539 8993 9548 9027
rect 9496 8984 9548 8993
rect 12716 9120 12768 9172
rect 16764 9120 16816 9172
rect 18236 9120 18288 9172
rect 19064 9120 19116 9172
rect 12256 8984 12308 9036
rect 13268 9052 13320 9104
rect 12440 9027 12492 9036
rect 12440 8993 12449 9027
rect 12449 8993 12483 9027
rect 12483 8993 12492 9027
rect 12440 8984 12492 8993
rect 7564 8848 7616 8900
rect 8852 8891 8904 8900
rect 8852 8857 8861 8891
rect 8861 8857 8895 8891
rect 8895 8857 8904 8891
rect 8852 8848 8904 8857
rect 4436 8780 4488 8832
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 8208 8780 8260 8832
rect 8944 8780 8996 8832
rect 11336 8848 11388 8900
rect 12532 8848 12584 8900
rect 12808 8984 12860 9036
rect 14556 8984 14608 9036
rect 15660 9027 15712 9036
rect 15660 8993 15669 9027
rect 15669 8993 15703 9027
rect 15703 8993 15712 9027
rect 15660 8984 15712 8993
rect 15936 9027 15988 9036
rect 15936 8993 15945 9027
rect 15945 8993 15979 9027
rect 15979 8993 15988 9027
rect 15936 8984 15988 8993
rect 16580 9052 16632 9104
rect 17960 9052 18012 9104
rect 20904 9120 20956 9172
rect 21640 9120 21692 9172
rect 23204 9163 23256 9172
rect 23204 9129 23213 9163
rect 23213 9129 23247 9163
rect 23247 9129 23256 9163
rect 23204 9120 23256 9129
rect 23848 9120 23900 9172
rect 26884 9163 26936 9172
rect 26884 9129 26893 9163
rect 26893 9129 26927 9163
rect 26927 9129 26936 9163
rect 26884 9120 26936 9129
rect 20076 9052 20128 9104
rect 23480 9052 23532 9104
rect 18236 8984 18288 9036
rect 19524 8984 19576 9036
rect 15752 8848 15804 8900
rect 17132 8916 17184 8968
rect 17684 8916 17736 8968
rect 18052 8959 18104 8968
rect 18052 8925 18061 8959
rect 18061 8925 18095 8959
rect 18095 8925 18104 8959
rect 18052 8916 18104 8925
rect 18696 8916 18748 8968
rect 21456 8984 21508 9036
rect 19800 8916 19852 8968
rect 21640 8916 21692 8968
rect 23388 8984 23440 9036
rect 23664 9027 23716 9036
rect 23664 8993 23673 9027
rect 23673 8993 23707 9027
rect 23707 8993 23716 9027
rect 23664 8984 23716 8993
rect 24124 8984 24176 9036
rect 25320 9052 25372 9104
rect 25872 9052 25924 9104
rect 24952 8984 25004 9036
rect 25412 8984 25464 9036
rect 24308 8959 24360 8968
rect 24308 8925 24317 8959
rect 24317 8925 24351 8959
rect 24351 8925 24360 8959
rect 24308 8916 24360 8925
rect 24400 8959 24452 8968
rect 24400 8925 24409 8959
rect 24409 8925 24443 8959
rect 24443 8925 24452 8959
rect 24400 8916 24452 8925
rect 23480 8848 23532 8900
rect 24124 8848 24176 8900
rect 24768 8848 24820 8900
rect 17776 8780 17828 8832
rect 21272 8780 21324 8832
rect 22468 8780 22520 8832
rect 24860 8780 24912 8832
rect 3756 8678 3808 8730
rect 3820 8678 3872 8730
rect 3884 8678 3936 8730
rect 3948 8678 4000 8730
rect 4012 8678 4064 8730
rect 10472 8678 10524 8730
rect 10536 8678 10588 8730
rect 10600 8678 10652 8730
rect 10664 8678 10716 8730
rect 10728 8678 10780 8730
rect 17188 8678 17240 8730
rect 17252 8678 17304 8730
rect 17316 8678 17368 8730
rect 17380 8678 17432 8730
rect 17444 8678 17496 8730
rect 23904 8678 23956 8730
rect 23968 8678 24020 8730
rect 24032 8678 24084 8730
rect 24096 8678 24148 8730
rect 24160 8678 24212 8730
rect 3608 8576 3660 8628
rect 7656 8619 7708 8628
rect 7656 8585 7665 8619
rect 7665 8585 7699 8619
rect 7699 8585 7708 8619
rect 7656 8576 7708 8585
rect 8392 8576 8444 8628
rect 8668 8576 8720 8628
rect 11796 8576 11848 8628
rect 12532 8576 12584 8628
rect 15936 8576 15988 8628
rect 3332 8508 3384 8560
rect 3884 8508 3936 8560
rect 2780 8440 2832 8492
rect 4436 8483 4488 8492
rect 4436 8449 4445 8483
rect 4445 8449 4479 8483
rect 4479 8449 4488 8483
rect 4436 8440 4488 8449
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 8576 8508 8628 8560
rect 8484 8440 8536 8492
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 2596 8304 2648 8356
rect 3148 8304 3200 8356
rect 4160 8415 4212 8424
rect 4160 8381 4169 8415
rect 4169 8381 4203 8415
rect 4203 8381 4212 8415
rect 4160 8372 4212 8381
rect 4988 8372 5040 8424
rect 5448 8415 5500 8424
rect 5448 8381 5457 8415
rect 5457 8381 5491 8415
rect 5491 8381 5500 8415
rect 5448 8372 5500 8381
rect 6920 8372 6972 8424
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8760 8372 8812 8381
rect 8852 8372 8904 8424
rect 9680 8440 9732 8492
rect 8668 8304 8720 8356
rect 3516 8236 3568 8288
rect 6092 8236 6144 8288
rect 7288 8236 7340 8288
rect 9404 8279 9456 8288
rect 9404 8245 9413 8279
rect 9413 8245 9447 8279
rect 9447 8245 9456 8279
rect 9404 8236 9456 8245
rect 12164 8508 12216 8560
rect 15660 8508 15712 8560
rect 17960 8551 18012 8560
rect 17960 8517 17969 8551
rect 17969 8517 18003 8551
rect 18003 8517 18012 8551
rect 17960 8508 18012 8517
rect 20076 8619 20128 8628
rect 20076 8585 20085 8619
rect 20085 8585 20119 8619
rect 20119 8585 20128 8619
rect 20076 8576 20128 8585
rect 20352 8576 20404 8628
rect 21732 8576 21784 8628
rect 22560 8576 22612 8628
rect 23664 8576 23716 8628
rect 23388 8508 23440 8560
rect 23848 8508 23900 8560
rect 24492 8619 24544 8628
rect 24492 8585 24501 8619
rect 24501 8585 24535 8619
rect 24535 8585 24544 8619
rect 24492 8576 24544 8585
rect 10232 8440 10284 8492
rect 10784 8440 10836 8492
rect 10968 8415 11020 8424
rect 10968 8381 10977 8415
rect 10977 8381 11011 8415
rect 11011 8381 11020 8415
rect 10968 8372 11020 8381
rect 11244 8415 11296 8424
rect 11244 8381 11253 8415
rect 11253 8381 11287 8415
rect 11287 8381 11296 8415
rect 11244 8372 11296 8381
rect 11336 8415 11388 8424
rect 11336 8381 11345 8415
rect 11345 8381 11379 8415
rect 11379 8381 11388 8415
rect 11336 8372 11388 8381
rect 12716 8440 12768 8492
rect 13360 8440 13412 8492
rect 11796 8415 11848 8424
rect 11796 8381 11810 8415
rect 11810 8381 11844 8415
rect 11844 8381 11848 8415
rect 11796 8372 11848 8381
rect 12164 8372 12216 8424
rect 12348 8372 12400 8424
rect 12900 8415 12952 8424
rect 12900 8381 12909 8415
rect 12909 8381 12943 8415
rect 12943 8381 12952 8415
rect 12900 8372 12952 8381
rect 11060 8304 11112 8356
rect 11612 8347 11664 8356
rect 11612 8313 11621 8347
rect 11621 8313 11655 8347
rect 11655 8313 11664 8347
rect 11612 8304 11664 8313
rect 11980 8304 12032 8356
rect 12624 8304 12676 8356
rect 13636 8372 13688 8424
rect 16304 8440 16356 8492
rect 16488 8483 16540 8492
rect 16488 8449 16497 8483
rect 16497 8449 16531 8483
rect 16531 8449 16540 8483
rect 16488 8440 16540 8449
rect 14372 8372 14424 8424
rect 16764 8415 16816 8424
rect 16764 8381 16773 8415
rect 16773 8381 16807 8415
rect 16807 8381 16816 8415
rect 16764 8372 16816 8381
rect 17592 8440 17644 8492
rect 20168 8440 20220 8492
rect 21732 8483 21784 8492
rect 21732 8449 21741 8483
rect 21741 8449 21775 8483
rect 21775 8449 21784 8483
rect 21732 8440 21784 8449
rect 22468 8440 22520 8492
rect 23756 8440 23808 8492
rect 24676 8551 24728 8560
rect 24676 8517 24685 8551
rect 24685 8517 24719 8551
rect 24719 8517 24728 8551
rect 24676 8508 24728 8517
rect 25412 8440 25464 8492
rect 17776 8372 17828 8424
rect 21824 8372 21876 8424
rect 16488 8304 16540 8356
rect 18788 8304 18840 8356
rect 21088 8304 21140 8356
rect 22008 8304 22060 8356
rect 11336 8236 11388 8288
rect 12072 8236 12124 8288
rect 12348 8279 12400 8288
rect 12348 8245 12357 8279
rect 12357 8245 12391 8279
rect 12391 8245 12400 8279
rect 12348 8236 12400 8245
rect 14188 8279 14240 8288
rect 14188 8245 14197 8279
rect 14197 8245 14231 8279
rect 14231 8245 14240 8279
rect 14188 8236 14240 8245
rect 14832 8236 14884 8288
rect 18328 8279 18380 8288
rect 18328 8245 18337 8279
rect 18337 8245 18371 8279
rect 18371 8245 18380 8279
rect 18328 8236 18380 8245
rect 18604 8236 18656 8288
rect 19524 8236 19576 8288
rect 21364 8236 21416 8288
rect 22468 8304 22520 8356
rect 22652 8415 22704 8424
rect 22652 8381 22661 8415
rect 22661 8381 22695 8415
rect 22695 8381 22704 8415
rect 22652 8372 22704 8381
rect 23480 8372 23532 8424
rect 23388 8236 23440 8288
rect 24768 8347 24820 8356
rect 24768 8313 24777 8347
rect 24777 8313 24811 8347
rect 24811 8313 24820 8347
rect 24768 8304 24820 8313
rect 24860 8304 24912 8356
rect 25412 8347 25464 8356
rect 25412 8313 25437 8347
rect 25437 8313 25464 8347
rect 25412 8304 25464 8313
rect 25596 8304 25648 8356
rect 26884 8304 26936 8356
rect 25780 8236 25832 8288
rect 7114 8134 7166 8186
rect 7178 8134 7230 8186
rect 7242 8134 7294 8186
rect 7306 8134 7358 8186
rect 7370 8134 7422 8186
rect 13830 8134 13882 8186
rect 13894 8134 13946 8186
rect 13958 8134 14010 8186
rect 14022 8134 14074 8186
rect 14086 8134 14138 8186
rect 20546 8134 20598 8186
rect 20610 8134 20662 8186
rect 20674 8134 20726 8186
rect 20738 8134 20790 8186
rect 20802 8134 20854 8186
rect 27262 8134 27314 8186
rect 27326 8134 27378 8186
rect 27390 8134 27442 8186
rect 27454 8134 27506 8186
rect 27518 8134 27570 8186
rect 2596 8075 2648 8084
rect 2596 8041 2605 8075
rect 2605 8041 2639 8075
rect 2639 8041 2648 8075
rect 2596 8032 2648 8041
rect 2780 8075 2832 8084
rect 2780 8041 2789 8075
rect 2789 8041 2823 8075
rect 2823 8041 2832 8075
rect 2780 8032 2832 8041
rect 8760 8032 8812 8084
rect 12808 8032 12860 8084
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 2780 7896 2832 7948
rect 2964 7939 3016 7948
rect 2964 7905 2973 7939
rect 2973 7905 3007 7939
rect 3007 7905 3016 7939
rect 2964 7896 3016 7905
rect 3148 7939 3200 7948
rect 3148 7905 3157 7939
rect 3157 7905 3191 7939
rect 3191 7905 3200 7939
rect 3148 7896 3200 7905
rect 3516 7939 3568 7948
rect 3516 7905 3525 7939
rect 3525 7905 3559 7939
rect 3559 7905 3568 7939
rect 3516 7896 3568 7905
rect 3608 7896 3660 7948
rect 3884 7896 3936 7948
rect 3332 7828 3384 7880
rect 4252 7939 4304 7948
rect 4252 7905 4261 7939
rect 4261 7905 4295 7939
rect 4295 7905 4304 7939
rect 4252 7896 4304 7905
rect 6460 7939 6512 7948
rect 6460 7905 6494 7939
rect 6494 7905 6512 7939
rect 6460 7896 6512 7905
rect 8300 7896 8352 7948
rect 8484 7939 8536 7948
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 8484 7896 8536 7905
rect 9680 7964 9732 8016
rect 5448 7828 5500 7880
rect 6184 7871 6236 7880
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6184 7828 6236 7837
rect 8208 7828 8260 7880
rect 8852 7939 8904 7948
rect 8852 7905 8861 7939
rect 8861 7905 8895 7939
rect 8895 7905 8904 7939
rect 8852 7896 8904 7905
rect 9404 7896 9456 7948
rect 13268 8007 13320 8016
rect 13268 7973 13277 8007
rect 13277 7973 13311 8007
rect 13311 7973 13320 8007
rect 13268 7964 13320 7973
rect 14372 8007 14424 8016
rect 14372 7973 14381 8007
rect 14381 7973 14415 8007
rect 14415 7973 14424 8007
rect 14372 7964 14424 7973
rect 14556 7964 14608 8016
rect 11796 7939 11848 7948
rect 11796 7905 11830 7939
rect 11830 7905 11848 7939
rect 11796 7896 11848 7905
rect 12072 7896 12124 7948
rect 12808 7828 12860 7880
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 13360 7760 13412 7812
rect 14740 7939 14792 7948
rect 14740 7905 14749 7939
rect 14749 7905 14783 7939
rect 14783 7905 14792 7939
rect 14740 7896 14792 7905
rect 14832 7939 14884 7948
rect 14832 7905 14841 7939
rect 14841 7905 14875 7939
rect 14875 7905 14884 7939
rect 14832 7896 14884 7905
rect 15200 7939 15252 7948
rect 18788 8075 18840 8084
rect 18788 8041 18797 8075
rect 18797 8041 18831 8075
rect 18831 8041 18840 8075
rect 18788 8032 18840 8041
rect 20168 8032 20220 8084
rect 20536 8032 20588 8084
rect 15200 7905 15215 7939
rect 15215 7905 15249 7939
rect 15249 7905 15252 7939
rect 15200 7896 15252 7905
rect 15476 7939 15528 7948
rect 15476 7905 15485 7939
rect 15485 7905 15519 7939
rect 15519 7905 15528 7939
rect 15476 7896 15528 7905
rect 16580 7964 16632 8016
rect 17592 7964 17644 8016
rect 20812 8007 20864 8016
rect 14740 7760 14792 7812
rect 3424 7735 3476 7744
rect 3424 7701 3433 7735
rect 3433 7701 3467 7735
rect 3467 7701 3476 7735
rect 3424 7692 3476 7701
rect 4160 7692 4212 7744
rect 7748 7692 7800 7744
rect 8116 7735 8168 7744
rect 8116 7701 8125 7735
rect 8125 7701 8159 7735
rect 8159 7701 8168 7735
rect 8116 7692 8168 7701
rect 8668 7692 8720 7744
rect 11336 7692 11388 7744
rect 11888 7692 11940 7744
rect 13176 7692 13228 7744
rect 15384 7692 15436 7744
rect 18604 7939 18656 7948
rect 18604 7905 18613 7939
rect 18613 7905 18647 7939
rect 18647 7905 18656 7939
rect 18604 7896 18656 7905
rect 20812 7973 20821 8007
rect 20821 7973 20855 8007
rect 20855 7973 20864 8007
rect 20812 7964 20864 7973
rect 19524 7939 19576 7948
rect 19524 7905 19533 7939
rect 19533 7905 19567 7939
rect 19567 7905 19576 7939
rect 19524 7896 19576 7905
rect 20076 7896 20128 7948
rect 18328 7828 18380 7880
rect 19800 7828 19852 7880
rect 18696 7760 18748 7812
rect 20628 7760 20680 7812
rect 21364 7896 21416 7948
rect 21640 7939 21692 7948
rect 21640 7905 21649 7939
rect 21649 7905 21683 7939
rect 21683 7905 21692 7939
rect 21640 7896 21692 7905
rect 22008 8007 22060 8016
rect 22008 7973 22017 8007
rect 22017 7973 22051 8007
rect 22051 7973 22060 8007
rect 22008 7964 22060 7973
rect 23388 7964 23440 8016
rect 21088 7871 21140 7880
rect 21088 7837 21097 7871
rect 21097 7837 21131 7871
rect 21131 7837 21140 7871
rect 21088 7828 21140 7837
rect 22560 7896 22612 7948
rect 23572 7896 23624 7948
rect 24032 8032 24084 8084
rect 24492 8032 24544 8084
rect 24952 8032 25004 8084
rect 24768 7964 24820 8016
rect 23848 7939 23900 7948
rect 23848 7905 23857 7939
rect 23857 7905 23891 7939
rect 23891 7905 23900 7939
rect 23848 7896 23900 7905
rect 24216 7939 24268 7948
rect 24216 7905 24225 7939
rect 24225 7905 24259 7939
rect 24259 7905 24268 7939
rect 24216 7896 24268 7905
rect 24676 7939 24728 7948
rect 24676 7905 24685 7939
rect 24685 7905 24719 7939
rect 24719 7905 24728 7939
rect 24676 7896 24728 7905
rect 22652 7828 22704 7880
rect 23756 7828 23808 7880
rect 22468 7760 22520 7812
rect 23480 7760 23532 7812
rect 25136 7939 25188 7948
rect 25136 7905 25145 7939
rect 25145 7905 25179 7939
rect 25179 7905 25188 7939
rect 25136 7896 25188 7905
rect 25228 7939 25280 7948
rect 25228 7905 25237 7939
rect 25237 7905 25271 7939
rect 25271 7905 25280 7939
rect 25228 7896 25280 7905
rect 17776 7692 17828 7744
rect 22008 7735 22060 7744
rect 22008 7701 22017 7735
rect 22017 7701 22051 7735
rect 22051 7701 22060 7735
rect 22008 7692 22060 7701
rect 23112 7735 23164 7744
rect 23112 7701 23121 7735
rect 23121 7701 23155 7735
rect 23155 7701 23164 7735
rect 23112 7692 23164 7701
rect 24308 7692 24360 7744
rect 24768 7692 24820 7744
rect 3756 7590 3808 7642
rect 3820 7590 3872 7642
rect 3884 7590 3936 7642
rect 3948 7590 4000 7642
rect 4012 7590 4064 7642
rect 10472 7590 10524 7642
rect 10536 7590 10588 7642
rect 10600 7590 10652 7642
rect 10664 7590 10716 7642
rect 10728 7590 10780 7642
rect 17188 7590 17240 7642
rect 17252 7590 17304 7642
rect 17316 7590 17368 7642
rect 17380 7590 17432 7642
rect 17444 7590 17496 7642
rect 23904 7590 23956 7642
rect 23968 7590 24020 7642
rect 24032 7590 24084 7642
rect 24096 7590 24148 7642
rect 24160 7590 24212 7642
rect 4252 7488 4304 7540
rect 5632 7488 5684 7540
rect 3240 7420 3292 7472
rect 3792 7420 3844 7472
rect 4160 7352 4212 7404
rect 6460 7531 6512 7540
rect 6460 7497 6469 7531
rect 6469 7497 6503 7531
rect 6503 7497 6512 7531
rect 6460 7488 6512 7497
rect 9128 7488 9180 7540
rect 11060 7488 11112 7540
rect 11796 7488 11848 7540
rect 13360 7531 13412 7540
rect 13360 7497 13369 7531
rect 13369 7497 13403 7531
rect 13403 7497 13412 7531
rect 13360 7488 13412 7497
rect 13728 7488 13780 7540
rect 15292 7488 15344 7540
rect 18972 7531 19024 7540
rect 13636 7420 13688 7472
rect 18972 7497 18981 7531
rect 18981 7497 19015 7531
rect 19015 7497 19024 7531
rect 18972 7488 19024 7497
rect 19800 7488 19852 7540
rect 21180 7488 21232 7540
rect 23480 7488 23532 7540
rect 24124 7488 24176 7540
rect 26884 7531 26936 7540
rect 26884 7497 26893 7531
rect 26893 7497 26927 7531
rect 26927 7497 26936 7531
rect 26884 7488 26936 7497
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 8852 7395 8904 7404
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 3516 7327 3568 7336
rect 3516 7293 3525 7327
rect 3525 7293 3559 7327
rect 3559 7293 3568 7327
rect 3516 7284 3568 7293
rect 3424 7216 3476 7268
rect 3700 7327 3752 7336
rect 3700 7293 3709 7327
rect 3709 7293 3743 7327
rect 3743 7293 3752 7327
rect 3700 7284 3752 7293
rect 3792 7327 3844 7336
rect 3792 7293 3801 7327
rect 3801 7293 3835 7327
rect 3835 7293 3844 7327
rect 3792 7284 3844 7293
rect 4620 7327 4672 7336
rect 4620 7293 4629 7327
rect 4629 7293 4663 7327
rect 4663 7293 4672 7327
rect 4620 7284 4672 7293
rect 4988 7327 5040 7336
rect 4988 7293 4997 7327
rect 4997 7293 5031 7327
rect 5031 7293 5040 7327
rect 4988 7284 5040 7293
rect 5632 7284 5684 7336
rect 5816 7216 5868 7268
rect 6092 7327 6144 7336
rect 6092 7293 6101 7327
rect 6101 7293 6135 7327
rect 6135 7293 6144 7327
rect 6092 7284 6144 7293
rect 2780 7148 2832 7200
rect 3332 7148 3384 7200
rect 4252 7148 4304 7200
rect 6000 7148 6052 7200
rect 6092 7148 6144 7200
rect 6736 7284 6788 7336
rect 8116 7284 8168 7336
rect 10784 7284 10836 7336
rect 10324 7216 10376 7268
rect 11060 7284 11112 7336
rect 11152 7284 11204 7336
rect 11428 7327 11480 7336
rect 11428 7293 11437 7327
rect 11437 7293 11471 7327
rect 11471 7293 11480 7327
rect 11428 7284 11480 7293
rect 11520 7327 11572 7336
rect 11520 7293 11529 7327
rect 11529 7293 11563 7327
rect 11563 7293 11572 7327
rect 11520 7284 11572 7293
rect 12348 7352 12400 7404
rect 12072 7284 12124 7336
rect 12624 7216 12676 7268
rect 7012 7148 7064 7200
rect 7472 7148 7524 7200
rect 8300 7148 8352 7200
rect 13176 7327 13228 7336
rect 13176 7293 13190 7327
rect 13190 7293 13224 7327
rect 13224 7293 13228 7327
rect 13176 7284 13228 7293
rect 14188 7284 14240 7336
rect 16580 7284 16632 7336
rect 13268 7216 13320 7268
rect 15384 7259 15436 7268
rect 15384 7225 15418 7259
rect 15418 7225 15436 7259
rect 18052 7420 18104 7472
rect 23572 7420 23624 7472
rect 24584 7420 24636 7472
rect 25320 7420 25372 7472
rect 17868 7395 17920 7404
rect 17868 7361 17877 7395
rect 17877 7361 17911 7395
rect 17911 7361 17920 7395
rect 17868 7352 17920 7361
rect 18236 7352 18288 7404
rect 19340 7395 19392 7404
rect 19340 7361 19349 7395
rect 19349 7361 19383 7395
rect 19383 7361 19392 7395
rect 19340 7352 19392 7361
rect 24768 7352 24820 7404
rect 16856 7327 16908 7336
rect 16856 7293 16865 7327
rect 16865 7293 16899 7327
rect 16899 7293 16908 7327
rect 16856 7284 16908 7293
rect 16948 7284 17000 7336
rect 19616 7284 19668 7336
rect 15384 7216 15436 7225
rect 13360 7148 13412 7200
rect 15016 7148 15068 7200
rect 16488 7191 16540 7200
rect 16488 7157 16497 7191
rect 16497 7157 16531 7191
rect 16531 7157 16540 7191
rect 16488 7148 16540 7157
rect 20076 7148 20128 7200
rect 20352 7216 20404 7268
rect 22008 7284 22060 7336
rect 22928 7327 22980 7336
rect 22928 7293 22937 7327
rect 22937 7293 22971 7327
rect 22971 7293 22980 7327
rect 22928 7284 22980 7293
rect 23112 7327 23164 7336
rect 23112 7293 23121 7327
rect 23121 7293 23155 7327
rect 23155 7293 23164 7327
rect 23112 7284 23164 7293
rect 23480 7284 23532 7336
rect 24216 7284 24268 7336
rect 24860 7284 24912 7336
rect 25780 7327 25832 7336
rect 25780 7293 25814 7327
rect 25814 7293 25832 7327
rect 21824 7216 21876 7268
rect 23664 7216 23716 7268
rect 24400 7259 24452 7268
rect 20536 7148 20588 7200
rect 21364 7148 21416 7200
rect 23756 7148 23808 7200
rect 24400 7225 24427 7259
rect 24427 7225 24452 7259
rect 24400 7216 24452 7225
rect 24492 7216 24544 7268
rect 25044 7216 25096 7268
rect 25780 7284 25832 7293
rect 25872 7216 25924 7268
rect 7114 7046 7166 7098
rect 7178 7046 7230 7098
rect 7242 7046 7294 7098
rect 7306 7046 7358 7098
rect 7370 7046 7422 7098
rect 13830 7046 13882 7098
rect 13894 7046 13946 7098
rect 13958 7046 14010 7098
rect 14022 7046 14074 7098
rect 14086 7046 14138 7098
rect 20546 7046 20598 7098
rect 20610 7046 20662 7098
rect 20674 7046 20726 7098
rect 20738 7046 20790 7098
rect 20802 7046 20854 7098
rect 27262 7046 27314 7098
rect 27326 7046 27378 7098
rect 27390 7046 27442 7098
rect 27454 7046 27506 7098
rect 27518 7046 27570 7098
rect 3700 6944 3752 6996
rect 4620 6944 4672 6996
rect 6092 6944 6144 6996
rect 8208 6987 8260 6996
rect 8208 6953 8217 6987
rect 8217 6953 8251 6987
rect 8251 6953 8260 6987
rect 8208 6944 8260 6953
rect 9404 6944 9456 6996
rect 11060 6944 11112 6996
rect 6184 6919 6236 6928
rect 1584 6808 1636 6860
rect 2780 6851 2832 6860
rect 2780 6817 2814 6851
rect 2814 6817 2832 6851
rect 6184 6885 6193 6919
rect 6193 6885 6227 6919
rect 6227 6885 6236 6919
rect 6184 6876 6236 6885
rect 7472 6876 7524 6928
rect 4160 6851 4212 6860
rect 2780 6808 2832 6817
rect 4160 6817 4169 6851
rect 4169 6817 4203 6851
rect 4203 6817 4212 6851
rect 4160 6808 4212 6817
rect 5724 6808 5776 6860
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 8392 6851 8444 6860
rect 8392 6817 8396 6851
rect 8396 6817 8430 6851
rect 8430 6817 8444 6851
rect 8392 6808 8444 6817
rect 8576 6851 8628 6860
rect 8576 6817 8585 6851
rect 8585 6817 8619 6851
rect 8619 6817 8628 6851
rect 8576 6808 8628 6817
rect 8668 6851 8720 6860
rect 8668 6817 8713 6851
rect 8713 6817 8720 6851
rect 8668 6808 8720 6817
rect 8852 6851 8904 6860
rect 8852 6817 8861 6851
rect 8861 6817 8895 6851
rect 8895 6817 8904 6851
rect 8852 6808 8904 6817
rect 8944 6808 8996 6860
rect 9956 6919 10008 6928
rect 9956 6885 9965 6919
rect 9965 6885 9999 6919
rect 9999 6885 10008 6919
rect 9956 6876 10008 6885
rect 10784 6876 10836 6928
rect 9128 6851 9180 6860
rect 9128 6817 9137 6851
rect 9137 6817 9171 6851
rect 9171 6817 9180 6851
rect 9128 6808 9180 6817
rect 9404 6851 9456 6860
rect 9404 6817 9413 6851
rect 9413 6817 9447 6851
rect 9447 6817 9456 6851
rect 9404 6808 9456 6817
rect 7012 6672 7064 6724
rect 5540 6647 5592 6656
rect 5540 6613 5549 6647
rect 5549 6613 5583 6647
rect 5583 6613 5592 6647
rect 5540 6604 5592 6613
rect 6276 6604 6328 6656
rect 9220 6672 9272 6724
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 11428 6944 11480 6996
rect 12256 6944 12308 6996
rect 12808 6944 12860 6996
rect 16488 6944 16540 6996
rect 20260 6944 20312 6996
rect 20628 6944 20680 6996
rect 12716 6876 12768 6928
rect 13176 6876 13228 6928
rect 17776 6876 17828 6928
rect 19616 6876 19668 6928
rect 9864 6740 9916 6792
rect 10416 6740 10468 6792
rect 11428 6740 11480 6792
rect 12900 6808 12952 6860
rect 19340 6808 19392 6860
rect 20076 6808 20128 6860
rect 20996 6876 21048 6928
rect 9588 6715 9640 6724
rect 9588 6681 9597 6715
rect 9597 6681 9631 6715
rect 9631 6681 9640 6715
rect 9588 6672 9640 6681
rect 11244 6672 11296 6724
rect 11704 6672 11756 6724
rect 13084 6783 13136 6792
rect 13084 6749 13093 6783
rect 13093 6749 13127 6783
rect 13127 6749 13136 6783
rect 13084 6740 13136 6749
rect 13452 6740 13504 6792
rect 17592 6783 17644 6792
rect 17592 6749 17601 6783
rect 17601 6749 17635 6783
rect 17635 6749 17644 6783
rect 17592 6740 17644 6749
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 20812 6851 20864 6860
rect 20812 6817 20821 6851
rect 20821 6817 20855 6851
rect 20855 6817 20864 6851
rect 20812 6808 20864 6817
rect 20904 6851 20956 6860
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 24400 6944 24452 6996
rect 25872 6987 25924 6996
rect 24308 6876 24360 6928
rect 25872 6953 25881 6987
rect 25881 6953 25915 6987
rect 25915 6953 25924 6987
rect 25872 6944 25924 6953
rect 20444 6740 20496 6792
rect 9496 6604 9548 6656
rect 10140 6647 10192 6656
rect 10140 6613 10149 6647
rect 10149 6613 10183 6647
rect 10183 6613 10192 6647
rect 10140 6604 10192 6613
rect 10232 6647 10284 6656
rect 10232 6613 10241 6647
rect 10241 6613 10275 6647
rect 10275 6613 10284 6647
rect 10232 6604 10284 6613
rect 10416 6604 10468 6656
rect 11060 6604 11112 6656
rect 12164 6604 12216 6656
rect 16304 6604 16356 6656
rect 18328 6604 18380 6656
rect 23572 6808 23624 6860
rect 24124 6851 24176 6860
rect 24124 6817 24133 6851
rect 24133 6817 24167 6851
rect 24167 6817 24176 6851
rect 24124 6808 24176 6817
rect 24584 6808 24636 6860
rect 24768 6851 24820 6860
rect 24768 6817 24802 6851
rect 24802 6817 24820 6851
rect 24768 6808 24820 6817
rect 25872 6740 25924 6792
rect 19340 6604 19392 6656
rect 19708 6604 19760 6656
rect 20076 6604 20128 6656
rect 20260 6604 20312 6656
rect 24400 6672 24452 6724
rect 22376 6604 22428 6656
rect 24308 6604 24360 6656
rect 3756 6502 3808 6554
rect 3820 6502 3872 6554
rect 3884 6502 3936 6554
rect 3948 6502 4000 6554
rect 4012 6502 4064 6554
rect 10472 6502 10524 6554
rect 10536 6502 10588 6554
rect 10600 6502 10652 6554
rect 10664 6502 10716 6554
rect 10728 6502 10780 6554
rect 17188 6502 17240 6554
rect 17252 6502 17304 6554
rect 17316 6502 17368 6554
rect 17380 6502 17432 6554
rect 17444 6502 17496 6554
rect 23904 6502 23956 6554
rect 23968 6502 24020 6554
rect 24032 6502 24084 6554
rect 24096 6502 24148 6554
rect 24160 6502 24212 6554
rect 4988 6443 5040 6452
rect 4988 6409 4997 6443
rect 4997 6409 5031 6443
rect 5031 6409 5040 6443
rect 4988 6400 5040 6409
rect 5448 6400 5500 6452
rect 5540 6375 5592 6384
rect 5540 6341 5549 6375
rect 5549 6341 5583 6375
rect 5583 6341 5592 6375
rect 5540 6332 5592 6341
rect 5816 6443 5868 6452
rect 5816 6409 5825 6443
rect 5825 6409 5859 6443
rect 5859 6409 5868 6443
rect 5816 6400 5868 6409
rect 9036 6400 9088 6452
rect 10048 6400 10100 6452
rect 10324 6443 10376 6452
rect 10324 6409 10333 6443
rect 10333 6409 10367 6443
rect 10367 6409 10376 6443
rect 10324 6400 10376 6409
rect 11244 6443 11296 6452
rect 11244 6409 11253 6443
rect 11253 6409 11287 6443
rect 11287 6409 11296 6443
rect 11244 6400 11296 6409
rect 11336 6400 11388 6452
rect 14556 6400 14608 6452
rect 17684 6443 17736 6452
rect 17684 6409 17693 6443
rect 17693 6409 17727 6443
rect 17727 6409 17736 6443
rect 17684 6400 17736 6409
rect 19616 6400 19668 6452
rect 6184 6332 6236 6384
rect 6276 6307 6328 6316
rect 6276 6273 6285 6307
rect 6285 6273 6319 6307
rect 6319 6273 6328 6307
rect 6276 6264 6328 6273
rect 3516 6196 3568 6248
rect 4620 6128 4672 6180
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 7564 6196 7616 6248
rect 7748 6196 7800 6248
rect 8208 6239 8260 6248
rect 8208 6205 8217 6239
rect 8217 6205 8251 6239
rect 8251 6205 8260 6239
rect 8208 6196 8260 6205
rect 9588 6332 9640 6384
rect 10232 6264 10284 6316
rect 10324 6264 10376 6316
rect 11060 6307 11112 6316
rect 11060 6273 11069 6307
rect 11069 6273 11103 6307
rect 11103 6273 11112 6307
rect 11060 6264 11112 6273
rect 9956 6196 10008 6248
rect 10048 6196 10100 6248
rect 10968 6196 11020 6248
rect 11336 6239 11388 6248
rect 11336 6205 11345 6239
rect 11345 6205 11379 6239
rect 11379 6205 11388 6239
rect 11336 6196 11388 6205
rect 19984 6332 20036 6384
rect 8576 6103 8628 6112
rect 8576 6069 8585 6103
rect 8585 6069 8619 6103
rect 8619 6069 8628 6103
rect 8576 6060 8628 6069
rect 9496 6060 9548 6112
rect 10784 6103 10836 6112
rect 10784 6069 10793 6103
rect 10793 6069 10827 6103
rect 10827 6069 10836 6103
rect 10784 6060 10836 6069
rect 13820 6196 13872 6248
rect 16396 6264 16448 6316
rect 17592 6264 17644 6316
rect 18144 6264 18196 6316
rect 21272 6400 21324 6452
rect 20904 6332 20956 6384
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 23480 6400 23532 6409
rect 23756 6400 23808 6452
rect 25228 6400 25280 6452
rect 25872 6443 25924 6452
rect 25872 6409 25881 6443
rect 25881 6409 25915 6443
rect 25915 6409 25924 6443
rect 25872 6400 25924 6409
rect 14280 6196 14332 6248
rect 16948 6196 17000 6248
rect 18052 6239 18104 6248
rect 18052 6205 18061 6239
rect 18061 6205 18095 6239
rect 18095 6205 18104 6239
rect 18052 6196 18104 6205
rect 11428 6060 11480 6112
rect 11520 6103 11572 6112
rect 11520 6069 11529 6103
rect 11529 6069 11563 6103
rect 11563 6069 11572 6103
rect 11520 6060 11572 6069
rect 11612 6060 11664 6112
rect 12256 6060 12308 6112
rect 15660 6128 15712 6180
rect 15844 6060 15896 6112
rect 16856 6128 16908 6180
rect 18328 6196 18380 6248
rect 18420 6239 18472 6248
rect 18420 6205 18429 6239
rect 18429 6205 18463 6239
rect 18463 6205 18472 6239
rect 18420 6196 18472 6205
rect 18604 6196 18656 6248
rect 20444 6239 20496 6248
rect 20444 6205 20453 6239
rect 20453 6205 20487 6239
rect 20487 6205 20496 6239
rect 20444 6196 20496 6205
rect 21272 6264 21324 6316
rect 23388 6307 23440 6316
rect 23388 6273 23397 6307
rect 23397 6273 23431 6307
rect 23431 6273 23440 6307
rect 23388 6264 23440 6273
rect 24492 6307 24544 6316
rect 24492 6273 24501 6307
rect 24501 6273 24535 6307
rect 24535 6273 24544 6307
rect 24492 6264 24544 6273
rect 20812 6239 20864 6248
rect 20812 6205 20821 6239
rect 20821 6205 20855 6239
rect 20855 6205 20864 6239
rect 20812 6196 20864 6205
rect 21364 6196 21416 6248
rect 21824 6196 21876 6248
rect 22376 6239 22428 6248
rect 22376 6205 22385 6239
rect 22385 6205 22419 6239
rect 22419 6205 22428 6239
rect 22376 6196 22428 6205
rect 23480 6196 23532 6248
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 21088 6128 21140 6180
rect 21272 6128 21324 6180
rect 22008 6128 22060 6180
rect 22744 6128 22796 6180
rect 22836 6128 22888 6180
rect 24308 6239 24360 6248
rect 24308 6205 24317 6239
rect 24317 6205 24351 6239
rect 24351 6205 24360 6239
rect 24308 6196 24360 6205
rect 24216 6128 24268 6180
rect 24584 6128 24636 6180
rect 24768 6171 24820 6180
rect 24768 6137 24802 6171
rect 24802 6137 24820 6171
rect 24768 6128 24820 6137
rect 17960 6060 18012 6112
rect 20628 6060 20680 6112
rect 22560 6060 22612 6112
rect 7114 5958 7166 6010
rect 7178 5958 7230 6010
rect 7242 5958 7294 6010
rect 7306 5958 7358 6010
rect 7370 5958 7422 6010
rect 13830 5958 13882 6010
rect 13894 5958 13946 6010
rect 13958 5958 14010 6010
rect 14022 5958 14074 6010
rect 14086 5958 14138 6010
rect 20546 5958 20598 6010
rect 20610 5958 20662 6010
rect 20674 5958 20726 6010
rect 20738 5958 20790 6010
rect 20802 5958 20854 6010
rect 27262 5958 27314 6010
rect 27326 5958 27378 6010
rect 27390 5958 27442 6010
rect 27454 5958 27506 6010
rect 27518 5958 27570 6010
rect 4344 5856 4396 5908
rect 5724 5856 5776 5908
rect 7748 5899 7800 5908
rect 7748 5865 7757 5899
rect 7757 5865 7791 5899
rect 7791 5865 7800 5899
rect 7748 5856 7800 5865
rect 9680 5856 9732 5908
rect 11336 5856 11388 5908
rect 12164 5856 12216 5908
rect 12256 5899 12308 5908
rect 12256 5865 12265 5899
rect 12265 5865 12299 5899
rect 12299 5865 12308 5899
rect 12256 5856 12308 5865
rect 12992 5856 13044 5908
rect 13820 5856 13872 5908
rect 14188 5856 14240 5908
rect 15108 5899 15160 5908
rect 15108 5865 15117 5899
rect 15117 5865 15151 5899
rect 15151 5865 15160 5899
rect 15108 5856 15160 5865
rect 16120 5856 16172 5908
rect 17684 5856 17736 5908
rect 6736 5788 6788 5840
rect 8208 5788 8260 5840
rect 10140 5788 10192 5840
rect 10876 5788 10928 5840
rect 4252 5720 4304 5772
rect 5172 5720 5224 5772
rect 5264 5720 5316 5772
rect 5448 5720 5500 5772
rect 6000 5763 6052 5772
rect 6000 5729 6009 5763
rect 6009 5729 6043 5763
rect 6043 5729 6052 5763
rect 6000 5720 6052 5729
rect 4528 5652 4580 5704
rect 5080 5652 5132 5704
rect 5356 5584 5408 5636
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 8852 5720 8904 5772
rect 9496 5720 9548 5772
rect 10968 5763 11020 5772
rect 10968 5729 10977 5763
rect 10977 5729 11011 5763
rect 11011 5729 11020 5763
rect 10968 5720 11020 5729
rect 12532 5788 12584 5840
rect 13360 5788 13412 5840
rect 15016 5788 15068 5840
rect 18420 5788 18472 5840
rect 19892 5856 19944 5908
rect 20352 5856 20404 5908
rect 21180 5856 21232 5908
rect 21364 5899 21416 5908
rect 21364 5865 21373 5899
rect 21373 5865 21407 5899
rect 21407 5865 21416 5899
rect 21364 5856 21416 5865
rect 9036 5652 9088 5704
rect 3332 5516 3384 5568
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 8852 5584 8904 5636
rect 10784 5584 10836 5636
rect 11612 5516 11664 5568
rect 11704 5559 11756 5568
rect 11704 5525 11713 5559
rect 11713 5525 11747 5559
rect 11747 5525 11756 5559
rect 11704 5516 11756 5525
rect 12808 5720 12860 5772
rect 13452 5763 13504 5772
rect 13452 5729 13461 5763
rect 13461 5729 13495 5763
rect 13495 5729 13504 5763
rect 13452 5720 13504 5729
rect 14188 5720 14240 5772
rect 14556 5720 14608 5772
rect 15384 5720 15436 5772
rect 15844 5720 15896 5772
rect 18052 5763 18104 5772
rect 18052 5729 18086 5763
rect 18086 5729 18104 5763
rect 18052 5720 18104 5729
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 12716 5652 12768 5661
rect 12992 5652 13044 5704
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 15200 5695 15252 5704
rect 15200 5661 15209 5695
rect 15209 5661 15243 5695
rect 15243 5661 15252 5695
rect 15200 5652 15252 5661
rect 15660 5652 15712 5704
rect 16856 5652 16908 5704
rect 14280 5516 14332 5568
rect 16856 5516 16908 5568
rect 19524 5720 19576 5772
rect 22744 5899 22796 5908
rect 22744 5865 22753 5899
rect 22753 5865 22787 5899
rect 22787 5865 22796 5899
rect 22744 5856 22796 5865
rect 24768 5856 24820 5908
rect 25136 5856 25188 5908
rect 24584 5788 24636 5840
rect 19984 5720 20036 5772
rect 20260 5720 20312 5772
rect 23572 5720 23624 5772
rect 24216 5720 24268 5772
rect 25136 5720 25188 5772
rect 21180 5652 21232 5704
rect 21916 5695 21968 5704
rect 21916 5661 21925 5695
rect 21925 5661 21959 5695
rect 21959 5661 21968 5695
rect 21916 5652 21968 5661
rect 20996 5584 21048 5636
rect 22376 5695 22428 5704
rect 22376 5661 22385 5695
rect 22385 5661 22419 5695
rect 22419 5661 22428 5695
rect 22376 5652 22428 5661
rect 18144 5516 18196 5568
rect 21456 5516 21508 5568
rect 22100 5516 22152 5568
rect 22560 5695 22612 5704
rect 22560 5661 22569 5695
rect 22569 5661 22603 5695
rect 22603 5661 22612 5695
rect 22560 5652 22612 5661
rect 26056 5720 26108 5772
rect 24216 5584 24268 5636
rect 23756 5516 23808 5568
rect 25136 5559 25188 5568
rect 25136 5525 25145 5559
rect 25145 5525 25179 5559
rect 25179 5525 25188 5559
rect 25136 5516 25188 5525
rect 3756 5414 3808 5466
rect 3820 5414 3872 5466
rect 3884 5414 3936 5466
rect 3948 5414 4000 5466
rect 4012 5414 4064 5466
rect 10472 5414 10524 5466
rect 10536 5414 10588 5466
rect 10600 5414 10652 5466
rect 10664 5414 10716 5466
rect 10728 5414 10780 5466
rect 17188 5414 17240 5466
rect 17252 5414 17304 5466
rect 17316 5414 17368 5466
rect 17380 5414 17432 5466
rect 17444 5414 17496 5466
rect 23904 5414 23956 5466
rect 23968 5414 24020 5466
rect 24032 5414 24084 5466
rect 24096 5414 24148 5466
rect 24160 5414 24212 5466
rect 6736 5312 6788 5364
rect 4160 5219 4212 5228
rect 4160 5185 4169 5219
rect 4169 5185 4203 5219
rect 4203 5185 4212 5219
rect 4160 5176 4212 5185
rect 5172 5176 5224 5228
rect 4712 5040 4764 5092
rect 6368 5108 6420 5160
rect 5540 5015 5592 5024
rect 5540 4981 5549 5015
rect 5549 4981 5583 5015
rect 5583 4981 5592 5015
rect 5540 4972 5592 4981
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 5632 4972 5684 4981
rect 8668 5312 8720 5364
rect 9956 5312 10008 5364
rect 10048 5355 10100 5364
rect 10048 5321 10057 5355
rect 10057 5321 10091 5355
rect 10091 5321 10100 5355
rect 10048 5312 10100 5321
rect 12900 5312 12952 5364
rect 13728 5312 13780 5364
rect 15752 5312 15804 5364
rect 8392 5108 8444 5160
rect 9128 5108 9180 5160
rect 9680 5108 9732 5160
rect 10876 5108 10928 5160
rect 8300 5040 8352 5092
rect 8576 5040 8628 5092
rect 11520 5040 11572 5092
rect 7748 4972 7800 5024
rect 8484 4972 8536 5024
rect 9404 4972 9456 5024
rect 16212 5244 16264 5296
rect 12624 5108 12676 5160
rect 14280 5108 14332 5160
rect 14464 5108 14516 5160
rect 15016 5108 15068 5160
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 12992 5040 13044 5092
rect 16028 5108 16080 5160
rect 18052 5312 18104 5364
rect 18144 5244 18196 5296
rect 17960 5176 18012 5228
rect 16856 5151 16908 5160
rect 16856 5117 16890 5151
rect 16890 5117 16908 5151
rect 16856 5108 16908 5117
rect 19892 5151 19944 5160
rect 19892 5117 19901 5151
rect 19901 5117 19935 5151
rect 19935 5117 19944 5151
rect 19892 5108 19944 5117
rect 20812 5312 20864 5364
rect 21916 5312 21968 5364
rect 23572 5355 23624 5364
rect 23572 5321 23581 5355
rect 23581 5321 23615 5355
rect 23615 5321 23624 5355
rect 23572 5312 23624 5321
rect 24492 5312 24544 5364
rect 26056 5312 26108 5364
rect 20996 5108 21048 5160
rect 21824 5108 21876 5160
rect 23756 5244 23808 5296
rect 23388 5219 23440 5228
rect 23388 5185 23397 5219
rect 23397 5185 23431 5219
rect 23431 5185 23440 5219
rect 23388 5176 23440 5185
rect 23480 5176 23532 5228
rect 11888 4972 11940 5024
rect 16672 5040 16724 5092
rect 23756 5108 23808 5160
rect 19156 4972 19208 5024
rect 25412 5040 25464 5092
rect 7114 4870 7166 4922
rect 7178 4870 7230 4922
rect 7242 4870 7294 4922
rect 7306 4870 7358 4922
rect 7370 4870 7422 4922
rect 13830 4870 13882 4922
rect 13894 4870 13946 4922
rect 13958 4870 14010 4922
rect 14022 4870 14074 4922
rect 14086 4870 14138 4922
rect 20546 4870 20598 4922
rect 20610 4870 20662 4922
rect 20674 4870 20726 4922
rect 20738 4870 20790 4922
rect 20802 4870 20854 4922
rect 27262 4870 27314 4922
rect 27326 4870 27378 4922
rect 27390 4870 27442 4922
rect 27454 4870 27506 4922
rect 27518 4870 27570 4922
rect 4528 4768 4580 4820
rect 4712 4811 4764 4820
rect 4712 4777 4721 4811
rect 4721 4777 4755 4811
rect 4755 4777 4764 4811
rect 4712 4768 4764 4777
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 8484 4811 8536 4820
rect 8484 4777 8493 4811
rect 8493 4777 8527 4811
rect 8527 4777 8536 4811
rect 8484 4768 8536 4777
rect 4160 4700 4212 4752
rect 3332 4675 3384 4684
rect 3332 4641 3366 4675
rect 3366 4641 3384 4675
rect 3332 4632 3384 4641
rect 5632 4700 5684 4752
rect 4344 4564 4396 4616
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 5264 4632 5316 4684
rect 6736 4564 6788 4616
rect 7472 4428 7524 4480
rect 7748 4675 7800 4684
rect 7748 4641 7757 4675
rect 7757 4641 7791 4675
rect 7791 4641 7800 4675
rect 7748 4632 7800 4641
rect 8392 4700 8444 4752
rect 10048 4632 10100 4684
rect 12072 4700 12124 4752
rect 12624 4768 12676 4820
rect 13176 4768 13228 4820
rect 14188 4768 14240 4820
rect 14372 4768 14424 4820
rect 13360 4700 13412 4752
rect 8668 4564 8720 4616
rect 9864 4564 9916 4616
rect 10784 4675 10836 4684
rect 10784 4641 10793 4675
rect 10793 4641 10827 4675
rect 10827 4641 10836 4675
rect 10784 4632 10836 4641
rect 10876 4632 10928 4684
rect 12164 4632 12216 4684
rect 12532 4632 12584 4684
rect 12900 4675 12952 4684
rect 12900 4641 12909 4675
rect 12909 4641 12943 4675
rect 12943 4641 12952 4675
rect 12900 4632 12952 4641
rect 14372 4632 14424 4684
rect 15384 4700 15436 4752
rect 16396 4743 16448 4752
rect 16396 4709 16405 4743
rect 16405 4709 16439 4743
rect 16439 4709 16448 4743
rect 16396 4700 16448 4709
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 15016 4564 15068 4616
rect 16580 4675 16632 4684
rect 16580 4641 16589 4675
rect 16589 4641 16623 4675
rect 16623 4641 16632 4675
rect 16580 4632 16632 4641
rect 19616 4768 19668 4820
rect 23756 4811 23808 4820
rect 23756 4777 23765 4811
rect 23765 4777 23799 4811
rect 23799 4777 23808 4811
rect 23756 4768 23808 4777
rect 24676 4768 24728 4820
rect 17040 4743 17092 4752
rect 17040 4709 17049 4743
rect 17049 4709 17083 4743
rect 17083 4709 17092 4743
rect 17040 4700 17092 4709
rect 17132 4743 17184 4752
rect 17132 4709 17141 4743
rect 17141 4709 17175 4743
rect 17175 4709 17184 4743
rect 17132 4700 17184 4709
rect 24584 4743 24636 4752
rect 24584 4709 24593 4743
rect 24593 4709 24627 4743
rect 24627 4709 24636 4743
rect 24584 4700 24636 4709
rect 8116 4539 8168 4548
rect 8116 4505 8125 4539
rect 8125 4505 8159 4539
rect 8159 4505 8168 4539
rect 8116 4496 8168 4505
rect 10784 4496 10836 4548
rect 18604 4607 18656 4616
rect 18604 4573 18613 4607
rect 18613 4573 18647 4607
rect 18647 4573 18656 4607
rect 18604 4564 18656 4573
rect 10140 4471 10192 4480
rect 10140 4437 10149 4471
rect 10149 4437 10183 4471
rect 10183 4437 10192 4471
rect 10140 4428 10192 4437
rect 10968 4428 11020 4480
rect 16764 4471 16816 4480
rect 16764 4437 16773 4471
rect 16773 4437 16807 4471
rect 16807 4437 16816 4471
rect 16764 4428 16816 4437
rect 24400 4675 24452 4684
rect 24400 4641 24409 4675
rect 24409 4641 24443 4675
rect 24443 4641 24452 4675
rect 24400 4632 24452 4641
rect 25412 4768 25464 4820
rect 19524 4496 19576 4548
rect 19340 4428 19392 4480
rect 25136 4428 25188 4480
rect 3756 4326 3808 4378
rect 3820 4326 3872 4378
rect 3884 4326 3936 4378
rect 3948 4326 4000 4378
rect 4012 4326 4064 4378
rect 10472 4326 10524 4378
rect 10536 4326 10588 4378
rect 10600 4326 10652 4378
rect 10664 4326 10716 4378
rect 10728 4326 10780 4378
rect 17188 4326 17240 4378
rect 17252 4326 17304 4378
rect 17316 4326 17368 4378
rect 17380 4326 17432 4378
rect 17444 4326 17496 4378
rect 23904 4326 23956 4378
rect 23968 4326 24020 4378
rect 24032 4326 24084 4378
rect 24096 4326 24148 4378
rect 24160 4326 24212 4378
rect 4160 4088 4212 4140
rect 2780 3952 2832 4004
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 4068 4063 4120 4072
rect 4068 4029 4077 4063
rect 4077 4029 4111 4063
rect 4111 4029 4120 4063
rect 4068 4020 4120 4029
rect 4528 4088 4580 4140
rect 5540 4224 5592 4276
rect 10048 4267 10100 4276
rect 10048 4233 10057 4267
rect 10057 4233 10091 4267
rect 10091 4233 10100 4267
rect 10048 4224 10100 4233
rect 12164 4267 12216 4276
rect 12164 4233 12173 4267
rect 12173 4233 12207 4267
rect 12207 4233 12216 4267
rect 12164 4224 12216 4233
rect 16580 4224 16632 4276
rect 17040 4224 17092 4276
rect 19616 4267 19668 4276
rect 19616 4233 19625 4267
rect 19625 4233 19659 4267
rect 19659 4233 19668 4267
rect 19616 4224 19668 4233
rect 19984 4224 20036 4276
rect 6920 4156 6972 4208
rect 8116 4156 8168 4208
rect 8668 4156 8720 4208
rect 12532 4156 12584 4208
rect 4620 4020 4672 4072
rect 4712 4063 4764 4072
rect 4712 4029 4721 4063
rect 4721 4029 4755 4063
rect 4755 4029 4764 4063
rect 4712 4020 4764 4029
rect 5540 4088 5592 4140
rect 5908 4088 5960 4140
rect 3424 3927 3476 3936
rect 3424 3893 3433 3927
rect 3433 3893 3467 3927
rect 3467 3893 3476 3927
rect 3424 3884 3476 3893
rect 5080 4063 5132 4072
rect 5080 4029 5089 4063
rect 5089 4029 5123 4063
rect 5123 4029 5132 4063
rect 5080 4020 5132 4029
rect 4988 3952 5040 4004
rect 6736 4063 6788 4072
rect 6736 4029 6745 4063
rect 6745 4029 6779 4063
rect 6779 4029 6788 4063
rect 6736 4020 6788 4029
rect 6920 4020 6972 4072
rect 7564 4020 7616 4072
rect 7656 4063 7708 4072
rect 7656 4029 7665 4063
rect 7665 4029 7699 4063
rect 7699 4029 7708 4063
rect 7656 4020 7708 4029
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 8668 4063 8720 4072
rect 8668 4029 8677 4063
rect 8677 4029 8711 4063
rect 8711 4029 8720 4063
rect 8668 4020 8720 4029
rect 10692 4063 10744 4072
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 10692 4020 10744 4029
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 10968 4063 11020 4072
rect 10968 4029 10977 4063
rect 10977 4029 11011 4063
rect 11011 4029 11020 4063
rect 10968 4020 11020 4029
rect 11060 4063 11112 4072
rect 11060 4029 11072 4063
rect 11072 4029 11106 4063
rect 11106 4029 11112 4063
rect 11060 4020 11112 4029
rect 12348 4088 12400 4140
rect 11520 4063 11572 4072
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 11704 4063 11756 4072
rect 11704 4029 11713 4063
rect 11713 4029 11747 4063
rect 11747 4029 11756 4063
rect 11704 4020 11756 4029
rect 11796 4063 11848 4072
rect 11796 4029 11805 4063
rect 11805 4029 11839 4063
rect 11839 4029 11848 4063
rect 11796 4020 11848 4029
rect 11888 4063 11940 4072
rect 11888 4029 11897 4063
rect 11897 4029 11931 4063
rect 11931 4029 11940 4063
rect 11888 4020 11940 4029
rect 16764 4156 16816 4208
rect 16396 4088 16448 4140
rect 16948 4156 17000 4208
rect 17316 4156 17368 4208
rect 17684 4156 17736 4208
rect 18604 4156 18656 4208
rect 14188 4020 14240 4072
rect 12072 3952 12124 4004
rect 12256 3952 12308 4004
rect 12348 3952 12400 4004
rect 14372 3952 14424 4004
rect 15108 4020 15160 4072
rect 15292 3952 15344 4004
rect 15660 3952 15712 4004
rect 17040 4063 17092 4072
rect 17040 4029 17049 4063
rect 17049 4029 17083 4063
rect 17083 4029 17092 4063
rect 17040 4020 17092 4029
rect 17316 4063 17368 4072
rect 17316 4029 17325 4063
rect 17325 4029 17359 4063
rect 17359 4029 17368 4063
rect 17316 4020 17368 4029
rect 16764 3952 16816 4004
rect 19340 4063 19392 4072
rect 19340 4029 19349 4063
rect 19349 4029 19383 4063
rect 19383 4029 19392 4063
rect 19340 4020 19392 4029
rect 20996 4131 21048 4140
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 24584 4020 24636 4072
rect 3976 3884 4028 3936
rect 5264 3927 5316 3936
rect 5264 3893 5273 3927
rect 5273 3893 5307 3927
rect 5307 3893 5316 3927
rect 5264 3884 5316 3893
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 9588 3884 9640 3936
rect 10784 3884 10836 3936
rect 11336 3884 11388 3936
rect 11428 3927 11480 3936
rect 11428 3893 11437 3927
rect 11437 3893 11471 3927
rect 11471 3893 11480 3927
rect 11428 3884 11480 3893
rect 12808 3884 12860 3936
rect 18052 3927 18104 3936
rect 18052 3893 18061 3927
rect 18061 3893 18095 3927
rect 18095 3893 18104 3927
rect 18052 3884 18104 3893
rect 19432 3884 19484 3936
rect 23020 3952 23072 4004
rect 7114 3782 7166 3834
rect 7178 3782 7230 3834
rect 7242 3782 7294 3834
rect 7306 3782 7358 3834
rect 7370 3782 7422 3834
rect 13830 3782 13882 3834
rect 13894 3782 13946 3834
rect 13958 3782 14010 3834
rect 14022 3782 14074 3834
rect 14086 3782 14138 3834
rect 20546 3782 20598 3834
rect 20610 3782 20662 3834
rect 20674 3782 20726 3834
rect 20738 3782 20790 3834
rect 20802 3782 20854 3834
rect 27262 3782 27314 3834
rect 27326 3782 27378 3834
rect 27390 3782 27442 3834
rect 27454 3782 27506 3834
rect 27518 3782 27570 3834
rect 2780 3723 2832 3732
rect 2780 3689 2789 3723
rect 2789 3689 2823 3723
rect 2823 3689 2832 3723
rect 2780 3680 2832 3689
rect 4068 3680 4120 3732
rect 4712 3680 4764 3732
rect 4804 3680 4856 3732
rect 7840 3680 7892 3732
rect 10692 3680 10744 3732
rect 10968 3680 11020 3732
rect 12256 3680 12308 3732
rect 12716 3680 12768 3732
rect 15108 3680 15160 3732
rect 15200 3723 15252 3732
rect 15200 3689 15209 3723
rect 15209 3689 15243 3723
rect 15243 3689 15252 3723
rect 15200 3680 15252 3689
rect 16028 3680 16080 3732
rect 16488 3723 16540 3732
rect 16488 3689 16497 3723
rect 16497 3689 16531 3723
rect 16531 3689 16540 3723
rect 16488 3680 16540 3689
rect 16764 3680 16816 3732
rect 4160 3612 4212 3664
rect 5448 3612 5500 3664
rect 3424 3544 3476 3596
rect 3976 3587 4028 3596
rect 3976 3553 3985 3587
rect 3985 3553 4019 3587
rect 4019 3553 4028 3587
rect 3976 3544 4028 3553
rect 5816 3544 5868 3596
rect 6368 3612 6420 3664
rect 9036 3544 9088 3596
rect 9128 3587 9180 3596
rect 9128 3553 9137 3587
rect 9137 3553 9171 3587
rect 9171 3553 9180 3587
rect 9404 3587 9456 3596
rect 9128 3544 9180 3553
rect 9404 3553 9413 3587
rect 9413 3553 9447 3587
rect 9447 3553 9456 3587
rect 9404 3544 9456 3553
rect 10140 3544 10192 3596
rect 11428 3612 11480 3664
rect 12072 3612 12124 3664
rect 13268 3612 13320 3664
rect 13636 3612 13688 3664
rect 15844 3612 15896 3664
rect 17040 3612 17092 3664
rect 11520 3544 11572 3596
rect 3792 3476 3844 3528
rect 12256 3544 12308 3596
rect 12716 3587 12768 3596
rect 12716 3553 12725 3587
rect 12725 3553 12759 3587
rect 12759 3553 12768 3587
rect 12716 3544 12768 3553
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 12992 3587 13044 3596
rect 12992 3553 13001 3587
rect 13001 3553 13035 3587
rect 13035 3553 13044 3587
rect 12992 3544 13044 3553
rect 3608 3340 3660 3392
rect 14004 3476 14056 3528
rect 14188 3519 14240 3528
rect 14188 3485 14197 3519
rect 14197 3485 14231 3519
rect 14231 3485 14240 3519
rect 14188 3476 14240 3485
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 15660 3519 15712 3528
rect 15660 3485 15669 3519
rect 15669 3485 15703 3519
rect 15703 3485 15712 3519
rect 15660 3476 15712 3485
rect 16948 3587 17000 3596
rect 16948 3553 16957 3587
rect 16957 3553 16991 3587
rect 16991 3553 17000 3587
rect 16948 3544 17000 3553
rect 7840 3408 7892 3460
rect 5356 3340 5408 3392
rect 5632 3383 5684 3392
rect 5632 3349 5641 3383
rect 5641 3349 5675 3383
rect 5675 3349 5684 3383
rect 5632 3340 5684 3349
rect 7656 3340 7708 3392
rect 7932 3340 7984 3392
rect 15476 3408 15528 3460
rect 16856 3476 16908 3528
rect 12348 3340 12400 3392
rect 12532 3340 12584 3392
rect 13176 3340 13228 3392
rect 16028 3408 16080 3460
rect 16396 3408 16448 3460
rect 16672 3408 16724 3460
rect 17776 3612 17828 3664
rect 18052 3612 18104 3664
rect 19524 3723 19576 3732
rect 19524 3689 19533 3723
rect 19533 3689 19567 3723
rect 19567 3689 19576 3723
rect 19524 3680 19576 3689
rect 19892 3612 19944 3664
rect 17960 3544 18012 3596
rect 19800 3544 19852 3596
rect 20444 3544 20496 3596
rect 20996 3587 21048 3596
rect 20996 3553 21005 3587
rect 21005 3553 21039 3587
rect 21039 3553 21048 3587
rect 20996 3544 21048 3553
rect 17684 3519 17736 3528
rect 17684 3485 17693 3519
rect 17693 3485 17727 3519
rect 17727 3485 17736 3519
rect 17684 3476 17736 3485
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 18328 3340 18380 3392
rect 3756 3238 3808 3290
rect 3820 3238 3872 3290
rect 3884 3238 3936 3290
rect 3948 3238 4000 3290
rect 4012 3238 4064 3290
rect 10472 3238 10524 3290
rect 10536 3238 10588 3290
rect 10600 3238 10652 3290
rect 10664 3238 10716 3290
rect 10728 3238 10780 3290
rect 17188 3238 17240 3290
rect 17252 3238 17304 3290
rect 17316 3238 17368 3290
rect 17380 3238 17432 3290
rect 17444 3238 17496 3290
rect 23904 3238 23956 3290
rect 23968 3238 24020 3290
rect 24032 3238 24084 3290
rect 24096 3238 24148 3290
rect 24160 3238 24212 3290
rect 4160 3136 4212 3188
rect 5080 3136 5132 3188
rect 5816 3136 5868 3188
rect 6736 3136 6788 3188
rect 8944 3136 8996 3188
rect 9036 3136 9088 3188
rect 4712 3068 4764 3120
rect 5724 3068 5776 3120
rect 6736 3000 6788 3052
rect 8852 3068 8904 3120
rect 9312 3068 9364 3120
rect 5632 2932 5684 2984
rect 5724 2975 5776 2984
rect 5724 2941 5733 2975
rect 5733 2941 5767 2975
rect 5767 2941 5776 2975
rect 5724 2932 5776 2941
rect 7196 2932 7248 2984
rect 7564 2932 7616 2984
rect 8944 3000 8996 3052
rect 7932 2975 7984 2984
rect 7932 2941 7941 2975
rect 7941 2941 7975 2975
rect 7975 2941 7984 2975
rect 7932 2932 7984 2941
rect 8300 2932 8352 2984
rect 9864 3000 9916 3052
rect 9588 2975 9640 2984
rect 9588 2941 9597 2975
rect 9597 2941 9631 2975
rect 9631 2941 9640 2975
rect 9588 2932 9640 2941
rect 9680 2932 9732 2984
rect 10324 3000 10376 3052
rect 12256 3136 12308 3188
rect 12440 3179 12492 3188
rect 12440 3145 12449 3179
rect 12449 3145 12483 3179
rect 12483 3145 12492 3179
rect 12440 3136 12492 3145
rect 13084 3136 13136 3188
rect 16212 3136 16264 3188
rect 16764 3136 16816 3188
rect 16948 3136 17000 3188
rect 20352 3136 20404 3188
rect 20444 3179 20496 3188
rect 20444 3145 20453 3179
rect 20453 3145 20487 3179
rect 20487 3145 20496 3179
rect 20444 3136 20496 3145
rect 11428 3068 11480 3120
rect 13176 3068 13228 3120
rect 13728 3068 13780 3120
rect 14004 3000 14056 3052
rect 14464 3000 14516 3052
rect 10968 2975 11020 2984
rect 10968 2941 10977 2975
rect 10977 2941 11011 2975
rect 11011 2941 11020 2975
rect 10968 2932 11020 2941
rect 11520 2932 11572 2984
rect 11612 2932 11664 2984
rect 12164 2975 12216 2984
rect 12164 2941 12173 2975
rect 12173 2941 12207 2975
rect 12207 2941 12216 2975
rect 12164 2932 12216 2941
rect 12256 2975 12308 2984
rect 12256 2941 12289 2975
rect 12289 2941 12308 2975
rect 12256 2932 12308 2941
rect 13728 2932 13780 2984
rect 13912 2975 13964 2984
rect 13912 2941 13921 2975
rect 13921 2941 13955 2975
rect 13955 2941 13964 2975
rect 13912 2932 13964 2941
rect 3700 2864 3752 2916
rect 5540 2907 5592 2916
rect 5540 2873 5549 2907
rect 5549 2873 5583 2907
rect 5583 2873 5592 2907
rect 5540 2864 5592 2873
rect 6644 2864 6696 2916
rect 12808 2864 12860 2916
rect 5172 2839 5224 2848
rect 5172 2805 5181 2839
rect 5181 2805 5215 2839
rect 5215 2805 5224 2839
rect 5172 2796 5224 2805
rect 8116 2796 8168 2848
rect 9680 2796 9732 2848
rect 9864 2839 9916 2848
rect 9864 2805 9873 2839
rect 9873 2805 9907 2839
rect 9907 2805 9916 2839
rect 9864 2796 9916 2805
rect 10508 2796 10560 2848
rect 11612 2796 11664 2848
rect 14188 2864 14240 2916
rect 15844 2975 15896 2984
rect 15844 2941 15853 2975
rect 15853 2941 15887 2975
rect 15887 2941 15896 2975
rect 15844 2932 15896 2941
rect 16580 3000 16632 3052
rect 16488 2975 16540 2984
rect 16488 2941 16497 2975
rect 16497 2941 16531 2975
rect 16531 2941 16540 2975
rect 16488 2932 16540 2941
rect 16764 2975 16816 2984
rect 16764 2941 16773 2975
rect 16773 2941 16807 2975
rect 16807 2941 16816 2975
rect 16764 2932 16816 2941
rect 18144 3000 18196 3052
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 19432 2932 19484 2984
rect 16028 2907 16080 2916
rect 16028 2873 16037 2907
rect 16037 2873 16071 2907
rect 16071 2873 16080 2907
rect 16028 2864 16080 2873
rect 16120 2907 16172 2916
rect 16120 2873 16129 2907
rect 16129 2873 16163 2907
rect 16163 2873 16172 2907
rect 16120 2864 16172 2873
rect 16672 2907 16724 2916
rect 16672 2873 16681 2907
rect 16681 2873 16715 2907
rect 16715 2873 16724 2907
rect 16672 2864 16724 2873
rect 14464 2839 14516 2848
rect 14464 2805 14473 2839
rect 14473 2805 14507 2839
rect 14507 2805 14516 2839
rect 14464 2796 14516 2805
rect 16488 2796 16540 2848
rect 16948 2796 17000 2848
rect 7114 2694 7166 2746
rect 7178 2694 7230 2746
rect 7242 2694 7294 2746
rect 7306 2694 7358 2746
rect 7370 2694 7422 2746
rect 13830 2694 13882 2746
rect 13894 2694 13946 2746
rect 13958 2694 14010 2746
rect 14022 2694 14074 2746
rect 14086 2694 14138 2746
rect 20546 2694 20598 2746
rect 20610 2694 20662 2746
rect 20674 2694 20726 2746
rect 20738 2694 20790 2746
rect 20802 2694 20854 2746
rect 27262 2694 27314 2746
rect 27326 2694 27378 2746
rect 27390 2694 27442 2746
rect 27454 2694 27506 2746
rect 27518 2694 27570 2746
rect 3700 2635 3752 2644
rect 3700 2601 3709 2635
rect 3709 2601 3743 2635
rect 3743 2601 3752 2635
rect 3700 2592 3752 2601
rect 7656 2592 7708 2644
rect 7748 2592 7800 2644
rect 6644 2524 6696 2576
rect 3608 2456 3660 2508
rect 5172 2499 5224 2508
rect 5172 2465 5181 2499
rect 5181 2465 5215 2499
rect 5215 2465 5224 2499
rect 5172 2456 5224 2465
rect 5356 2499 5408 2508
rect 5356 2465 5365 2499
rect 5365 2465 5399 2499
rect 5399 2465 5408 2499
rect 5356 2456 5408 2465
rect 5816 2456 5868 2508
rect 7380 2456 7432 2508
rect 8392 2524 8444 2576
rect 9588 2592 9640 2644
rect 14280 2592 14332 2644
rect 16212 2592 16264 2644
rect 20076 2592 20128 2644
rect 11428 2524 11480 2576
rect 7840 2499 7892 2508
rect 7840 2465 7849 2499
rect 7849 2465 7883 2499
rect 7883 2465 7892 2499
rect 7840 2456 7892 2465
rect 8116 2456 8168 2508
rect 9864 2456 9916 2508
rect 10508 2499 10560 2508
rect 10508 2465 10517 2499
rect 10517 2465 10551 2499
rect 10551 2465 10560 2499
rect 10508 2456 10560 2465
rect 12532 2524 12584 2576
rect 15292 2524 15344 2576
rect 12440 2499 12492 2508
rect 12440 2465 12449 2499
rect 12449 2465 12483 2499
rect 12483 2465 12492 2499
rect 12440 2456 12492 2465
rect 14372 2456 14424 2508
rect 14464 2456 14516 2508
rect 6092 2388 6144 2440
rect 7748 2388 7800 2440
rect 5356 2320 5408 2372
rect 9956 2320 10008 2372
rect 12716 2388 12768 2440
rect 5080 2252 5132 2304
rect 6368 2252 6420 2304
rect 8484 2295 8536 2304
rect 8484 2261 8493 2295
rect 8493 2261 8527 2295
rect 8527 2261 8536 2295
rect 8484 2252 8536 2261
rect 10324 2295 10376 2304
rect 10324 2261 10333 2295
rect 10333 2261 10367 2295
rect 10367 2261 10376 2295
rect 10324 2252 10376 2261
rect 11520 2252 11572 2304
rect 14464 2320 14516 2372
rect 16488 2499 16540 2508
rect 16488 2465 16497 2499
rect 16497 2465 16531 2499
rect 16531 2465 16540 2499
rect 16488 2456 16540 2465
rect 16948 2499 17000 2508
rect 16948 2465 16957 2499
rect 16957 2465 16991 2499
rect 16991 2465 17000 2499
rect 16948 2456 17000 2465
rect 19800 2499 19852 2508
rect 19800 2465 19809 2499
rect 19809 2465 19843 2499
rect 19843 2465 19852 2499
rect 19800 2456 19852 2465
rect 19984 2499 20036 2508
rect 19984 2465 19993 2499
rect 19993 2465 20027 2499
rect 20027 2465 20036 2499
rect 19984 2456 20036 2465
rect 20076 2456 20128 2508
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 21824 2388 21876 2440
rect 21456 2320 21508 2372
rect 14740 2252 14792 2304
rect 16120 2252 16172 2304
rect 17592 2252 17644 2304
rect 17776 2252 17828 2304
rect 3756 2150 3808 2202
rect 3820 2150 3872 2202
rect 3884 2150 3936 2202
rect 3948 2150 4000 2202
rect 4012 2150 4064 2202
rect 10472 2150 10524 2202
rect 10536 2150 10588 2202
rect 10600 2150 10652 2202
rect 10664 2150 10716 2202
rect 10728 2150 10780 2202
rect 17188 2150 17240 2202
rect 17252 2150 17304 2202
rect 17316 2150 17368 2202
rect 17380 2150 17432 2202
rect 17444 2150 17496 2202
rect 23904 2150 23956 2202
rect 23968 2150 24020 2202
rect 24032 2150 24084 2202
rect 24096 2150 24148 2202
rect 24160 2150 24212 2202
rect 6552 2048 6604 2100
rect 7656 2048 7708 2100
rect 8300 2048 8352 2100
rect 9036 2048 9088 2100
rect 9588 2048 9640 2100
rect 5724 1980 5776 2032
rect 6736 1912 6788 1964
rect 7748 1912 7800 1964
rect 4528 1887 4580 1896
rect 4528 1853 4537 1887
rect 4537 1853 4571 1887
rect 4571 1853 4580 1887
rect 4528 1844 4580 1853
rect 5356 1844 5408 1896
rect 6368 1887 6420 1896
rect 6368 1853 6377 1887
rect 6377 1853 6411 1887
rect 6411 1853 6420 1887
rect 6368 1844 6420 1853
rect 7564 1887 7616 1896
rect 7564 1853 7573 1887
rect 7573 1853 7607 1887
rect 7607 1853 7616 1887
rect 7564 1844 7616 1853
rect 15660 2048 15712 2100
rect 13728 1980 13780 2032
rect 4896 1776 4948 1828
rect 4344 1708 4396 1760
rect 6644 1751 6696 1760
rect 6644 1717 6653 1751
rect 6653 1717 6687 1751
rect 6687 1717 6696 1751
rect 6644 1708 6696 1717
rect 8116 1887 8168 1896
rect 8116 1853 8125 1887
rect 8125 1853 8159 1887
rect 8159 1853 8168 1887
rect 8116 1844 8168 1853
rect 9404 1844 9456 1896
rect 8484 1776 8536 1828
rect 12808 1912 12860 1964
rect 10324 1844 10376 1896
rect 11520 1887 11572 1896
rect 11520 1853 11529 1887
rect 11529 1853 11563 1887
rect 11563 1853 11572 1887
rect 11520 1844 11572 1853
rect 12716 1844 12768 1896
rect 16580 1980 16632 2032
rect 9680 1776 9732 1828
rect 12900 1776 12952 1828
rect 10232 1751 10284 1760
rect 10232 1717 10241 1751
rect 10241 1717 10275 1751
rect 10275 1717 10284 1751
rect 10232 1708 10284 1717
rect 11336 1751 11388 1760
rect 11336 1717 11345 1751
rect 11345 1717 11379 1751
rect 11379 1717 11388 1751
rect 11336 1708 11388 1717
rect 12808 1751 12860 1760
rect 12808 1717 12817 1751
rect 12817 1717 12851 1751
rect 12851 1717 12860 1751
rect 12808 1708 12860 1717
rect 14464 1887 14516 1896
rect 14464 1853 14473 1887
rect 14473 1853 14507 1887
rect 14507 1853 14516 1887
rect 14464 1844 14516 1853
rect 19064 1912 19116 1964
rect 20536 1912 20588 1964
rect 15568 1844 15620 1896
rect 15936 1887 15988 1896
rect 15936 1853 15945 1887
rect 15945 1853 15979 1887
rect 15979 1853 15988 1887
rect 15936 1844 15988 1853
rect 16120 1887 16172 1896
rect 16120 1853 16134 1887
rect 16134 1853 16168 1887
rect 16168 1853 16172 1887
rect 16120 1844 16172 1853
rect 17776 1887 17828 1896
rect 17776 1853 17794 1887
rect 17794 1853 17828 1887
rect 17776 1844 17828 1853
rect 18052 1887 18104 1896
rect 18052 1853 18061 1887
rect 18061 1853 18095 1887
rect 18095 1853 18104 1887
rect 18052 1844 18104 1853
rect 18144 1844 18196 1896
rect 13912 1776 13964 1828
rect 16396 1776 16448 1828
rect 19156 1887 19208 1896
rect 19156 1853 19165 1887
rect 19165 1853 19199 1887
rect 19199 1853 19208 1887
rect 19156 1844 19208 1853
rect 19708 1844 19760 1896
rect 20444 1887 20496 1896
rect 20444 1853 20453 1887
rect 20453 1853 20487 1887
rect 20487 1853 20496 1887
rect 20444 1844 20496 1853
rect 20628 1844 20680 1896
rect 19800 1776 19852 1828
rect 27068 1776 27120 1828
rect 14372 1708 14424 1760
rect 15108 1751 15160 1760
rect 15108 1717 15117 1751
rect 15117 1717 15151 1751
rect 15151 1717 15160 1751
rect 15108 1708 15160 1717
rect 15844 1708 15896 1760
rect 17868 1708 17920 1760
rect 25320 1708 25372 1760
rect 7114 1606 7166 1658
rect 7178 1606 7230 1658
rect 7242 1606 7294 1658
rect 7306 1606 7358 1658
rect 7370 1606 7422 1658
rect 13830 1606 13882 1658
rect 13894 1606 13946 1658
rect 13958 1606 14010 1658
rect 14022 1606 14074 1658
rect 14086 1606 14138 1658
rect 20546 1606 20598 1658
rect 20610 1606 20662 1658
rect 20674 1606 20726 1658
rect 20738 1606 20790 1658
rect 20802 1606 20854 1658
rect 27262 1606 27314 1658
rect 27326 1606 27378 1658
rect 27390 1606 27442 1658
rect 27454 1606 27506 1658
rect 27518 1606 27570 1658
rect 4896 1547 4948 1556
rect 4896 1513 4905 1547
rect 4905 1513 4939 1547
rect 4939 1513 4948 1547
rect 4896 1504 4948 1513
rect 7472 1504 7524 1556
rect 9220 1504 9272 1556
rect 9496 1504 9548 1556
rect 848 1436 900 1488
rect 5080 1411 5132 1420
rect 5080 1377 5089 1411
rect 5089 1377 5123 1411
rect 5123 1377 5132 1411
rect 5080 1368 5132 1377
rect 6644 1436 6696 1488
rect 8944 1411 8996 1420
rect 8944 1377 8953 1411
rect 8953 1377 8987 1411
rect 8987 1377 8996 1411
rect 8944 1368 8996 1377
rect 9772 1504 9824 1556
rect 10324 1504 10376 1556
rect 11428 1504 11480 1556
rect 12992 1504 13044 1556
rect 14188 1504 14240 1556
rect 10232 1436 10284 1488
rect 11336 1436 11388 1488
rect 12808 1479 12860 1488
rect 12808 1445 12842 1479
rect 12842 1445 12860 1479
rect 12808 1436 12860 1445
rect 12900 1436 12952 1488
rect 16212 1504 16264 1556
rect 16396 1504 16448 1556
rect 17960 1504 18012 1556
rect 18512 1504 18564 1556
rect 19064 1504 19116 1556
rect 15108 1479 15160 1488
rect 15108 1445 15126 1479
rect 15126 1445 15160 1479
rect 15108 1436 15160 1445
rect 17592 1436 17644 1488
rect 4528 1300 4580 1352
rect 5448 1300 5500 1352
rect 8852 1343 8904 1352
rect 8852 1309 8861 1343
rect 8861 1309 8895 1343
rect 8895 1309 8904 1343
rect 8852 1300 8904 1309
rect 9404 1343 9456 1352
rect 9404 1309 9413 1343
rect 9413 1309 9447 1343
rect 9447 1309 9456 1343
rect 9404 1300 9456 1309
rect 9036 1232 9088 1284
rect 13912 1300 13964 1352
rect 14556 1368 14608 1420
rect 15568 1368 15620 1420
rect 17960 1411 18012 1420
rect 17960 1377 17969 1411
rect 17969 1377 18003 1411
rect 18003 1377 18012 1411
rect 17960 1368 18012 1377
rect 12716 1164 12768 1216
rect 14372 1164 14424 1216
rect 15568 1207 15620 1216
rect 15568 1173 15577 1207
rect 15577 1173 15611 1207
rect 15611 1173 15620 1207
rect 15568 1164 15620 1173
rect 17868 1300 17920 1352
rect 18144 1411 18196 1420
rect 18144 1377 18158 1411
rect 18158 1377 18192 1411
rect 18192 1377 18196 1411
rect 18144 1368 18196 1377
rect 19248 1411 19300 1420
rect 19248 1377 19257 1411
rect 19257 1377 19291 1411
rect 19291 1377 19300 1411
rect 19248 1368 19300 1377
rect 19340 1411 19392 1420
rect 19340 1377 19349 1411
rect 19349 1377 19383 1411
rect 19383 1377 19392 1411
rect 19340 1368 19392 1377
rect 19800 1411 19852 1420
rect 19800 1377 19809 1411
rect 19809 1377 19843 1411
rect 19843 1377 19852 1411
rect 19800 1368 19852 1377
rect 19892 1368 19944 1420
rect 21456 1436 21508 1488
rect 23572 1368 23624 1420
rect 18052 1232 18104 1284
rect 18328 1207 18380 1216
rect 18328 1173 18337 1207
rect 18337 1173 18371 1207
rect 18371 1173 18380 1207
rect 18328 1164 18380 1173
rect 20076 1164 20128 1216
rect 3756 1062 3808 1114
rect 3820 1062 3872 1114
rect 3884 1062 3936 1114
rect 3948 1062 4000 1114
rect 4012 1062 4064 1114
rect 10472 1062 10524 1114
rect 10536 1062 10588 1114
rect 10600 1062 10652 1114
rect 10664 1062 10716 1114
rect 10728 1062 10780 1114
rect 17188 1062 17240 1114
rect 17252 1062 17304 1114
rect 17316 1062 17368 1114
rect 17380 1062 17432 1114
rect 17444 1062 17496 1114
rect 23904 1062 23956 1114
rect 23968 1062 24020 1114
rect 24032 1062 24084 1114
rect 24096 1062 24148 1114
rect 24160 1062 24212 1114
rect 7840 892 7892 944
rect 7748 867 7800 876
rect 7748 833 7757 867
rect 7757 833 7791 867
rect 7791 833 7800 867
rect 9036 892 9088 944
rect 9588 892 9640 944
rect 7748 824 7800 833
rect 7656 799 7708 808
rect 7656 765 7665 799
rect 7665 765 7699 799
rect 7699 765 7708 799
rect 7656 756 7708 765
rect 2596 688 2648 740
rect 7472 688 7524 740
rect 8116 756 8168 808
rect 8852 824 8904 876
rect 8760 799 8812 808
rect 8760 765 8769 799
rect 8769 765 8803 799
rect 8803 765 8812 799
rect 8760 756 8812 765
rect 9036 799 9088 808
rect 9036 765 9045 799
rect 9045 765 9079 799
rect 9079 765 9088 799
rect 10324 824 10376 876
rect 11336 935 11388 944
rect 11336 901 11345 935
rect 11345 901 11379 935
rect 11379 901 11388 935
rect 11336 892 11388 901
rect 12716 892 12768 944
rect 12992 892 13044 944
rect 13084 935 13136 944
rect 13084 901 13093 935
rect 13093 901 13127 935
rect 13127 901 13136 935
rect 13084 892 13136 901
rect 9036 756 9088 765
rect 9220 688 9272 740
rect 9956 688 10008 740
rect 11612 799 11664 808
rect 11612 765 11621 799
rect 11621 765 11655 799
rect 11655 765 11664 799
rect 11612 756 11664 765
rect 11152 688 11204 740
rect 14740 892 14792 944
rect 14832 935 14884 944
rect 14832 901 14841 935
rect 14841 901 14875 935
rect 14875 901 14884 935
rect 14832 892 14884 901
rect 15568 824 15620 876
rect 14372 756 14424 808
rect 14740 799 14792 808
rect 14740 765 14743 799
rect 14743 765 14792 799
rect 14740 756 14792 765
rect 13912 688 13964 740
rect 19708 620 19760 672
rect 7114 518 7166 570
rect 7178 518 7230 570
rect 7242 518 7294 570
rect 7306 518 7358 570
rect 7370 518 7422 570
rect 13830 518 13882 570
rect 13894 518 13946 570
rect 13958 518 14010 570
rect 14022 518 14074 570
rect 14086 518 14138 570
rect 20546 518 20598 570
rect 20610 518 20662 570
rect 20674 518 20726 570
rect 20738 518 20790 570
rect 20802 518 20854 570
rect 27262 518 27314 570
rect 27326 518 27378 570
rect 27390 518 27442 570
rect 27454 518 27506 570
rect 27518 518 27570 570
<< metal2 >>
rect 754 17762 810 18000
rect 1398 17762 1454 18000
rect 754 17734 888 17762
rect 754 17600 810 17734
rect 860 17338 888 17734
rect 1398 17734 1532 17762
rect 1398 17600 1454 17734
rect 1504 17338 1532 17734
rect 2042 17600 2098 18000
rect 2686 17600 2742 18000
rect 3330 17762 3386 18000
rect 3974 17762 4030 18000
rect 3330 17734 3464 17762
rect 3330 17600 3386 17734
rect 848 17332 900 17338
rect 848 17274 900 17280
rect 1492 17332 1544 17338
rect 1492 17274 1544 17280
rect 2056 16522 2084 17600
rect 2700 17202 2728 17600
rect 3436 17202 3464 17734
rect 3620 17734 4030 17762
rect 3620 17338 3648 17734
rect 3974 17600 4030 17734
rect 4618 17762 4674 18000
rect 4618 17734 4752 17762
rect 4618 17600 4674 17734
rect 3756 17436 4064 17445
rect 3756 17434 3762 17436
rect 3818 17434 3842 17436
rect 3898 17434 3922 17436
rect 3978 17434 4002 17436
rect 4058 17434 4064 17436
rect 3818 17382 3820 17434
rect 4000 17382 4002 17434
rect 3756 17380 3762 17382
rect 3818 17380 3842 17382
rect 3898 17380 3922 17382
rect 3978 17380 4002 17382
rect 4058 17380 4064 17382
rect 3756 17371 4064 17380
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 4724 17202 4752 17734
rect 5262 17600 5318 18000
rect 5906 17600 5962 18000
rect 6550 17600 6606 18000
rect 7194 17600 7250 18000
rect 7838 17600 7894 18000
rect 8482 17600 8538 18000
rect 9126 17600 9182 18000
rect 9770 17762 9826 18000
rect 9692 17734 9826 17762
rect 5276 17202 5304 17600
rect 5920 17338 5948 17600
rect 6564 17338 6592 17600
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 7208 17270 7236 17600
rect 7196 17264 7248 17270
rect 7196 17206 7248 17212
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 2044 16516 2096 16522
rect 2044 16458 2096 16464
rect 3756 16348 4064 16357
rect 3756 16346 3762 16348
rect 3818 16346 3842 16348
rect 3898 16346 3922 16348
rect 3978 16346 4002 16348
rect 4058 16346 4064 16348
rect 3818 16294 3820 16346
rect 4000 16294 4002 16346
rect 3756 16292 3762 16294
rect 3818 16292 3842 16294
rect 3898 16292 3922 16294
rect 3978 16292 4002 16294
rect 4058 16292 4064 16294
rect 3756 16283 4064 16292
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 14958 1440 15438
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 14414 1440 14894
rect 3436 14618 3464 15506
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 3756 15260 4064 15269
rect 3756 15258 3762 15260
rect 3818 15258 3842 15260
rect 3898 15258 3922 15260
rect 3978 15258 4002 15260
rect 4058 15258 4064 15260
rect 3818 15206 3820 15258
rect 4000 15206 4002 15258
rect 3756 15204 3762 15206
rect 3818 15204 3842 15206
rect 3898 15204 3922 15206
rect 3978 15204 4002 15206
rect 4058 15204 4064 15206
rect 3756 15195 4064 15204
rect 4264 14958 4292 15302
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3804 14482 3832 14758
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 12782 1440 14350
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 3068 13802 3096 14214
rect 3252 14074 3280 14418
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 3344 13818 3372 13942
rect 3436 13938 3464 14214
rect 3756 14172 4064 14181
rect 3756 14170 3762 14172
rect 3818 14170 3842 14172
rect 3898 14170 3922 14172
rect 3978 14170 4002 14172
rect 4058 14170 4064 14172
rect 3818 14118 3820 14170
rect 4000 14118 4002 14170
rect 3756 14116 3762 14118
rect 3818 14116 3842 14118
rect 3898 14116 3922 14118
rect 3978 14116 4002 14118
rect 4058 14116 4064 14118
rect 3756 14107 4064 14116
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3516 13864 3568 13870
rect 3056 13796 3108 13802
rect 3344 13790 3464 13818
rect 3516 13806 3568 13812
rect 3056 13738 3108 13744
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 12374 1440 12718
rect 1400 12368 1452 12374
rect 1400 12310 1452 12316
rect 2056 12306 2084 13126
rect 3068 12782 3096 13738
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2700 11218 2728 12378
rect 3068 11694 3096 12718
rect 3160 12102 3188 12718
rect 3252 12238 3280 13262
rect 3436 12646 3464 13790
rect 3528 13462 3556 13806
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 3606 13560 3662 13569
rect 3606 13495 3662 13504
rect 3516 13456 3568 13462
rect 3516 13398 3568 13404
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3344 12306 3372 12582
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3436 12238 3464 12582
rect 3620 12374 3648 13495
rect 3790 13424 3846 13433
rect 3790 13359 3792 13368
rect 3844 13359 3846 13368
rect 3792 13330 3844 13336
rect 4080 13326 4108 13670
rect 4172 13530 4200 14418
rect 4264 13870 4292 14894
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 4356 14618 4384 14826
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4344 14000 4396 14006
rect 4344 13942 4396 13948
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4356 13569 4384 13942
rect 4342 13560 4398 13569
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4252 13524 4304 13530
rect 4342 13495 4398 13504
rect 4252 13466 4304 13472
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 3756 13084 4064 13093
rect 3756 13082 3762 13084
rect 3818 13082 3842 13084
rect 3898 13082 3922 13084
rect 3978 13082 4002 13084
rect 4058 13082 4064 13084
rect 3818 13030 3820 13082
rect 4000 13030 4002 13082
rect 3756 13028 3762 13030
rect 3818 13028 3842 13030
rect 3898 13028 3922 13030
rect 3978 13028 4002 13030
rect 4058 13028 4064 13030
rect 3756 13019 4064 13028
rect 4172 12986 4200 13194
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 3804 12238 3832 12786
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2700 10130 2728 11154
rect 3160 10606 3188 12038
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2884 9722 2912 10066
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1596 8430 1624 8910
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1596 6866 1624 8366
rect 2596 8356 2648 8362
rect 2596 8298 2648 8304
rect 2608 8090 2636 8298
rect 2792 8090 2820 8434
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2792 7954 2820 8026
rect 2976 7954 3004 9318
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3160 7954 3188 8298
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3252 7478 3280 9386
rect 3344 8566 3372 9454
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3332 7880 3384 7886
rect 3436 7868 3464 12174
rect 4080 12170 4108 12650
rect 4172 12374 4200 12922
rect 4264 12850 4292 13466
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 4356 13258 4384 13330
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4356 12374 4384 13194
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4344 12368 4396 12374
rect 4344 12310 4396 12316
rect 4448 12170 4476 14010
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4540 13802 4568 13874
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4526 13424 4582 13433
rect 4526 13359 4582 13368
rect 4540 12306 4568 13359
rect 4632 12850 4660 16594
rect 5276 15162 5304 16594
rect 5920 16522 5948 17070
rect 6000 17060 6052 17066
rect 6000 17002 6052 17008
rect 5908 16516 5960 16522
rect 5908 16458 5960 16464
rect 5920 16250 5948 16458
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5908 15972 5960 15978
rect 5908 15914 5960 15920
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 4816 14482 4844 15098
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 5092 13938 5120 14826
rect 5368 14618 5396 14894
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5276 14498 5304 14554
rect 5552 14550 5580 14894
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5540 14544 5592 14550
rect 5276 14470 5396 14498
rect 5540 14486 5592 14492
rect 5368 14414 5396 14470
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5276 13530 5304 13806
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 4436 12164 4488 12170
rect 4436 12106 4488 12112
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11898 3648 12038
rect 3756 11996 4064 12005
rect 3756 11994 3762 11996
rect 3818 11994 3842 11996
rect 3898 11994 3922 11996
rect 3978 11994 4002 11996
rect 4058 11994 4064 11996
rect 3818 11942 3820 11994
rect 4000 11942 4002 11994
rect 3756 11940 3762 11942
rect 3818 11940 3842 11942
rect 3898 11940 3922 11942
rect 3978 11940 4002 11942
rect 4058 11940 4064 11942
rect 3756 11931 4064 11940
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 4724 11694 4752 13466
rect 4804 13456 4856 13462
rect 4802 13424 4804 13433
rect 4856 13424 4858 13433
rect 4802 13359 4858 13368
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4816 12442 4844 12718
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4816 12170 4844 12242
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4816 11762 4844 12106
rect 4908 11898 4936 12650
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4816 11506 4844 11698
rect 4724 11478 4844 11506
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4448 11218 4476 11290
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 3756 10908 4064 10917
rect 3756 10906 3762 10908
rect 3818 10906 3842 10908
rect 3898 10906 3922 10908
rect 3978 10906 4002 10908
rect 4058 10906 4064 10908
rect 3818 10854 3820 10906
rect 4000 10854 4002 10906
rect 3756 10852 3762 10854
rect 3818 10852 3842 10854
rect 3898 10852 3922 10854
rect 3978 10852 4002 10854
rect 4058 10852 4064 10854
rect 3756 10843 4064 10852
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 4068 10124 4120 10130
rect 4172 10112 4200 10474
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4120 10084 4200 10112
rect 4068 10066 4120 10072
rect 4356 10062 4384 10406
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 3756 9820 4064 9829
rect 3756 9818 3762 9820
rect 3818 9818 3842 9820
rect 3898 9818 3922 9820
rect 3978 9818 4002 9820
rect 4058 9818 4064 9820
rect 3818 9766 3820 9818
rect 4000 9766 4002 9818
rect 3756 9764 3762 9766
rect 3818 9764 3842 9766
rect 3898 9764 3922 9766
rect 3978 9764 4002 9766
rect 4058 9764 4064 9766
rect 3756 9755 4064 9764
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3620 8634 3648 8978
rect 3756 8732 4064 8741
rect 3756 8730 3762 8732
rect 3818 8730 3842 8732
rect 3898 8730 3922 8732
rect 3978 8730 4002 8732
rect 4058 8730 4064 8732
rect 3818 8678 3820 8730
rect 4000 8678 4002 8730
rect 3756 8676 3762 8678
rect 3818 8676 3842 8678
rect 3898 8676 3922 8678
rect 3978 8676 4002 8678
rect 4058 8676 4064 8678
rect 3756 8667 4064 8676
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3528 7954 3556 8230
rect 3896 7954 3924 8502
rect 4172 8430 4200 9590
rect 4264 9518 4292 9862
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 3384 7840 3464 7868
rect 3332 7822 3384 7828
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 3344 7206 3372 7822
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3436 7274 3464 7686
rect 3620 7562 3648 7890
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 3756 7644 4064 7653
rect 3756 7642 3762 7644
rect 3818 7642 3842 7644
rect 3898 7642 3922 7644
rect 3978 7642 4002 7644
rect 4058 7642 4064 7644
rect 3818 7590 3820 7642
rect 4000 7590 4002 7642
rect 3756 7588 3762 7590
rect 3818 7588 3842 7590
rect 3898 7588 3922 7590
rect 3978 7588 4002 7590
rect 4058 7588 4064 7590
rect 3756 7579 4064 7588
rect 3528 7534 3648 7562
rect 3528 7342 3556 7534
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3804 7342 3832 7414
rect 4172 7410 4200 7686
rect 4264 7546 4292 7890
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 2792 6866 2820 7142
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 3528 6254 3556 7278
rect 3712 7002 3740 7278
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 3756 6556 4064 6565
rect 3756 6554 3762 6556
rect 3818 6554 3842 6556
rect 3898 6554 3922 6556
rect 3978 6554 4002 6556
rect 4058 6554 4064 6556
rect 3818 6502 3820 6554
rect 4000 6502 4002 6554
rect 3756 6500 3762 6502
rect 3818 6500 3842 6502
rect 3898 6500 3922 6502
rect 3978 6500 4002 6502
rect 4058 6500 4064 6502
rect 3756 6491 4064 6500
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3344 4690 3372 5510
rect 3756 5468 4064 5477
rect 3756 5466 3762 5468
rect 3818 5466 3842 5468
rect 3898 5466 3922 5468
rect 3978 5466 4002 5468
rect 4058 5466 4064 5468
rect 3818 5414 3820 5466
rect 4000 5414 4002 5466
rect 3756 5412 3762 5414
rect 3818 5412 3842 5414
rect 3898 5412 3922 5414
rect 3978 5412 4002 5414
rect 4058 5412 4064 5414
rect 3756 5403 4064 5412
rect 4172 5234 4200 6802
rect 4264 5778 4292 7142
rect 4356 5914 4384 9862
rect 4448 9450 4476 11154
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4632 10266 4660 10542
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4448 9081 4476 9386
rect 4434 9072 4490 9081
rect 4434 9007 4490 9016
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 8498 4476 8774
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4632 7002 4660 7278
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4632 6186 4660 6938
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4172 4758 4200 5170
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3756 4380 4064 4389
rect 3756 4378 3762 4380
rect 3818 4378 3842 4380
rect 3898 4378 3922 4380
rect 3978 4378 4002 4380
rect 4058 4378 4064 4380
rect 3818 4326 3820 4378
rect 4000 4326 4002 4378
rect 3756 4324 3762 4326
rect 3818 4324 3842 4326
rect 3898 4324 3922 4326
rect 3978 4324 4002 4326
rect 4058 4324 4064 4326
rect 3756 4315 4064 4324
rect 4172 4146 4200 4694
rect 4356 4622 4384 5850
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4540 4826 4568 5646
rect 4724 5522 4752 11478
rect 5000 11354 5028 13126
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 5184 11218 5212 12310
rect 5368 12170 5396 14350
rect 5828 14074 5856 14758
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5644 13462 5672 13806
rect 5632 13456 5684 13462
rect 5828 13433 5856 14010
rect 5632 13398 5684 13404
rect 5814 13424 5870 13433
rect 5814 13359 5870 13368
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 5828 12434 5856 13194
rect 5644 12406 5856 12434
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 5368 11694 5396 12106
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5172 11212 5224 11218
rect 5356 11212 5408 11218
rect 5172 11154 5224 11160
rect 5276 11172 5356 11200
rect 5000 10674 5028 11154
rect 5184 11014 5212 11154
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4816 10062 4844 10474
rect 5000 10130 5028 10610
rect 5184 10554 5212 10950
rect 5092 10538 5212 10554
rect 5080 10532 5212 10538
rect 5132 10526 5212 10532
rect 5080 10474 5132 10480
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4816 9518 4844 9998
rect 5092 9518 5120 10474
rect 5276 10266 5304 11172
rect 5356 11154 5408 11160
rect 5460 11200 5488 12174
rect 5644 12102 5672 12406
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5540 11212 5592 11218
rect 5460 11172 5540 11200
rect 5460 10470 5488 11172
rect 5540 11154 5592 11160
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5276 10130 5304 10202
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5368 9602 5396 10406
rect 5460 10266 5488 10406
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5552 9654 5580 10950
rect 5276 9574 5396 9602
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4908 8498 4936 8910
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 5000 8430 5028 9386
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5000 6458 5028 7278
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 5000 5692 5028 6394
rect 5276 6118 5304 9574
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5276 5778 5304 6054
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5080 5704 5132 5710
rect 5000 5664 5080 5692
rect 5080 5646 5132 5652
rect 5184 5658 5212 5714
rect 5184 5630 5304 5658
rect 5368 5642 5396 9454
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5460 7886 5488 8366
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5644 7546 5672 12038
rect 5920 11898 5948 15914
rect 6012 15638 6040 17002
rect 7114 16892 7422 16901
rect 7114 16890 7120 16892
rect 7176 16890 7200 16892
rect 7256 16890 7280 16892
rect 7336 16890 7360 16892
rect 7416 16890 7422 16892
rect 7176 16838 7178 16890
rect 7358 16838 7360 16890
rect 7114 16836 7120 16838
rect 7176 16836 7200 16838
rect 7256 16836 7280 16838
rect 7336 16836 7360 16838
rect 7416 16836 7422 16838
rect 7114 16827 7422 16836
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 6380 16250 6408 16594
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6656 15706 6684 15982
rect 6840 15706 6868 15982
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6000 15632 6052 15638
rect 6000 15574 6052 15580
rect 6012 15162 6040 15574
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6656 15366 6684 15506
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6840 14958 6868 15438
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6472 14618 6500 14758
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 6012 13870 6040 14486
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6288 13870 6316 14418
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6288 13530 6316 13806
rect 6656 13734 6684 14894
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6288 13190 6316 13330
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6564 12782 6592 13398
rect 6748 13394 6776 14758
rect 6840 14550 6868 14894
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 7024 14414 7052 15982
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7114 15804 7422 15813
rect 7114 15802 7120 15804
rect 7176 15802 7200 15804
rect 7256 15802 7280 15804
rect 7336 15802 7360 15804
rect 7416 15802 7422 15804
rect 7176 15750 7178 15802
rect 7358 15750 7360 15802
rect 7114 15748 7120 15750
rect 7176 15748 7200 15750
rect 7256 15748 7280 15750
rect 7336 15748 7360 15750
rect 7416 15748 7422 15750
rect 7114 15739 7422 15748
rect 7380 15564 7432 15570
rect 7484 15552 7512 15846
rect 7432 15524 7512 15552
rect 7380 15506 7432 15512
rect 7114 14716 7422 14725
rect 7114 14714 7120 14716
rect 7176 14714 7200 14716
rect 7256 14714 7280 14716
rect 7336 14714 7360 14716
rect 7416 14714 7422 14716
rect 7176 14662 7178 14714
rect 7358 14662 7360 14714
rect 7114 14660 7120 14662
rect 7176 14660 7200 14662
rect 7256 14660 7280 14662
rect 7336 14660 7360 14662
rect 7416 14660 7422 14662
rect 7114 14651 7422 14660
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7484 13938 7512 14350
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7114 13628 7422 13637
rect 7114 13626 7120 13628
rect 7176 13626 7200 13628
rect 7256 13626 7280 13628
rect 7336 13626 7360 13628
rect 7416 13626 7422 13628
rect 7176 13574 7178 13626
rect 7358 13574 7360 13626
rect 7114 13572 7120 13574
rect 7176 13572 7200 13574
rect 7256 13572 7280 13574
rect 7336 13572 7360 13574
rect 7416 13572 7422 13574
rect 7114 13563 7422 13572
rect 7576 13394 7604 14486
rect 7760 13938 7788 16594
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 6748 12918 6776 13330
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 7024 12850 7052 13262
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6564 12084 6592 12718
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6642 12336 6698 12345
rect 6642 12271 6644 12280
rect 6696 12271 6698 12280
rect 6644 12242 6696 12248
rect 6644 12096 6696 12102
rect 6564 12056 6644 12084
rect 6644 12038 6696 12044
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 6656 11694 6684 12038
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6012 11218 6040 11630
rect 6932 11218 6960 12378
rect 7024 11762 7052 12786
rect 7484 12782 7512 12922
rect 7576 12889 7604 13330
rect 7562 12880 7618 12889
rect 7562 12815 7618 12824
rect 7576 12782 7604 12815
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7114 12540 7422 12549
rect 7114 12538 7120 12540
rect 7176 12538 7200 12540
rect 7256 12538 7280 12540
rect 7336 12538 7360 12540
rect 7416 12538 7422 12540
rect 7176 12486 7178 12538
rect 7358 12486 7360 12538
rect 7114 12484 7120 12486
rect 7176 12484 7200 12486
rect 7256 12484 7280 12486
rect 7336 12484 7360 12486
rect 7416 12484 7422 12486
rect 7114 12475 7422 12484
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7114 11452 7422 11461
rect 7114 11450 7120 11452
rect 7176 11450 7200 11452
rect 7256 11450 7280 11452
rect 7336 11450 7360 11452
rect 7416 11450 7422 11452
rect 7176 11398 7178 11450
rect 7358 11398 7360 11450
rect 7114 11396 7120 11398
rect 7176 11396 7200 11398
rect 7256 11396 7280 11398
rect 7336 11396 7360 11398
rect 7416 11396 7422 11398
rect 7114 11387 7422 11396
rect 7484 11336 7512 12582
rect 7760 12442 7788 13874
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7484 11308 7696 11336
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 5736 9654 5764 11154
rect 6012 10606 6040 11154
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5736 7392 5764 9590
rect 5828 9586 5856 9862
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 6840 9518 6868 10542
rect 6932 10062 6960 11154
rect 7484 10674 7512 11308
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 5736 7364 5948 7392
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5460 5778 5488 6394
rect 5552 6390 5580 6598
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 4724 5494 5028 5522
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4724 4826 4752 5034
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4540 4146 4568 4762
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4632 4134 4844 4162
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2792 3738 2820 3946
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 3436 3602 3464 3878
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3804 3534 3832 4014
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3988 3602 4016 3878
rect 4080 3738 4108 4014
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4172 3670 4200 4082
rect 4632 4078 4660 4134
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4724 3738 4752 4014
rect 4816 3738 4844 4134
rect 5000 4010 5028 5494
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5184 4690 5212 5170
rect 5276 4690 5304 5630
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5540 5568 5592 5574
rect 5644 5522 5672 7278
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5736 5914 5764 6802
rect 5828 6458 5856 7210
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5592 5516 5764 5522
rect 5540 5510 5764 5516
rect 5552 5494 5764 5510
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5552 4282 5580 4966
rect 5644 4758 5672 4966
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3620 2514 3648 3334
rect 3756 3292 4064 3301
rect 3756 3290 3762 3292
rect 3818 3290 3842 3292
rect 3898 3290 3922 3292
rect 3978 3290 4002 3292
rect 4058 3290 4064 3292
rect 3818 3238 3820 3290
rect 4000 3238 4002 3290
rect 3756 3236 3762 3238
rect 3818 3236 3842 3238
rect 3898 3236 3922 3238
rect 3978 3236 4002 3238
rect 4058 3236 4064 3238
rect 3756 3227 4064 3236
rect 4172 3194 4200 3606
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4724 3126 4752 3674
rect 5092 3641 5120 4014
rect 5264 3936 5316 3942
rect 5316 3896 5396 3924
rect 5264 3878 5316 3884
rect 5078 3632 5134 3641
rect 5078 3567 5134 3576
rect 5092 3194 5120 3567
rect 5368 3398 5396 3896
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 3700 2916 3752 2922
rect 3700 2858 3752 2864
rect 3712 2650 3740 2858
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 5184 2514 5212 2790
rect 5368 2514 5396 3334
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5368 2378 5396 2450
rect 5356 2372 5408 2378
rect 5356 2314 5408 2320
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 3756 2204 4064 2213
rect 3756 2202 3762 2204
rect 3818 2202 3842 2204
rect 3898 2202 3922 2204
rect 3978 2202 4002 2204
rect 4058 2202 4064 2204
rect 3818 2150 3820 2202
rect 4000 2150 4002 2202
rect 3756 2148 3762 2150
rect 3818 2148 3842 2150
rect 3898 2148 3922 2150
rect 3978 2148 4002 2150
rect 4058 2148 4064 2150
rect 3756 2139 4064 2148
rect 4528 1896 4580 1902
rect 4528 1838 4580 1844
rect 4344 1760 4396 1766
rect 4344 1702 4396 1708
rect 848 1488 900 1494
rect 848 1430 900 1436
rect 860 400 888 1430
rect 3756 1116 4064 1125
rect 3756 1114 3762 1116
rect 3818 1114 3842 1116
rect 3898 1114 3922 1116
rect 3978 1114 4002 1116
rect 4058 1114 4064 1116
rect 3818 1062 3820 1114
rect 4000 1062 4002 1114
rect 3756 1060 3762 1062
rect 3818 1060 3842 1062
rect 3898 1060 3922 1062
rect 3978 1060 4002 1062
rect 4058 1060 4064 1062
rect 3756 1051 4064 1060
rect 2596 740 2648 746
rect 2596 682 2648 688
rect 2608 400 2636 682
rect 4356 400 4384 1702
rect 4540 1358 4568 1838
rect 4896 1828 4948 1834
rect 4896 1770 4948 1776
rect 4908 1562 4936 1770
rect 4896 1556 4948 1562
rect 4896 1498 4948 1504
rect 5092 1426 5120 2246
rect 5368 1902 5396 2314
rect 5356 1896 5408 1902
rect 5356 1838 5408 1844
rect 5080 1420 5132 1426
rect 5080 1362 5132 1368
rect 5460 1358 5488 3606
rect 5552 2922 5580 4082
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5644 2990 5672 3334
rect 5736 3126 5764 5494
rect 5920 4146 5948 7364
rect 6104 7342 6132 8230
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6012 5778 6040 7142
rect 6104 7002 6132 7142
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6196 6934 6224 7822
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 6196 6390 6224 6870
rect 6288 6746 6316 9318
rect 6380 9110 6408 9454
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6472 7546 6500 7890
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6288 6718 6408 6746
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6184 6384 6236 6390
rect 6184 6326 6236 6332
rect 6288 6322 6316 6598
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 6380 5166 6408 6718
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6380 3670 6408 3878
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5828 3194 5856 3538
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5724 3120 5776 3126
rect 5776 3068 5856 3074
rect 5724 3062 5856 3068
rect 5736 3046 5856 3062
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5736 2038 5764 2926
rect 5828 2514 5856 3046
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 5724 2032 5776 2038
rect 5724 1974 5776 1980
rect 4528 1352 4580 1358
rect 4528 1294 4580 1300
rect 5448 1352 5500 1358
rect 5448 1294 5500 1300
rect 6104 400 6132 2382
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 6380 1902 6408 2246
rect 6564 2106 6592 9386
rect 6656 9042 6684 9454
rect 6840 9160 6868 9454
rect 6748 9132 6868 9160
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6748 7342 6776 9132
rect 6932 9110 6960 9862
rect 7024 9722 7052 10542
rect 7114 10364 7422 10373
rect 7114 10362 7120 10364
rect 7176 10362 7200 10364
rect 7256 10362 7280 10364
rect 7336 10362 7360 10364
rect 7416 10362 7422 10364
rect 7176 10310 7178 10362
rect 7358 10310 7360 10362
rect 7114 10308 7120 10310
rect 7176 10308 7200 10310
rect 7256 10308 7280 10310
rect 7336 10308 7360 10310
rect 7416 10308 7422 10310
rect 7114 10299 7422 10308
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 7392 9466 7420 9522
rect 7484 9466 7512 10610
rect 7576 10470 7604 11154
rect 7668 11014 7696 11308
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7852 10810 7880 17600
rect 8496 17202 8524 17600
rect 9140 17338 9168 17600
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 8036 16114 8064 16390
rect 8496 16250 8524 16594
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8482 15600 8538 15609
rect 8312 14890 8340 15574
rect 8482 15535 8484 15544
rect 8536 15535 8538 15544
rect 8484 15506 8536 15512
rect 8208 14884 8260 14890
rect 8208 14826 8260 14832
rect 8300 14884 8352 14890
rect 8300 14826 8352 14832
rect 8220 14278 8248 14826
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8220 14074 8248 14214
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7944 12646 7972 13262
rect 8220 13190 8248 13738
rect 8312 13326 8340 14826
rect 8588 14822 8616 16594
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9508 16046 9536 16390
rect 9692 16182 9720 17734
rect 9770 17600 9826 17734
rect 10414 17600 10470 18000
rect 11058 17600 11114 18000
rect 11702 17600 11758 18000
rect 12346 17600 12402 18000
rect 12990 17600 13046 18000
rect 13634 17600 13690 18000
rect 14278 17600 14334 18000
rect 14922 17600 14978 18000
rect 15566 17600 15622 18000
rect 16210 17600 16266 18000
rect 16854 17600 16910 18000
rect 17498 17600 17554 18000
rect 18142 17600 18198 18000
rect 18786 17600 18842 18000
rect 19430 17600 19486 18000
rect 20074 17600 20130 18000
rect 20718 17600 20774 18000
rect 21362 17762 21418 18000
rect 21362 17734 21680 17762
rect 21362 17600 21418 17734
rect 10428 17524 10456 17600
rect 10336 17496 10456 17524
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9784 16726 9812 16934
rect 9772 16720 9824 16726
rect 9772 16662 9824 16668
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9772 16108 9824 16114
rect 9876 16096 9904 17138
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10152 16794 10180 17070
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 9824 16068 9904 16096
rect 9772 16050 9824 16056
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 9496 16040 9548 16046
rect 9784 16017 9812 16050
rect 10152 16046 10180 16730
rect 10244 16250 10272 17070
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10140 16040 10192 16046
rect 9496 15982 9548 15988
rect 9770 16008 9826 16017
rect 8864 15706 8892 15982
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8404 13462 8432 14214
rect 8496 13530 8524 14486
rect 8588 14482 8616 14758
rect 8852 14544 8904 14550
rect 8852 14486 8904 14492
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8680 13530 8708 13806
rect 8772 13734 8800 14214
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8864 13530 8892 14486
rect 8956 14278 8984 15302
rect 9324 15162 9352 15506
rect 9508 15502 9536 15982
rect 10140 15982 10192 15988
rect 9770 15943 9826 15952
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9496 15496 9548 15502
rect 9496 15438 9548 15444
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 9508 14958 9536 15438
rect 9692 15434 9720 15506
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9692 15162 9720 15370
rect 9784 15366 9812 15506
rect 9864 15428 9916 15434
rect 9864 15370 9916 15376
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8850 13424 8906 13433
rect 8576 13388 8628 13394
rect 8496 13348 8576 13376
rect 8300 13320 8352 13326
rect 8496 13308 8524 13348
rect 8956 13410 8984 14214
rect 8906 13382 8984 13410
rect 8850 13359 8852 13368
rect 8576 13330 8628 13336
rect 8904 13359 8906 13368
rect 8852 13330 8904 13336
rect 8352 13280 8524 13308
rect 8760 13320 8812 13326
rect 8300 13262 8352 13268
rect 8760 13262 8812 13268
rect 9140 13274 9168 14758
rect 9232 13394 9260 14758
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9416 13818 9444 13874
rect 9600 13870 9628 14758
rect 9876 14618 9904 15370
rect 10336 15094 10364 17496
rect 10472 17436 10780 17445
rect 10472 17434 10478 17436
rect 10534 17434 10558 17436
rect 10614 17434 10638 17436
rect 10694 17434 10718 17436
rect 10774 17434 10780 17436
rect 10534 17382 10536 17434
rect 10716 17382 10718 17434
rect 10472 17380 10478 17382
rect 10534 17380 10558 17382
rect 10614 17380 10638 17382
rect 10694 17380 10718 17382
rect 10774 17380 10780 17382
rect 10472 17371 10780 17380
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10704 16522 10732 17070
rect 11072 16658 11100 17600
rect 11716 16794 11744 17600
rect 12360 16794 12388 17600
rect 13004 17338 13032 17600
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 13648 17270 13676 17600
rect 14292 17338 14320 17600
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14936 17270 14964 17600
rect 15580 17338 15608 17600
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 13636 17264 13688 17270
rect 13636 17206 13688 17212
rect 14924 17264 14976 17270
rect 14924 17206 14976 17212
rect 16224 17134 16252 17600
rect 16580 17264 16632 17270
rect 16580 17206 16632 17212
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 12438 16688 12494 16697
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10692 16516 10744 16522
rect 10692 16458 10744 16464
rect 10472 16348 10780 16357
rect 10472 16346 10478 16348
rect 10534 16346 10558 16348
rect 10614 16346 10638 16348
rect 10694 16346 10718 16348
rect 10774 16346 10780 16348
rect 10534 16294 10536 16346
rect 10716 16294 10718 16346
rect 10472 16292 10478 16294
rect 10534 16292 10558 16294
rect 10614 16292 10638 16294
rect 10694 16292 10718 16294
rect 10774 16292 10780 16294
rect 10472 16283 10780 16292
rect 10888 16250 10916 16594
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10520 15706 10548 15846
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10508 15564 10560 15570
rect 10612 15552 10640 15982
rect 10704 15570 10732 16050
rect 10888 16046 10916 16186
rect 10980 16182 11008 16458
rect 11164 16250 11192 16662
rect 11888 16652 11940 16658
rect 11716 16612 11888 16640
rect 11244 16516 11296 16522
rect 11244 16458 11296 16464
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 10980 16046 11008 16118
rect 11256 16046 11284 16458
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11060 15972 11112 15978
rect 11060 15914 11112 15920
rect 10560 15524 10640 15552
rect 10692 15564 10744 15570
rect 10508 15506 10560 15512
rect 10744 15524 10916 15552
rect 10692 15506 10744 15512
rect 10472 15260 10780 15269
rect 10472 15258 10478 15260
rect 10534 15258 10558 15260
rect 10614 15258 10638 15260
rect 10694 15258 10718 15260
rect 10774 15258 10780 15260
rect 10534 15206 10536 15258
rect 10716 15206 10718 15258
rect 10472 15204 10478 15206
rect 10534 15204 10558 15206
rect 10614 15204 10638 15206
rect 10694 15204 10718 15206
rect 10774 15204 10780 15206
rect 10472 15195 10780 15204
rect 10888 15162 10916 15524
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10324 15088 10376 15094
rect 10324 15030 10376 15036
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9968 14618 9996 14894
rect 10324 14884 10376 14890
rect 10324 14826 10376 14832
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10048 14544 10100 14550
rect 9876 14492 10048 14498
rect 9876 14486 10100 14492
rect 9876 14482 10088 14486
rect 9864 14476 10088 14482
rect 9916 14470 10088 14476
rect 9864 14418 9916 14424
rect 9324 13790 9444 13818
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9324 13274 9352 13790
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9416 13394 9444 13670
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 8036 12442 8064 13126
rect 8220 12782 8248 13126
rect 8772 12782 8800 13262
rect 9140 13246 9352 13274
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 8036 10742 8064 12378
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8588 12102 8616 12242
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8496 11626 8524 12038
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8404 11354 8432 11562
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 8312 10606 8340 11154
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 9722 7604 10066
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 8312 9518 8340 10406
rect 8404 9518 8432 11290
rect 8680 11218 8708 12718
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 7024 9178 7052 9454
rect 7392 9438 7512 9466
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 7114 9276 7422 9285
rect 7114 9274 7120 9276
rect 7176 9274 7200 9276
rect 7256 9274 7280 9276
rect 7336 9274 7360 9276
rect 7416 9274 7422 9276
rect 7176 9222 7178 9274
rect 7358 9222 7360 9274
rect 7114 9220 7120 9222
rect 7176 9220 7200 9222
rect 7256 9220 7280 9222
rect 7336 9220 7360 9222
rect 7416 9220 7422 9222
rect 7114 9211 7422 9220
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 7288 9036 7340 9042
rect 7484 9024 7512 9438
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7576 9042 7604 9318
rect 7340 8996 7512 9024
rect 7564 9036 7616 9042
rect 7288 8978 7340 8984
rect 7564 8978 7616 8984
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8484 9036 8536 9042
rect 8588 9024 8616 10610
rect 8772 10606 8800 12718
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 8864 12374 8892 12582
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8956 12306 8984 12582
rect 9048 12306 9076 12582
rect 9232 12306 9260 12650
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9048 11558 9076 12038
rect 9324 11694 9352 13246
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9416 12986 9444 13194
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9508 12782 9536 13670
rect 9600 13462 9628 13806
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9876 13394 9904 14418
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10244 13394 10272 14214
rect 10336 13870 10364 14826
rect 11072 14618 11100 15914
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 10472 14172 10780 14181
rect 10472 14170 10478 14172
rect 10534 14170 10558 14172
rect 10614 14170 10638 14172
rect 10694 14170 10718 14172
rect 10774 14170 10780 14172
rect 10534 14118 10536 14170
rect 10716 14118 10718 14170
rect 10472 14116 10478 14118
rect 10534 14116 10558 14118
rect 10614 14116 10638 14118
rect 10694 14116 10718 14118
rect 10774 14116 10780 14118
rect 10472 14107 10780 14116
rect 11348 14074 11376 14350
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 9864 13388 9916 13394
rect 9692 13348 9864 13376
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9508 12306 9536 12718
rect 9692 12306 9720 13348
rect 9864 13330 9916 13336
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9416 11812 9444 12038
rect 9588 11824 9640 11830
rect 9416 11784 9588 11812
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8680 10266 8708 10542
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8772 9602 8800 10542
rect 9140 10130 9168 11630
rect 9416 10674 9444 11784
rect 9588 11766 9640 11772
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9600 10606 9628 11494
rect 9784 11370 9812 13126
rect 10244 12782 10272 13330
rect 10336 12782 10364 13806
rect 10966 13424 11022 13433
rect 10966 13359 11022 13368
rect 10472 13084 10780 13093
rect 10472 13082 10478 13084
rect 10534 13082 10558 13084
rect 10614 13082 10638 13084
rect 10694 13082 10718 13084
rect 10774 13082 10780 13084
rect 10534 13030 10536 13082
rect 10716 13030 10718 13082
rect 10472 13028 10478 13030
rect 10534 13028 10558 13030
rect 10614 13028 10638 13030
rect 10694 13028 10718 13030
rect 10774 13028 10780 13030
rect 10472 13019 10780 13028
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 9876 12306 9904 12718
rect 10152 12434 10180 12718
rect 9968 12406 10180 12434
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9968 12238 9996 12406
rect 10704 12238 10732 12718
rect 10980 12714 11008 13359
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10244 11898 10272 12174
rect 10472 11996 10780 12005
rect 10472 11994 10478 11996
rect 10534 11994 10558 11996
rect 10614 11994 10638 11996
rect 10694 11994 10718 11996
rect 10774 11994 10780 11996
rect 10534 11942 10536 11994
rect 10716 11942 10718 11994
rect 10472 11940 10478 11942
rect 10534 11940 10558 11942
rect 10614 11940 10638 11942
rect 10694 11940 10718 11942
rect 10774 11940 10780 11942
rect 10472 11931 10780 11940
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 9968 11778 9996 11834
rect 9968 11750 10180 11778
rect 10046 11656 10102 11665
rect 9864 11620 9916 11626
rect 10152 11626 10180 11750
rect 10046 11591 10102 11600
rect 10140 11620 10192 11626
rect 9864 11562 9916 11568
rect 9692 11342 9812 11370
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9232 9908 9260 10406
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 8680 9574 8800 9602
rect 9140 9880 9260 9908
rect 8680 9042 8708 9574
rect 9140 9518 9168 9880
rect 9416 9722 9444 10066
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 8536 8996 8616 9024
rect 8484 8978 8536 8984
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6748 5370 6776 5782
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6748 4078 6776 4558
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6748 3194 6776 4014
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6748 3058 6776 3130
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 6656 2582 6684 2858
rect 6840 2774 6868 8978
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8430 6960 8774
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 7300 8294 7328 8978
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7114 8188 7422 8197
rect 7114 8186 7120 8188
rect 7176 8186 7200 8188
rect 7256 8186 7280 8188
rect 7336 8186 7360 8188
rect 7416 8186 7422 8188
rect 7176 8134 7178 8186
rect 7358 8134 7360 8186
rect 7114 8132 7120 8134
rect 7176 8132 7200 8134
rect 7256 8132 7280 8134
rect 7336 8132 7360 8134
rect 7416 8132 7422 8134
rect 7114 8123 7422 8132
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7024 6730 7052 7142
rect 7114 7100 7422 7109
rect 7114 7098 7120 7100
rect 7176 7098 7200 7100
rect 7256 7098 7280 7100
rect 7336 7098 7360 7100
rect 7416 7098 7422 7100
rect 7176 7046 7178 7098
rect 7358 7046 7360 7098
rect 7114 7044 7120 7046
rect 7176 7044 7200 7046
rect 7256 7044 7280 7046
rect 7336 7044 7360 7046
rect 7416 7044 7422 7046
rect 7114 7035 7422 7044
rect 7484 6934 7512 7142
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7576 6254 7604 8842
rect 7668 8634 7696 8910
rect 8220 8838 8248 8978
rect 8312 8945 8340 8978
rect 8298 8936 8354 8945
rect 8298 8871 8354 8880
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 7760 7410 7788 7686
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 8128 7342 8156 7686
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8220 7002 8248 7822
rect 8312 7206 8340 7890
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 7838 6896 7894 6905
rect 7838 6831 7840 6840
rect 7892 6831 7894 6840
rect 7840 6802 7892 6808
rect 7838 6760 7894 6769
rect 7838 6695 7894 6704
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7114 6012 7422 6021
rect 7114 6010 7120 6012
rect 7176 6010 7200 6012
rect 7256 6010 7280 6012
rect 7336 6010 7360 6012
rect 7416 6010 7422 6012
rect 7176 5958 7178 6010
rect 7358 5958 7360 6010
rect 7114 5956 7120 5958
rect 7176 5956 7200 5958
rect 7256 5956 7280 5958
rect 7336 5956 7360 5958
rect 7416 5956 7422 5958
rect 7114 5947 7422 5956
rect 7760 5914 7788 6190
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7748 5704 7800 5710
rect 7852 5692 7880 6695
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8220 5846 8248 6190
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 7800 5664 7880 5692
rect 7748 5646 7800 5652
rect 7930 5536 7986 5545
rect 7930 5471 7986 5480
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7114 4924 7422 4933
rect 7114 4922 7120 4924
rect 7176 4922 7200 4924
rect 7256 4922 7280 4924
rect 7336 4922 7360 4924
rect 7416 4922 7422 4924
rect 7176 4870 7178 4922
rect 7358 4870 7360 4922
rect 7114 4868 7120 4870
rect 7176 4868 7200 4870
rect 7256 4868 7280 4870
rect 7336 4868 7360 4870
rect 7416 4868 7422 4870
rect 7114 4859 7422 4868
rect 7760 4690 7788 4966
rect 7944 4826 7972 5471
rect 8312 5098 8340 7142
rect 8404 6866 8432 8570
rect 8588 8566 8616 8996
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8680 8634 8708 8978
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8496 7954 8524 8434
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8588 6866 8616 8502
rect 8772 8430 8800 9454
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8864 8430 8892 8842
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8680 7750 8708 8298
rect 8772 8090 8800 8366
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8680 6866 8708 7686
rect 8864 7410 8892 7890
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8956 7290 8984 8774
rect 9140 7546 9168 8978
rect 9324 8945 9352 9454
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9416 9042 9444 9318
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9310 8936 9366 8945
rect 9310 8871 9366 8880
rect 9508 8401 9536 8978
rect 9494 8392 9550 8401
rect 9494 8327 9550 8336
rect 9404 8288 9456 8294
rect 9600 8276 9628 10542
rect 9692 9586 9720 11342
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9784 10470 9812 11154
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9692 9217 9720 9522
rect 9678 9208 9734 9217
rect 9678 9143 9734 9152
rect 9692 8498 9720 9143
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9404 8230 9456 8236
rect 9508 8248 9628 8276
rect 9416 7954 9444 8230
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8864 7262 8984 7290
rect 8864 6866 8892 7262
rect 9140 6866 9168 7482
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9416 6866 9444 6938
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8404 4758 8432 5102
rect 8588 5098 8616 6054
rect 8680 5370 8708 6802
rect 8956 6746 8984 6802
rect 9508 6746 9536 8248
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 8864 6718 8984 6746
rect 9220 6724 9272 6730
rect 8864 5778 8892 6718
rect 9220 6666 9272 6672
rect 9416 6718 9536 6746
rect 9588 6724 9640 6730
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8864 5642 8892 5714
rect 9048 5710 9076 6394
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 8576 5092 8628 5098
rect 8576 5034 8628 5040
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8496 4826 8524 4966
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6932 4078 6960 4150
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 7114 3836 7422 3845
rect 7114 3834 7120 3836
rect 7176 3834 7200 3836
rect 7256 3834 7280 3836
rect 7336 3834 7360 3836
rect 7416 3834 7422 3836
rect 7176 3782 7178 3834
rect 7358 3782 7360 3834
rect 7114 3780 7120 3782
rect 7176 3780 7200 3782
rect 7256 3780 7280 3782
rect 7336 3780 7360 3782
rect 7416 3780 7422 3782
rect 7114 3771 7422 3780
rect 7196 2984 7248 2990
rect 7484 2972 7512 4422
rect 8128 4214 8156 4490
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 8404 4078 8432 4694
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8680 4214 8708 4558
rect 8668 4208 8720 4214
rect 8668 4150 8720 4156
rect 8680 4078 8708 4150
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 7576 2990 7604 4014
rect 7668 3398 7696 4014
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7852 3466 7880 3674
rect 8758 3632 8814 3641
rect 9140 3602 9168 5102
rect 8758 3567 8814 3576
rect 9036 3596 9088 3602
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7248 2944 7512 2972
rect 7564 2984 7616 2990
rect 7562 2952 7564 2961
rect 7616 2952 7618 2961
rect 7196 2926 7248 2932
rect 7562 2887 7618 2896
rect 6748 2746 6868 2774
rect 7114 2748 7422 2757
rect 7114 2746 7120 2748
rect 7176 2746 7200 2748
rect 7256 2746 7280 2748
rect 7336 2746 7360 2748
rect 7416 2746 7422 2748
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 6552 2100 6604 2106
rect 6552 2042 6604 2048
rect 6748 1970 6776 2746
rect 7176 2694 7178 2746
rect 7358 2694 7360 2746
rect 7114 2692 7120 2694
rect 7176 2692 7200 2694
rect 7256 2692 7280 2694
rect 7336 2692 7360 2694
rect 7416 2692 7422 2694
rect 7114 2683 7422 2692
rect 7668 2650 7696 3334
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 7760 2530 7788 2586
rect 7392 2514 7788 2530
rect 7852 2514 7880 3402
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7944 2990 7972 3334
rect 7932 2984 7984 2990
rect 8300 2984 8352 2990
rect 7932 2926 7984 2932
rect 8114 2952 8170 2961
rect 8300 2926 8352 2932
rect 8114 2887 8170 2896
rect 8128 2854 8156 2887
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 7380 2508 7788 2514
rect 7432 2502 7788 2508
rect 7840 2508 7892 2514
rect 7380 2450 7432 2456
rect 6736 1964 6788 1970
rect 6736 1906 6788 1912
rect 6368 1896 6420 1902
rect 6368 1838 6420 1844
rect 6644 1760 6696 1766
rect 6644 1702 6696 1708
rect 6656 1494 6684 1702
rect 7114 1660 7422 1669
rect 7114 1658 7120 1660
rect 7176 1658 7200 1660
rect 7256 1658 7280 1660
rect 7336 1658 7360 1660
rect 7416 1658 7422 1660
rect 7176 1606 7178 1658
rect 7358 1606 7360 1658
rect 7114 1604 7120 1606
rect 7176 1604 7200 1606
rect 7256 1604 7280 1606
rect 7336 1604 7360 1606
rect 7416 1604 7422 1606
rect 7114 1595 7422 1604
rect 7484 1562 7512 2502
rect 7840 2450 7892 2456
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7562 2000 7618 2009
rect 7562 1935 7618 1944
rect 7576 1902 7604 1935
rect 7564 1896 7616 1902
rect 7668 1873 7696 2042
rect 7760 1970 7788 2382
rect 7748 1964 7800 1970
rect 7748 1906 7800 1912
rect 7564 1838 7616 1844
rect 7654 1864 7710 1873
rect 7654 1799 7710 1808
rect 7472 1556 7524 1562
rect 7472 1498 7524 1504
rect 6644 1488 6696 1494
rect 6644 1430 6696 1436
rect 7484 746 7512 1498
rect 7668 814 7696 1799
rect 7760 882 7788 1906
rect 8128 1902 8156 2450
rect 8312 2106 8340 2926
rect 8392 2576 8444 2582
rect 8390 2544 8392 2553
rect 8444 2544 8446 2553
rect 8390 2479 8446 2488
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8300 2100 8352 2106
rect 8300 2042 8352 2048
rect 8116 1896 8168 1902
rect 8116 1838 8168 1844
rect 7840 944 7892 950
rect 7840 886 7892 892
rect 7748 876 7800 882
rect 7748 818 7800 824
rect 7656 808 7708 814
rect 7656 750 7708 756
rect 7472 740 7524 746
rect 7472 682 7524 688
rect 7114 572 7422 581
rect 7114 570 7120 572
rect 7176 570 7200 572
rect 7256 570 7280 572
rect 7336 570 7360 572
rect 7416 570 7422 572
rect 7176 518 7178 570
rect 7358 518 7360 570
rect 7114 516 7120 518
rect 7176 516 7200 518
rect 7256 516 7280 518
rect 7336 516 7360 518
rect 7416 516 7422 518
rect 7114 507 7422 516
rect 7852 400 7880 886
rect 8128 814 8156 1838
rect 8496 1834 8524 2246
rect 8484 1828 8536 1834
rect 8484 1770 8536 1776
rect 8772 814 8800 3567
rect 9036 3538 9088 3544
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9048 3194 9076 3538
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 8852 3120 8904 3126
rect 8850 3088 8852 3097
rect 8904 3088 8906 3097
rect 8956 3058 8984 3130
rect 8850 3023 8906 3032
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 9036 2100 9088 2106
rect 9036 2042 9088 2048
rect 9048 1986 9076 2042
rect 8956 1958 9076 1986
rect 8956 1426 8984 1958
rect 9232 1562 9260 6666
rect 9416 5030 9444 6718
rect 9588 6666 9640 6672
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6118 9536 6598
rect 9600 6390 9628 6666
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5778 9536 6054
rect 9692 5914 9720 7958
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9692 5166 9720 5850
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9312 3120 9364 3126
rect 9310 3088 9312 3097
rect 9364 3088 9366 3097
rect 9310 3023 9366 3032
rect 9416 1902 9444 3538
rect 9600 2990 9628 3878
rect 9678 3088 9734 3097
rect 9678 3023 9734 3032
rect 9692 2990 9720 3023
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9692 2854 9720 2926
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9600 2106 9628 2586
rect 9588 2100 9640 2106
rect 9588 2042 9640 2048
rect 9404 1896 9456 1902
rect 9404 1838 9456 1844
rect 9220 1556 9272 1562
rect 9220 1498 9272 1504
rect 8944 1420 8996 1426
rect 8944 1362 8996 1368
rect 8852 1352 8904 1358
rect 8852 1294 8904 1300
rect 8864 882 8892 1294
rect 9036 1284 9088 1290
rect 9036 1226 9088 1232
rect 9048 950 9076 1226
rect 9036 944 9088 950
rect 9036 886 9088 892
rect 8852 876 8904 882
rect 8852 818 8904 824
rect 9048 814 9076 886
rect 8116 808 8168 814
rect 8116 750 8168 756
rect 8760 808 8812 814
rect 8760 750 8812 756
rect 9036 808 9088 814
rect 9036 750 9088 756
rect 9232 746 9260 1498
rect 9416 1358 9444 1838
rect 9508 1834 9720 1850
rect 9508 1828 9732 1834
rect 9508 1822 9680 1828
rect 9508 1562 9536 1822
rect 9680 1770 9732 1776
rect 9784 1562 9812 10406
rect 9876 10169 9904 11562
rect 10060 11286 10088 11591
rect 10140 11562 10192 11568
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10060 10742 10088 11222
rect 10048 10736 10100 10742
rect 10048 10678 10100 10684
rect 9862 10160 9918 10169
rect 9862 10095 9918 10104
rect 10244 8498 10272 11290
rect 10336 10674 10364 11494
rect 10888 11286 10916 12378
rect 10966 12336 11022 12345
rect 10966 12271 10968 12280
rect 11020 12271 11022 12280
rect 11060 12300 11112 12306
rect 10968 12242 11020 12248
rect 11060 12242 11112 12248
rect 11072 12186 11100 12242
rect 10980 12158 11100 12186
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 10980 11626 11008 12158
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10472 10908 10780 10917
rect 10472 10906 10478 10908
rect 10534 10906 10558 10908
rect 10614 10906 10638 10908
rect 10694 10906 10718 10908
rect 10774 10906 10780 10908
rect 10534 10854 10536 10906
rect 10716 10854 10718 10906
rect 10472 10852 10478 10854
rect 10534 10852 10558 10854
rect 10614 10852 10638 10854
rect 10694 10852 10718 10854
rect 10774 10852 10780 10854
rect 10472 10843 10780 10852
rect 11072 10674 11100 11562
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10336 10198 10364 10610
rect 10324 10192 10376 10198
rect 10324 10134 10376 10140
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10336 9518 10364 9862
rect 10472 9820 10780 9829
rect 10472 9818 10478 9820
rect 10534 9818 10558 9820
rect 10614 9818 10638 9820
rect 10694 9818 10718 9820
rect 10774 9818 10780 9820
rect 10534 9766 10536 9818
rect 10716 9766 10718 9818
rect 10472 9764 10478 9766
rect 10534 9764 10558 9766
rect 10614 9764 10638 9766
rect 10694 9764 10718 9766
rect 10774 9764 10780 9766
rect 10472 9755 10780 9764
rect 11072 9518 11100 10610
rect 11256 10606 11284 12174
rect 11348 11218 11376 12582
rect 11624 12374 11652 12718
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11624 11354 11652 11562
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11256 10146 11284 10542
rect 11520 10192 11572 10198
rect 11256 10118 11376 10146
rect 11520 10134 11572 10140
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11256 9722 11284 9998
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10336 8401 10364 9454
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11164 9178 11192 9386
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11348 8906 11376 10118
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 10472 8732 10780 8741
rect 10472 8730 10478 8732
rect 10534 8730 10558 8732
rect 10614 8730 10638 8732
rect 10694 8730 10718 8732
rect 10774 8730 10780 8732
rect 10534 8678 10536 8730
rect 10716 8678 10718 8730
rect 10472 8676 10478 8678
rect 10534 8676 10558 8678
rect 10614 8676 10638 8678
rect 10694 8676 10718 8678
rect 10774 8676 10780 8678
rect 10472 8667 10780 8676
rect 11242 8528 11298 8537
rect 10784 8492 10836 8498
rect 10836 8452 10916 8480
rect 11242 8463 11298 8472
rect 10784 8434 10836 8440
rect 10322 8392 10378 8401
rect 10322 8327 10378 8336
rect 10472 7644 10780 7653
rect 10472 7642 10478 7644
rect 10534 7642 10558 7644
rect 10614 7642 10638 7644
rect 10694 7642 10718 7644
rect 10774 7642 10780 7644
rect 10534 7590 10536 7642
rect 10716 7590 10718 7642
rect 10472 7588 10478 7590
rect 10534 7588 10558 7590
rect 10614 7588 10638 7590
rect 10694 7588 10718 7590
rect 10774 7588 10780 7590
rect 10472 7579 10780 7588
rect 10888 7426 10916 8452
rect 11256 8430 11284 8463
rect 11348 8430 11376 8842
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 10796 7398 10916 7426
rect 10796 7342 10824 7398
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9876 4842 9904 6734
rect 9968 6254 9996 6870
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 6458 10088 6802
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 9968 5370 9996 6190
rect 10060 5370 10088 6190
rect 10152 5846 10180 6598
rect 10244 6322 10272 6598
rect 10336 6458 10364 7210
rect 10796 6934 10824 7278
rect 10784 6928 10836 6934
rect 10784 6870 10836 6876
rect 10874 6896 10930 6905
rect 10874 6831 10930 6840
rect 10416 6792 10468 6798
rect 10414 6760 10416 6769
rect 10468 6760 10470 6769
rect 10414 6695 10470 6704
rect 10428 6662 10456 6695
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10472 6556 10780 6565
rect 10472 6554 10478 6556
rect 10534 6554 10558 6556
rect 10614 6554 10638 6556
rect 10694 6554 10718 6556
rect 10774 6554 10780 6556
rect 10534 6502 10536 6554
rect 10716 6502 10718 6554
rect 10472 6500 10478 6502
rect 10534 6500 10558 6502
rect 10614 6500 10638 6502
rect 10694 6500 10718 6502
rect 10774 6500 10780 6502
rect 10472 6491 10780 6500
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 9876 4814 9996 4842
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9876 4049 9904 4558
rect 9862 4040 9918 4049
rect 9862 3975 9918 3984
rect 9876 3058 9904 3975
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9876 2514 9904 2790
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9968 2378 9996 4814
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10060 4282 10088 4626
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10152 3602 10180 4422
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10336 3058 10364 6258
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10796 5642 10824 6054
rect 10888 5846 10916 6831
rect 10980 6254 11008 8366
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 11072 7546 11100 8298
rect 11348 8294 11376 8366
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11072 7342 11100 7482
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11072 7002 11100 7278
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6322 11100 6598
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10980 5778 11008 6190
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10472 5468 10780 5477
rect 10472 5466 10478 5468
rect 10534 5466 10558 5468
rect 10614 5466 10638 5468
rect 10694 5466 10718 5468
rect 10774 5466 10780 5468
rect 10534 5414 10536 5466
rect 10716 5414 10718 5466
rect 10472 5412 10478 5414
rect 10534 5412 10558 5414
rect 10614 5412 10638 5414
rect 10694 5412 10718 5414
rect 10774 5412 10780 5414
rect 10472 5403 10780 5412
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 10888 4690 10916 5102
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10796 4570 10824 4626
rect 10796 4554 10916 4570
rect 10784 4548 10916 4554
rect 10836 4542 10916 4548
rect 10784 4490 10836 4496
rect 10472 4380 10780 4389
rect 10472 4378 10478 4380
rect 10534 4378 10558 4380
rect 10614 4378 10638 4380
rect 10694 4378 10718 4380
rect 10774 4378 10780 4380
rect 10534 4326 10536 4378
rect 10716 4326 10718 4378
rect 10472 4324 10478 4326
rect 10534 4324 10558 4326
rect 10614 4324 10638 4326
rect 10694 4324 10718 4326
rect 10774 4324 10780 4326
rect 10472 4315 10780 4324
rect 10888 4196 10916 4542
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10796 4168 10916 4196
rect 10796 4078 10824 4168
rect 10980 4078 11008 4422
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10968 4072 11020 4078
rect 11060 4072 11112 4078
rect 10968 4014 11020 4020
rect 11058 4040 11060 4049
rect 11112 4040 11114 4049
rect 10704 3738 10732 4014
rect 10796 3942 10824 4014
rect 11058 3975 11114 3984
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10472 3292 10780 3301
rect 10472 3290 10478 3292
rect 10534 3290 10558 3292
rect 10614 3290 10638 3292
rect 10694 3290 10718 3292
rect 10774 3290 10780 3292
rect 10534 3238 10536 3290
rect 10716 3238 10718 3290
rect 10472 3236 10478 3238
rect 10534 3236 10558 3238
rect 10614 3236 10638 3238
rect 10694 3236 10718 3238
rect 10774 3236 10780 3238
rect 10472 3227 10780 3236
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10980 2990 11008 3674
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10520 2514 10548 2790
rect 11164 2553 11192 7278
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11256 6458 11284 6666
rect 11348 6458 11376 7686
rect 11532 7342 11560 10134
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11624 8265 11652 8298
rect 11610 8256 11666 8265
rect 11610 8191 11666 8200
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11440 7002 11468 7278
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 11348 5914 11376 6190
rect 11440 6118 11468 6734
rect 11716 6730 11744 16612
rect 11888 16594 11940 16600
rect 12348 16652 12400 16658
rect 12438 16623 12440 16632
rect 12348 16594 12400 16600
rect 12492 16623 12494 16632
rect 12440 16594 12492 16600
rect 12164 16176 12216 16182
rect 12162 16144 12164 16153
rect 12216 16144 12218 16153
rect 12162 16079 12218 16088
rect 11980 16040 12032 16046
rect 11978 16008 11980 16017
rect 12032 16008 12034 16017
rect 11978 15943 12034 15952
rect 12164 15972 12216 15978
rect 11992 15706 12020 15943
rect 12216 15932 12296 15960
rect 12164 15914 12216 15920
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12268 15570 12296 15932
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12268 15094 12296 15506
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11900 13530 11928 14350
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11992 12782 12020 13398
rect 12176 13394 12204 14418
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12268 13870 12296 14214
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11808 12238 11836 12718
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 12084 11626 12112 12582
rect 12072 11620 12124 11626
rect 12072 11562 12124 11568
rect 12268 11286 12296 12582
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11992 10266 12020 10474
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 12176 10198 12204 10950
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 12268 10130 12296 10474
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11808 8430 11836 8570
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11808 8072 11836 8366
rect 11992 8362 12020 9862
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 12084 9178 12112 9386
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 12176 8566 12204 9930
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 11808 8044 11928 8072
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11808 7546 11836 7890
rect 11900 7750 11928 8044
rect 12084 7954 12112 8230
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 12084 7342 12112 7890
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 12176 6662 12204 8366
rect 12268 7002 12296 8978
rect 12360 8430 12388 16594
rect 12544 16046 12572 16934
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12636 16250 12664 16594
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12532 16040 12584 16046
rect 12716 16040 12768 16046
rect 12532 15982 12584 15988
rect 12714 16008 12716 16017
rect 12768 16008 12770 16017
rect 12714 15943 12770 15952
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12544 15162 12572 15506
rect 12820 15502 12848 16526
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 12918 12480 14894
rect 12820 14074 12848 15438
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12820 13938 12848 14010
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12544 12714 12572 12854
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12544 12594 12572 12650
rect 12452 12566 12572 12594
rect 12452 11218 12480 12566
rect 12728 12424 12756 13262
rect 12636 12396 12756 12424
rect 12636 11354 12664 12396
rect 12820 12374 12848 13874
rect 12808 12368 12860 12374
rect 12808 12310 12860 12316
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12728 11830 12756 12106
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12452 9674 12480 11154
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12544 10130 12572 10202
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12452 9646 12572 9674
rect 12544 9382 12572 9646
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12438 9208 12494 9217
rect 12438 9143 12494 9152
rect 12452 9042 12480 9143
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12544 8634 12572 8842
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12636 8362 12664 11290
rect 12728 11082 12756 11766
rect 12820 11218 12848 12106
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12820 9926 12848 10066
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12728 9178 12756 9862
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12820 9042 12848 9318
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12348 8288 12400 8294
rect 12348 8230 12400 8236
rect 12360 7410 12388 8230
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12636 7274 12664 8298
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12268 6118 12296 6938
rect 12728 6934 12756 8434
rect 12820 8090 12848 8978
rect 12912 8514 12940 17070
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13004 14958 13032 16050
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 13096 14634 13124 17070
rect 13188 16250 13492 16266
rect 13176 16244 13492 16250
rect 13228 16238 13492 16244
rect 13176 16186 13228 16192
rect 13188 15910 13216 16186
rect 13464 16182 13492 16238
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13556 14770 13584 17070
rect 13830 16892 14138 16901
rect 13830 16890 13836 16892
rect 13892 16890 13916 16892
rect 13972 16890 13996 16892
rect 14052 16890 14076 16892
rect 14132 16890 14138 16892
rect 13892 16838 13894 16890
rect 14074 16838 14076 16890
rect 13830 16836 13836 16838
rect 13892 16836 13916 16838
rect 13972 16836 13996 16838
rect 14052 16836 14076 16838
rect 14132 16836 14138 16838
rect 13830 16827 14138 16836
rect 14384 16794 14412 17070
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14568 16726 14596 17070
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14556 16720 14608 16726
rect 14556 16662 14608 16668
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13740 16046 13768 16390
rect 14646 16144 14702 16153
rect 14646 16079 14702 16088
rect 14660 16046 14688 16079
rect 14752 16046 14780 16934
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15292 16720 15344 16726
rect 15292 16662 15344 16668
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15212 16250 15240 16594
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 13728 16040 13780 16046
rect 14188 16040 14240 16046
rect 13728 15982 13780 15988
rect 14186 16008 14188 16017
rect 14372 16040 14424 16046
rect 14240 16008 14242 16017
rect 14372 15982 14424 15988
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14186 15943 14242 15952
rect 14200 15910 14228 15943
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 13648 15570 13676 15846
rect 13830 15804 14138 15813
rect 13830 15802 13836 15804
rect 13892 15802 13916 15804
rect 13972 15802 13996 15804
rect 14052 15802 14076 15804
rect 14132 15802 14138 15804
rect 13892 15750 13894 15802
rect 14074 15750 14076 15802
rect 13830 15748 13836 15750
rect 13892 15748 13916 15750
rect 13972 15748 13996 15750
rect 14052 15748 14076 15750
rect 14132 15748 14138 15750
rect 13830 15739 14138 15748
rect 14200 15706 14228 15846
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 14200 14958 14228 15642
rect 14384 15638 14412 15982
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 13556 14742 13768 14770
rect 13096 14606 13584 14634
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 13188 13394 13216 13670
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13280 12782 13308 14486
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13004 10674 13032 12650
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 13096 11354 13124 12174
rect 13188 11898 13216 12650
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13188 11218 13216 11562
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12912 8486 13032 8514
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12912 8090 12940 8366
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12820 7002 12848 7822
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11612 6112 11664 6118
rect 12256 6112 12308 6118
rect 11612 6054 11664 6060
rect 12176 6060 12256 6066
rect 12176 6054 12308 6060
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11532 5098 11560 6054
rect 11624 5574 11652 6054
rect 12176 6038 12296 6054
rect 12176 5914 12204 6038
rect 12254 5944 12310 5953
rect 12164 5908 12216 5914
rect 12254 5879 12256 5888
rect 12164 5850 12216 5856
rect 12308 5879 12310 5888
rect 12256 5850 12308 5856
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11716 4078 11744 5510
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11900 4078 11928 4966
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 12084 4162 12112 4694
rect 12544 4690 12572 5782
rect 12820 5778 12848 6938
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12636 4826 12664 5102
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12176 4282 12204 4626
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12544 4214 12572 4626
rect 12532 4208 12584 4214
rect 12084 4146 12388 4162
rect 12532 4150 12584 4156
rect 12084 4140 12400 4146
rect 12084 4134 12348 4140
rect 12348 4082 12400 4088
rect 11520 4072 11572 4078
rect 11348 4020 11520 4026
rect 11348 4014 11572 4020
rect 11704 4072 11756 4078
rect 11796 4072 11848 4078
rect 11704 4014 11756 4020
rect 11794 4040 11796 4049
rect 11888 4072 11940 4078
rect 11848 4040 11850 4049
rect 11348 3998 11560 4014
rect 11348 3942 11376 3998
rect 11888 4014 11940 4020
rect 11794 3975 11850 3984
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 12256 4004 12308 4010
rect 12256 3946 12308 3952
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3670 11468 3878
rect 12084 3670 12112 3946
rect 12268 3738 12296 3946
rect 12256 3732 12308 3738
rect 12176 3692 12256 3720
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11440 2582 11468 3062
rect 11532 2990 11560 3538
rect 12176 2990 12204 3692
rect 12256 3674 12308 3680
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12268 3194 12296 3538
rect 12360 3398 12388 3946
rect 12636 3584 12664 4762
rect 12728 3738 12756 5646
rect 12820 3942 12848 5714
rect 12912 5370 12940 6802
rect 13004 5914 13032 8486
rect 13096 7018 13124 11018
rect 13188 9722 13216 11018
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13188 9217 13216 9658
rect 13280 9654 13308 12718
rect 13372 11014 13400 12718
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13464 12209 13492 12582
rect 13450 12200 13506 12209
rect 13450 12135 13506 12144
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13464 11354 13492 11834
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13464 10266 13492 11154
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13372 9994 13400 10066
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13268 9648 13320 9654
rect 13464 9602 13492 9998
rect 13268 9590 13320 9596
rect 13174 9208 13230 9217
rect 13174 9143 13230 9152
rect 13280 9110 13308 9590
rect 13372 9574 13492 9602
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13372 8498 13400 9574
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13266 8256 13322 8265
rect 13266 8191 13322 8200
rect 13280 8022 13308 8191
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13188 7342 13216 7686
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13280 7274 13308 7958
rect 13360 7812 13412 7818
rect 13360 7754 13412 7760
rect 13372 7546 13400 7754
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13268 7268 13320 7274
rect 13268 7210 13320 7216
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13096 6990 13308 7018
rect 13176 6928 13228 6934
rect 13176 6870 13228 6876
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 13004 5250 13032 5646
rect 12912 5222 13032 5250
rect 12912 4690 12940 5222
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 13004 3602 13032 5034
rect 12716 3596 12768 3602
rect 12636 3556 12716 3584
rect 12716 3538 12768 3544
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12268 2990 12296 3130
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 11428 2576 11480 2582
rect 11150 2544 11206 2553
rect 10508 2508 10560 2514
rect 11428 2518 11480 2524
rect 11150 2479 11206 2488
rect 10508 2450 10560 2456
rect 9956 2372 10008 2378
rect 9956 2314 10008 2320
rect 9496 1556 9548 1562
rect 9496 1498 9548 1504
rect 9772 1556 9824 1562
rect 9772 1498 9824 1504
rect 9404 1352 9456 1358
rect 9404 1294 9456 1300
rect 9588 944 9640 950
rect 9588 886 9640 892
rect 9220 740 9272 746
rect 9220 682 9272 688
rect 9600 400 9628 886
rect 9968 746 9996 2314
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10336 1902 10364 2246
rect 10472 2204 10780 2213
rect 10472 2202 10478 2204
rect 10534 2202 10558 2204
rect 10614 2202 10638 2204
rect 10694 2202 10718 2204
rect 10774 2202 10780 2204
rect 10534 2150 10536 2202
rect 10716 2150 10718 2202
rect 10472 2148 10478 2150
rect 10534 2148 10558 2150
rect 10614 2148 10638 2150
rect 10694 2148 10718 2150
rect 10774 2148 10780 2150
rect 10472 2139 10780 2148
rect 10324 1896 10376 1902
rect 10324 1838 10376 1844
rect 10232 1760 10284 1766
rect 10232 1702 10284 1708
rect 10244 1494 10272 1702
rect 10324 1556 10376 1562
rect 10324 1498 10376 1504
rect 10232 1488 10284 1494
rect 10232 1430 10284 1436
rect 10336 882 10364 1498
rect 10472 1116 10780 1125
rect 10472 1114 10478 1116
rect 10534 1114 10558 1116
rect 10614 1114 10638 1116
rect 10694 1114 10718 1116
rect 10774 1114 10780 1116
rect 10534 1062 10536 1114
rect 10716 1062 10718 1114
rect 10472 1060 10478 1062
rect 10534 1060 10558 1062
rect 10614 1060 10638 1062
rect 10694 1060 10718 1062
rect 10774 1060 10780 1062
rect 10472 1051 10780 1060
rect 10324 876 10376 882
rect 10324 818 10376 824
rect 11164 746 11192 2479
rect 11532 2394 11560 2926
rect 11624 2854 11652 2926
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11440 2366 11560 2394
rect 11336 1760 11388 1766
rect 11336 1702 11388 1708
rect 11348 1494 11376 1702
rect 11440 1562 11468 2366
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11532 1902 11560 2246
rect 11520 1896 11572 1902
rect 11520 1838 11572 1844
rect 11428 1556 11480 1562
rect 11428 1498 11480 1504
rect 11336 1488 11388 1494
rect 11336 1430 11388 1436
rect 11336 944 11388 950
rect 11336 886 11388 892
rect 9956 740 10008 746
rect 9956 682 10008 688
rect 11152 740 11204 746
rect 11152 682 11204 688
rect 11348 400 11376 886
rect 11624 814 11652 2790
rect 12452 2514 12480 3130
rect 12544 2582 12572 3334
rect 12820 2922 12848 3538
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 12728 1902 12756 2382
rect 12820 1970 12848 2858
rect 12808 1964 12860 1970
rect 12808 1906 12860 1912
rect 12716 1896 12768 1902
rect 12716 1838 12768 1844
rect 12900 1828 12952 1834
rect 12900 1770 12952 1776
rect 12808 1760 12860 1766
rect 12808 1702 12860 1708
rect 12820 1494 12848 1702
rect 12912 1494 12940 1770
rect 13004 1562 13032 3538
rect 13096 3194 13124 6734
rect 13188 4826 13216 6870
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13280 3670 13308 6990
rect 13372 6610 13400 7142
rect 13464 6798 13492 9454
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13372 6582 13492 6610
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13372 4758 13400 5782
rect 13464 5778 13492 6582
rect 13556 5930 13584 14606
rect 13740 12434 13768 14742
rect 13830 14716 14138 14725
rect 13830 14714 13836 14716
rect 13892 14714 13916 14716
rect 13972 14714 13996 14716
rect 14052 14714 14076 14716
rect 14132 14714 14138 14716
rect 13892 14662 13894 14714
rect 14074 14662 14076 14714
rect 13830 14660 13836 14662
rect 13892 14660 13916 14662
rect 13972 14660 13996 14662
rect 14052 14660 14076 14662
rect 14132 14660 14138 14662
rect 13830 14651 14138 14660
rect 15212 14550 15240 15302
rect 15304 14890 15332 16662
rect 15396 16046 15424 16730
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13832 13870 13860 14214
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 13830 13628 14138 13637
rect 13830 13626 13836 13628
rect 13892 13626 13916 13628
rect 13972 13626 13996 13628
rect 14052 13626 14076 13628
rect 14132 13626 14138 13628
rect 13892 13574 13894 13626
rect 14074 13574 14076 13626
rect 13830 13572 13836 13574
rect 13892 13572 13916 13574
rect 13972 13572 13996 13574
rect 14052 13572 14076 13574
rect 14132 13572 14138 13574
rect 13830 13563 14138 13572
rect 14292 13530 14320 13670
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14384 13462 14412 13738
rect 14372 13456 14424 13462
rect 14372 13398 14424 13404
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 13830 12540 14138 12549
rect 13830 12538 13836 12540
rect 13892 12538 13916 12540
rect 13972 12538 13996 12540
rect 14052 12538 14076 12540
rect 14132 12538 14138 12540
rect 13892 12486 13894 12538
rect 14074 12486 14076 12538
rect 13830 12484 13836 12486
rect 13892 12484 13916 12486
rect 13972 12484 13996 12486
rect 14052 12484 14076 12486
rect 14132 12484 14138 12486
rect 13830 12475 14138 12484
rect 13648 12406 13768 12434
rect 13648 8650 13676 12406
rect 14200 12374 14228 12922
rect 14292 12714 14320 13330
rect 14476 13326 14504 14418
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 15120 14074 15148 14350
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 15120 13462 15148 14010
rect 15200 13864 15252 13870
rect 15304 13852 15332 14826
rect 15252 13824 15332 13852
rect 15200 13806 15252 13812
rect 15108 13456 15160 13462
rect 15108 13398 15160 13404
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14752 12442 14780 13262
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14844 12306 14872 12582
rect 14936 12442 14964 13262
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15120 12782 15148 13126
rect 15212 12850 15240 13806
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 15014 12200 15070 12209
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13740 11898 13768 12038
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13832 11694 13860 12038
rect 14568 11898 14596 12174
rect 15014 12135 15070 12144
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13830 11452 14138 11461
rect 13830 11450 13836 11452
rect 13892 11450 13916 11452
rect 13972 11450 13996 11452
rect 14052 11450 14076 11452
rect 14132 11450 14138 11452
rect 13892 11398 13894 11450
rect 14074 11398 14076 11450
rect 13830 11396 13836 11398
rect 13892 11396 13916 11398
rect 13972 11396 13996 11398
rect 14052 11396 14076 11398
rect 14132 11396 14138 11398
rect 13830 11387 14138 11396
rect 14568 11150 14596 11834
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14844 11218 14872 11290
rect 14832 11212 14884 11218
rect 14752 11172 14832 11200
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14752 10674 14780 11172
rect 15028 11200 15056 12135
rect 15120 11336 15148 12242
rect 15212 11694 15240 12786
rect 15304 12782 15332 12922
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15488 11354 15516 12718
rect 15476 11348 15528 11354
rect 15120 11308 15240 11336
rect 15108 11212 15160 11218
rect 15028 11172 15108 11200
rect 14832 11154 14884 11160
rect 15108 11154 15160 11160
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10112 13768 10406
rect 13830 10364 14138 10373
rect 13830 10362 13836 10364
rect 13892 10362 13916 10364
rect 13972 10362 13996 10364
rect 14052 10362 14076 10364
rect 14132 10362 14138 10364
rect 13892 10310 13894 10362
rect 14074 10310 14076 10362
rect 13830 10308 13836 10310
rect 13892 10308 13916 10310
rect 13972 10308 13996 10310
rect 14052 10308 14076 10310
rect 14132 10308 14138 10310
rect 13830 10299 14138 10308
rect 14844 10130 14872 10610
rect 15212 10266 15240 11308
rect 15476 11290 15528 11296
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15396 10130 15424 10406
rect 13820 10124 13872 10130
rect 13740 10084 13820 10112
rect 13820 10066 13872 10072
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 14200 9994 14228 10066
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14278 9616 14334 9625
rect 14278 9551 14280 9560
rect 14332 9551 14334 9560
rect 14280 9522 14332 9528
rect 13830 9276 14138 9285
rect 13830 9274 13836 9276
rect 13892 9274 13916 9276
rect 13972 9274 13996 9276
rect 14052 9274 14076 9276
rect 14132 9274 14138 9276
rect 13892 9222 13894 9274
rect 14074 9222 14076 9274
rect 13830 9220 13836 9222
rect 13892 9220 13916 9222
rect 13972 9220 13996 9222
rect 14052 9220 14076 9222
rect 14132 9220 14138 9222
rect 13830 9211 14138 9220
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 13648 8622 13768 8650
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13648 7478 13676 8366
rect 13740 7970 13768 8622
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 13830 8188 14138 8197
rect 13830 8186 13836 8188
rect 13892 8186 13916 8188
rect 13972 8186 13996 8188
rect 14052 8186 14076 8188
rect 14132 8186 14138 8188
rect 13892 8134 13894 8186
rect 14074 8134 14076 8186
rect 13830 8132 13836 8134
rect 13892 8132 13916 8134
rect 13972 8132 13996 8134
rect 14052 8132 14076 8134
rect 14132 8132 14138 8134
rect 13830 8123 14138 8132
rect 13740 7942 13860 7970
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13740 7546 13768 7822
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13636 7472 13688 7478
rect 13832 7426 13860 7942
rect 13636 7414 13688 7420
rect 13740 7398 13860 7426
rect 13740 6100 13768 7398
rect 14200 7342 14228 8230
rect 14384 8022 14412 8366
rect 14568 8022 14596 8978
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 14556 8016 14608 8022
rect 14556 7958 14608 7964
rect 14844 7954 14872 8230
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14752 7818 14780 7890
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 15028 7206 15056 9998
rect 15396 9450 15424 10066
rect 15488 9722 15516 11154
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15384 9444 15436 9450
rect 15384 9386 15436 9392
rect 15106 8392 15162 8401
rect 15106 8327 15162 8336
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 13830 7100 14138 7109
rect 13830 7098 13836 7100
rect 13892 7098 13916 7100
rect 13972 7098 13996 7100
rect 14052 7098 14076 7100
rect 14132 7098 14138 7100
rect 13892 7046 13894 7098
rect 14074 7046 14076 7098
rect 13830 7044 13836 7046
rect 13892 7044 13916 7046
rect 13972 7044 13996 7046
rect 14052 7044 14076 7046
rect 14132 7044 14138 7046
rect 13830 7035 14138 7044
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 13832 6310 14504 6338
rect 13832 6254 13860 6310
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 13740 6072 14228 6100
rect 13830 6012 14138 6021
rect 13830 6010 13836 6012
rect 13892 6010 13916 6012
rect 13972 6010 13996 6012
rect 14052 6010 14076 6012
rect 14132 6010 14138 6012
rect 13892 5958 13894 6010
rect 14074 5958 14076 6010
rect 13830 5956 13836 5958
rect 13892 5956 13916 5958
rect 13972 5956 13996 5958
rect 14052 5956 14076 5958
rect 14132 5956 14138 5958
rect 13830 5947 14138 5956
rect 13556 5902 13676 5930
rect 14200 5914 14228 6072
rect 13648 5896 13676 5902
rect 13820 5908 13872 5914
rect 13648 5868 13820 5896
rect 13820 5850 13872 5856
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 13464 5273 13492 5714
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13450 5264 13506 5273
rect 13450 5199 13506 5208
rect 13360 4752 13412 4758
rect 13360 4694 13412 4700
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13636 3664 13688 3670
rect 13636 3606 13688 3612
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13188 3126 13216 3334
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13648 1816 13676 3606
rect 13740 3126 13768 5306
rect 13830 4924 14138 4933
rect 13830 4922 13836 4924
rect 13892 4922 13916 4924
rect 13972 4922 13996 4924
rect 14052 4922 14076 4924
rect 14132 4922 14138 4924
rect 13892 4870 13894 4922
rect 14074 4870 14076 4922
rect 13830 4868 13836 4870
rect 13892 4868 13916 4870
rect 13972 4868 13996 4870
rect 14052 4868 14076 4870
rect 14132 4868 14138 4870
rect 13830 4859 14138 4868
rect 14200 4826 14228 5714
rect 14292 5574 14320 6190
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14292 5166 14320 5510
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14384 4826 14412 5646
rect 14476 5166 14504 6310
rect 14568 5778 14596 6394
rect 15028 5846 15056 7142
rect 15120 5914 15148 8327
rect 15488 7954 15516 9658
rect 15200 7948 15252 7954
rect 15476 7948 15528 7954
rect 15252 7908 15332 7936
rect 15200 7890 15252 7896
rect 15304 7546 15332 7908
rect 15476 7890 15528 7896
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15396 7274 15424 7686
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15016 5840 15068 5846
rect 15016 5782 15068 5788
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 13830 3836 14138 3845
rect 13830 3834 13836 3836
rect 13892 3834 13916 3836
rect 13972 3834 13996 3836
rect 14052 3834 14076 3836
rect 14132 3834 14138 3836
rect 13892 3782 13894 3834
rect 14074 3782 14076 3834
rect 13830 3780 13836 3782
rect 13892 3780 13916 3782
rect 13972 3780 13996 3782
rect 14052 3780 14076 3782
rect 14132 3780 14138 3782
rect 13830 3771 14138 3780
rect 14200 3534 14228 4014
rect 14292 3641 14320 4558
rect 14384 4010 14412 4626
rect 15028 4622 15056 5102
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14278 3632 14334 3641
rect 14278 3567 14334 3576
rect 14004 3528 14056 3534
rect 13910 3496 13966 3505
rect 14004 3470 14056 3476
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 13910 3431 13966 3440
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13740 2990 13768 3062
rect 13924 2990 13952 3431
rect 14016 3058 14044 3470
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13740 2038 13768 2926
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 13830 2748 14138 2757
rect 13830 2746 13836 2748
rect 13892 2746 13916 2748
rect 13972 2746 13996 2748
rect 14052 2746 14076 2748
rect 14132 2746 14138 2748
rect 13892 2694 13894 2746
rect 14074 2694 14076 2746
rect 13830 2692 13836 2694
rect 13892 2692 13916 2694
rect 13972 2692 13996 2694
rect 14052 2692 14076 2694
rect 14132 2692 14138 2694
rect 13830 2683 14138 2692
rect 13728 2032 13780 2038
rect 13728 1974 13780 1980
rect 13912 1828 13964 1834
rect 13648 1788 13912 1816
rect 13912 1770 13964 1776
rect 13830 1660 14138 1669
rect 13830 1658 13836 1660
rect 13892 1658 13916 1660
rect 13972 1658 13996 1660
rect 14052 1658 14076 1660
rect 14132 1658 14138 1660
rect 13892 1606 13894 1658
rect 14074 1606 14076 1658
rect 13830 1604 13836 1606
rect 13892 1604 13916 1606
rect 13972 1604 13996 1606
rect 14052 1604 14076 1606
rect 14132 1604 14138 1606
rect 13830 1595 14138 1604
rect 14200 1562 14228 2858
rect 14292 2650 14320 3470
rect 14476 3058 14504 4558
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15120 3738 15148 4014
rect 15212 3738 15240 5646
rect 15396 4758 15424 5714
rect 15580 5114 15608 17002
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15672 14482 15700 14758
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15764 12345 15792 12650
rect 15750 12336 15806 12345
rect 15750 12271 15806 12280
rect 15764 11218 15792 12271
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15672 10130 15700 10542
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15672 8566 15700 8978
rect 15764 8906 15792 10066
rect 15752 8900 15804 8906
rect 15752 8842 15804 8848
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 15856 6202 15884 17070
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15948 14618 15976 14894
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 16040 11558 16068 16662
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16224 15026 16252 15506
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 16132 13530 16160 13738
rect 16224 13734 16252 14962
rect 16408 14618 16436 15506
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16408 13394 16436 14554
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16500 14074 16528 14350
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16592 13546 16620 17206
rect 16868 17134 16896 17600
rect 17512 17542 17540 17600
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17188 17436 17496 17445
rect 17188 17434 17194 17436
rect 17250 17434 17274 17436
rect 17330 17434 17354 17436
rect 17410 17434 17434 17436
rect 17490 17434 17496 17436
rect 17250 17382 17252 17434
rect 17432 17382 17434 17434
rect 17188 17380 17194 17382
rect 17250 17380 17274 17382
rect 17330 17380 17354 17382
rect 17410 17380 17434 17382
rect 17490 17380 17496 17382
rect 17188 17371 17496 17380
rect 17788 17134 17816 17478
rect 19444 17134 19472 17600
rect 21652 17134 21680 17734
rect 22006 17600 22062 18000
rect 22650 17600 22706 18000
rect 23294 17600 23350 18000
rect 23938 17762 23994 18000
rect 23768 17734 23994 17762
rect 22020 17134 22048 17600
rect 22664 17134 22692 17600
rect 23308 17134 23336 17600
rect 23768 17134 23796 17734
rect 23938 17600 23994 17734
rect 24582 17600 24638 18000
rect 25226 17600 25282 18000
rect 25870 17600 25926 18000
rect 26514 17600 26570 18000
rect 27158 17600 27214 18000
rect 23904 17436 24212 17445
rect 23904 17434 23910 17436
rect 23966 17434 23990 17436
rect 24046 17434 24070 17436
rect 24126 17434 24150 17436
rect 24206 17434 24212 17436
rect 23966 17382 23968 17434
rect 24148 17382 24150 17434
rect 23904 17380 23910 17382
rect 23966 17380 23990 17382
rect 24046 17380 24070 17382
rect 24126 17380 24150 17382
rect 24206 17380 24212 17382
rect 23904 17371 24212 17380
rect 24596 17134 24624 17600
rect 25240 17202 25268 17600
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 22008 17128 22060 17134
rect 22008 17070 22060 17076
rect 22652 17128 22704 17134
rect 22652 17070 22704 17076
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23756 17128 23808 17134
rect 23756 17070 23808 17076
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 25780 17128 25832 17134
rect 25780 17070 25832 17076
rect 19524 17060 19576 17066
rect 19524 17002 19576 17008
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 16684 16726 16712 16934
rect 16672 16720 16724 16726
rect 16672 16662 16724 16668
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16684 14822 16712 15506
rect 16776 15162 16804 15506
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16776 13954 16804 15098
rect 16500 13518 16620 13546
rect 16684 13926 16804 13954
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16316 12238 16344 12922
rect 16500 12866 16528 13518
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16408 12838 16528 12866
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16132 11626 16160 12038
rect 16408 11898 16436 12838
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16500 12442 16528 12718
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16304 10192 16356 10198
rect 16304 10134 16356 10140
rect 16316 10062 16344 10134
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16316 9722 16344 9998
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16026 9480 16082 9489
rect 16026 9415 16028 9424
rect 16080 9415 16082 9424
rect 16028 9386 16080 9392
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15948 8634 15976 8978
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 16500 8498 16528 11562
rect 16592 10810 16620 13330
rect 16684 13258 16712 13926
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16776 13258 16804 13330
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16684 12850 16712 13194
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16684 12306 16712 12650
rect 16776 12374 16804 13194
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16580 9104 16632 9110
rect 16580 9046 16632 9052
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16316 6662 16344 8434
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16500 7206 16528 8298
rect 16592 8022 16620 9046
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16592 7342 16620 7958
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16500 7002 16528 7142
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15764 6174 15884 6202
rect 15672 5710 15700 6122
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15672 5234 15700 5646
rect 15764 5370 15792 6174
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15856 5778 15884 6054
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15488 5086 15608 5114
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14476 2514 14504 2790
rect 15304 2582 15332 3946
rect 15488 3466 15516 5086
rect 15672 4010 15700 5170
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 16040 3738 16068 5102
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14464 2508 14516 2514
rect 14516 2468 14596 2496
rect 14464 2450 14516 2456
rect 14384 1766 14412 2450
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 14476 1902 14504 2314
rect 14464 1896 14516 1902
rect 14464 1838 14516 1844
rect 14372 1760 14424 1766
rect 14372 1702 14424 1708
rect 12992 1556 13044 1562
rect 12992 1498 13044 1504
rect 14188 1556 14240 1562
rect 14188 1498 14240 1504
rect 12808 1488 12860 1494
rect 12808 1430 12860 1436
rect 12900 1488 12952 1494
rect 12900 1430 12952 1436
rect 12716 1216 12768 1222
rect 12716 1158 12768 1164
rect 12728 950 12756 1158
rect 13004 950 13032 1498
rect 13912 1352 13964 1358
rect 13912 1294 13964 1300
rect 12716 944 12768 950
rect 12716 886 12768 892
rect 12992 944 13044 950
rect 12992 886 13044 892
rect 13084 944 13136 950
rect 13084 886 13136 892
rect 11612 808 11664 814
rect 11612 750 11664 756
rect 13096 400 13124 886
rect 13924 746 13952 1294
rect 14384 1222 14412 1702
rect 14568 1426 14596 2468
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14556 1420 14608 1426
rect 14556 1362 14608 1368
rect 14372 1216 14424 1222
rect 14372 1158 14424 1164
rect 14384 814 14412 1158
rect 14752 950 14780 2246
rect 15672 2106 15700 3470
rect 15856 2990 15884 3606
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15660 2100 15712 2106
rect 15660 2042 15712 2048
rect 15568 1896 15620 1902
rect 15568 1838 15620 1844
rect 15108 1760 15160 1766
rect 15108 1702 15160 1708
rect 15120 1494 15148 1702
rect 15108 1488 15160 1494
rect 15108 1430 15160 1436
rect 15580 1426 15608 1838
rect 15856 1766 15884 2926
rect 16040 2922 16068 3402
rect 16132 2922 16160 5850
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 16224 3194 16252 5238
rect 16408 4758 16436 6258
rect 16684 5098 16712 10202
rect 16868 10010 16896 16594
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16960 13530 16988 15438
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16960 12782 16988 13262
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16960 11898 16988 12174
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 17052 10266 17080 16934
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 17144 16697 17172 16730
rect 17130 16688 17186 16697
rect 17130 16623 17186 16632
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 18144 16516 18196 16522
rect 18144 16458 18196 16464
rect 17188 16348 17496 16357
rect 17188 16346 17194 16348
rect 17250 16346 17274 16348
rect 17330 16346 17354 16348
rect 17410 16346 17434 16348
rect 17490 16346 17496 16348
rect 17250 16294 17252 16346
rect 17432 16294 17434 16346
rect 17188 16292 17194 16294
rect 17250 16292 17274 16294
rect 17330 16292 17354 16294
rect 17410 16292 17434 16294
rect 17490 16292 17496 16294
rect 17188 16283 17496 16292
rect 17696 16182 17724 16458
rect 18156 16250 18184 16458
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17958 15600 18014 15609
rect 17958 15535 18014 15544
rect 17776 15360 17828 15366
rect 17828 15320 17908 15348
rect 17776 15302 17828 15308
rect 17188 15260 17496 15269
rect 17188 15258 17194 15260
rect 17250 15258 17274 15260
rect 17330 15258 17354 15260
rect 17410 15258 17434 15260
rect 17490 15258 17496 15260
rect 17250 15206 17252 15258
rect 17432 15206 17434 15258
rect 17188 15204 17194 15206
rect 17250 15204 17274 15206
rect 17330 15204 17354 15206
rect 17410 15204 17434 15206
rect 17490 15204 17496 15206
rect 17188 15195 17496 15204
rect 17684 14884 17736 14890
rect 17684 14826 17736 14832
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17236 14482 17264 14758
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 17188 14172 17496 14181
rect 17188 14170 17194 14172
rect 17250 14170 17274 14172
rect 17330 14170 17354 14172
rect 17410 14170 17434 14172
rect 17490 14170 17496 14172
rect 17250 14118 17252 14170
rect 17432 14118 17434 14170
rect 17188 14116 17194 14118
rect 17250 14116 17274 14118
rect 17330 14116 17354 14118
rect 17410 14116 17434 14118
rect 17490 14116 17496 14118
rect 17188 14107 17496 14116
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17512 13308 17540 14010
rect 17696 13530 17724 14826
rect 17880 14414 17908 15320
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17880 13870 17908 14350
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17774 13560 17830 13569
rect 17684 13524 17736 13530
rect 17774 13495 17776 13504
rect 17684 13466 17736 13472
rect 17828 13495 17830 13504
rect 17776 13466 17828 13472
rect 17684 13388 17736 13394
rect 17736 13348 17816 13376
rect 17684 13330 17736 13336
rect 17592 13320 17644 13326
rect 17512 13280 17592 13308
rect 17592 13262 17644 13268
rect 17188 13084 17496 13093
rect 17188 13082 17194 13084
rect 17250 13082 17274 13084
rect 17330 13082 17354 13084
rect 17410 13082 17434 13084
rect 17490 13082 17496 13084
rect 17250 13030 17252 13082
rect 17432 13030 17434 13082
rect 17188 13028 17194 13030
rect 17250 13028 17274 13030
rect 17330 13028 17354 13030
rect 17410 13028 17434 13030
rect 17490 13028 17496 13030
rect 17188 13019 17496 13028
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17188 11996 17496 12005
rect 17188 11994 17194 11996
rect 17250 11994 17274 11996
rect 17330 11994 17354 11996
rect 17410 11994 17434 11996
rect 17490 11994 17496 11996
rect 17250 11942 17252 11994
rect 17432 11942 17434 11994
rect 17188 11940 17194 11942
rect 17250 11940 17274 11942
rect 17330 11940 17354 11942
rect 17410 11940 17434 11942
rect 17490 11940 17496 11942
rect 17188 11931 17496 11940
rect 17604 11082 17632 12242
rect 17696 11694 17724 12582
rect 17684 11688 17736 11694
rect 17684 11630 17736 11636
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17188 10908 17496 10917
rect 17188 10906 17194 10908
rect 17250 10906 17274 10908
rect 17330 10906 17354 10908
rect 17410 10906 17434 10908
rect 17490 10906 17496 10908
rect 17250 10854 17252 10906
rect 17432 10854 17434 10906
rect 17188 10852 17194 10854
rect 17250 10852 17274 10854
rect 17330 10852 17354 10854
rect 17410 10852 17434 10854
rect 17490 10852 17496 10854
rect 17188 10843 17496 10852
rect 17592 10532 17644 10538
rect 17592 10474 17644 10480
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 16868 9982 16988 10010
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16868 9518 16896 9862
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16776 9178 16804 9318
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16776 8430 16804 9114
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16960 7342 16988 9982
rect 17052 9160 17080 10066
rect 17188 9820 17496 9829
rect 17188 9818 17194 9820
rect 17250 9818 17274 9820
rect 17330 9818 17354 9820
rect 17410 9818 17434 9820
rect 17490 9818 17496 9820
rect 17250 9766 17252 9818
rect 17432 9766 17434 9818
rect 17188 9764 17194 9766
rect 17250 9764 17274 9766
rect 17330 9764 17354 9766
rect 17410 9764 17434 9766
rect 17490 9764 17496 9766
rect 17188 9755 17496 9764
rect 17604 9654 17632 10474
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17696 10266 17724 10406
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17052 9132 17172 9160
rect 17144 8974 17172 9132
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17188 8732 17496 8741
rect 17188 8730 17194 8732
rect 17250 8730 17274 8732
rect 17330 8730 17354 8732
rect 17410 8730 17434 8732
rect 17490 8730 17496 8732
rect 17250 8678 17252 8730
rect 17432 8678 17434 8730
rect 17188 8676 17194 8678
rect 17250 8676 17274 8678
rect 17330 8676 17354 8678
rect 17410 8676 17434 8678
rect 17490 8676 17496 8678
rect 17188 8667 17496 8676
rect 17604 8498 17632 9454
rect 17696 8974 17724 9862
rect 17788 9654 17816 13348
rect 17880 12918 17908 13806
rect 17972 13410 18000 15535
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18064 14550 18092 14894
rect 18144 14884 18196 14890
rect 18144 14826 18196 14832
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 18156 14006 18184 14826
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 17972 13382 18092 13410
rect 18248 13397 18276 13738
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 17972 12764 18000 13262
rect 17880 12736 18000 12764
rect 17880 12306 17908 12736
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17880 11286 17908 12242
rect 17972 11354 18000 12242
rect 18064 11626 18092 13382
rect 18236 13391 18288 13397
rect 18236 13333 18288 13339
rect 18420 13388 18472 13394
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18156 12306 18184 13126
rect 18248 12986 18276 13333
rect 18420 13330 18472 13336
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18052 11620 18104 11626
rect 18052 11562 18104 11568
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18064 10606 18092 10950
rect 18144 10804 18196 10810
rect 18144 10746 18196 10752
rect 18156 10606 18184 10746
rect 18248 10674 18276 12650
rect 18340 12442 18368 12718
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18432 12374 18460 13330
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18432 11898 18460 12310
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 17880 10266 17908 10542
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17880 9450 17908 9862
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 18156 9330 18184 10542
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18248 9586 18276 9998
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 17880 9302 18184 9330
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17604 8022 17632 8434
rect 17788 8430 17816 8774
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17592 8016 17644 8022
rect 17592 7958 17644 7964
rect 17188 7644 17496 7653
rect 17188 7642 17194 7644
rect 17250 7642 17274 7644
rect 17330 7642 17354 7644
rect 17410 7642 17434 7644
rect 17490 7642 17496 7644
rect 17250 7590 17252 7642
rect 17432 7590 17434 7642
rect 17188 7588 17194 7590
rect 17250 7588 17274 7590
rect 17330 7588 17354 7590
rect 17410 7588 17434 7590
rect 17490 7588 17496 7590
rect 17188 7579 17496 7588
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16868 6186 16896 7278
rect 16960 6254 16988 7278
rect 17604 6798 17632 7958
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17788 6934 17816 7686
rect 17880 7410 17908 9302
rect 18248 9178 18276 9522
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 18050 9072 18106 9081
rect 17972 8566 18000 9046
rect 18248 9042 18276 9114
rect 18050 9007 18106 9016
rect 18236 9036 18288 9042
rect 18064 8974 18092 9007
rect 18236 8978 18288 8984
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 18340 7886 18368 8230
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17776 6928 17828 6934
rect 17776 6870 17828 6876
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17188 6556 17496 6565
rect 17188 6554 17194 6556
rect 17250 6554 17274 6556
rect 17330 6554 17354 6556
rect 17410 6554 17434 6556
rect 17490 6554 17496 6556
rect 17250 6502 17252 6554
rect 17432 6502 17434 6554
rect 17188 6500 17194 6502
rect 17250 6500 17274 6502
rect 17330 6500 17354 6502
rect 17410 6500 17434 6502
rect 17490 6500 17496 6502
rect 17188 6491 17496 6500
rect 17604 6322 17632 6734
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16868 5710 16896 6122
rect 17696 5914 17724 6394
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 16856 5704 16908 5710
rect 16908 5664 16988 5692
rect 16856 5646 16908 5652
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16868 5166 16896 5510
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16672 5092 16724 5098
rect 16672 5034 16724 5040
rect 16684 4842 16712 5034
rect 16684 4814 16896 4842
rect 16396 4752 16448 4758
rect 16394 4720 16396 4729
rect 16448 4720 16450 4729
rect 16394 4655 16450 4664
rect 16580 4684 16632 4690
rect 16408 4146 16436 4655
rect 16580 4626 16632 4632
rect 16592 4282 16620 4626
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16408 3466 16436 4082
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16396 3460 16448 3466
rect 16396 3402 16448 3408
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16500 2990 16528 3674
rect 16592 3058 16620 4218
rect 16776 4214 16804 4422
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16776 3738 16804 3946
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16868 3534 16896 4814
rect 16960 4214 16988 5664
rect 17188 5468 17496 5477
rect 17188 5466 17194 5468
rect 17250 5466 17274 5468
rect 17330 5466 17354 5468
rect 17410 5466 17434 5468
rect 17490 5466 17496 5468
rect 17250 5414 17252 5466
rect 17432 5414 17434 5466
rect 17188 5412 17194 5414
rect 17250 5412 17274 5414
rect 17330 5412 17354 5414
rect 17410 5412 17434 5414
rect 17490 5412 17496 5414
rect 17188 5403 17496 5412
rect 17130 5264 17186 5273
rect 17130 5199 17186 5208
rect 17144 4758 17172 5199
rect 17040 4752 17092 4758
rect 17038 4720 17040 4729
rect 17132 4752 17184 4758
rect 17092 4720 17094 4729
rect 17132 4694 17184 4700
rect 17038 4655 17094 4664
rect 17188 4380 17496 4389
rect 17188 4378 17194 4380
rect 17250 4378 17274 4380
rect 17330 4378 17354 4380
rect 17410 4378 17434 4380
rect 17490 4378 17496 4380
rect 17250 4326 17252 4378
rect 17432 4326 17434 4378
rect 17188 4324 17194 4326
rect 17250 4324 17274 4326
rect 17330 4324 17354 4326
rect 17410 4324 17434 4326
rect 17490 4324 17496 4326
rect 17188 4315 17496 4324
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 16948 4208 17000 4214
rect 16948 4150 17000 4156
rect 17052 4078 17080 4218
rect 17316 4208 17368 4214
rect 17316 4150 17368 4156
rect 17684 4208 17736 4214
rect 17684 4150 17736 4156
rect 17328 4078 17356 4150
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17052 3670 17080 4014
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16856 3528 16908 3534
rect 16960 3505 16988 3538
rect 17696 3534 17724 4150
rect 17788 3670 17816 6870
rect 18064 6254 18092 7414
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 17960 6112 18012 6118
rect 17960 6054 18012 6060
rect 17972 5234 18000 6054
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18064 5370 18092 5714
rect 18156 5574 18184 6258
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 18156 5302 18184 5510
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18064 3670 18092 3878
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 18052 3664 18104 3670
rect 18052 3606 18104 3612
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17684 3528 17736 3534
rect 16856 3470 16908 3476
rect 16946 3496 17002 3505
rect 16672 3460 16724 3466
rect 17684 3470 17736 3476
rect 16946 3431 17002 3440
rect 16672 3402 16724 3408
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16488 2984 16540 2990
rect 16408 2944 16488 2972
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 16120 2916 16172 2922
rect 16120 2858 16172 2864
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 15934 2000 15990 2009
rect 15934 1935 15990 1944
rect 15948 1902 15976 1935
rect 16132 1902 16160 2246
rect 15936 1896 15988 1902
rect 15936 1838 15988 1844
rect 16120 1896 16172 1902
rect 16120 1838 16172 1844
rect 15844 1760 15896 1766
rect 15844 1702 15896 1708
rect 16224 1562 16252 2586
rect 16408 1834 16436 2944
rect 16488 2926 16540 2932
rect 16684 2922 16712 3402
rect 16960 3194 16988 3431
rect 17188 3292 17496 3301
rect 17188 3290 17194 3292
rect 17250 3290 17274 3292
rect 17330 3290 17354 3292
rect 17410 3290 17434 3292
rect 17490 3290 17496 3292
rect 17250 3238 17252 3290
rect 17432 3238 17434 3290
rect 17188 3236 17194 3238
rect 17250 3236 17274 3238
rect 17330 3236 17354 3238
rect 17410 3236 17434 3238
rect 17490 3236 17496 3238
rect 17188 3227 17496 3236
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16776 2990 16804 3130
rect 17972 3097 18000 3538
rect 18156 3534 18184 5238
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 17958 3088 18014 3097
rect 18156 3058 18184 3470
rect 18144 3052 18196 3058
rect 17958 3023 18014 3032
rect 18064 3012 18144 3040
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 16488 2848 16540 2854
rect 16488 2790 16540 2796
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16500 2514 16528 2790
rect 16960 2514 16988 2790
rect 16488 2508 16540 2514
rect 16488 2450 16540 2456
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17188 2204 17496 2213
rect 17188 2202 17194 2204
rect 17250 2202 17274 2204
rect 17330 2202 17354 2204
rect 17410 2202 17434 2204
rect 17490 2202 17496 2204
rect 17250 2150 17252 2202
rect 17432 2150 17434 2202
rect 17188 2148 17194 2150
rect 17250 2148 17274 2150
rect 17330 2148 17354 2150
rect 17410 2148 17434 2150
rect 17490 2148 17496 2150
rect 17188 2139 17496 2148
rect 16580 2032 16632 2038
rect 16580 1974 16632 1980
rect 16396 1828 16448 1834
rect 16396 1770 16448 1776
rect 16408 1562 16436 1770
rect 16212 1556 16264 1562
rect 16212 1498 16264 1504
rect 16396 1556 16448 1562
rect 16396 1498 16448 1504
rect 15568 1420 15620 1426
rect 15568 1362 15620 1368
rect 15580 1222 15608 1362
rect 15568 1216 15620 1222
rect 15568 1158 15620 1164
rect 14740 944 14792 950
rect 14740 886 14792 892
rect 14832 944 14884 950
rect 14832 886 14884 892
rect 14752 814 14780 886
rect 14372 808 14424 814
rect 14372 750 14424 756
rect 14740 808 14792 814
rect 14740 750 14792 756
rect 13912 740 13964 746
rect 13912 682 13964 688
rect 13830 572 14138 581
rect 13830 570 13836 572
rect 13892 570 13916 572
rect 13972 570 13996 572
rect 14052 570 14076 572
rect 14132 570 14138 572
rect 13892 518 13894 570
rect 14074 518 14076 570
rect 13830 516 13836 518
rect 13892 516 13916 518
rect 13972 516 13996 518
rect 14052 516 14076 518
rect 14132 516 14138 518
rect 13830 507 14138 516
rect 14844 400 14872 886
rect 15580 882 15608 1158
rect 15568 876 15620 882
rect 15568 818 15620 824
rect 16592 400 16620 1974
rect 17604 1494 17632 2246
rect 17788 1902 17816 2246
rect 17958 2000 18014 2009
rect 17958 1935 18014 1944
rect 17776 1896 17828 1902
rect 17776 1838 17828 1844
rect 17868 1760 17920 1766
rect 17868 1702 17920 1708
rect 17592 1488 17644 1494
rect 17592 1430 17644 1436
rect 17880 1358 17908 1702
rect 17972 1562 18000 1935
rect 18064 1902 18092 3012
rect 18144 2994 18196 3000
rect 18248 2774 18276 7346
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18340 6254 18368 6598
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18432 5846 18460 6190
rect 18420 5840 18472 5846
rect 18420 5782 18472 5788
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18340 2990 18368 3334
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18156 2746 18276 2774
rect 18156 1902 18184 2746
rect 18052 1896 18104 1902
rect 18052 1838 18104 1844
rect 18144 1896 18196 1902
rect 18144 1838 18196 1844
rect 17960 1556 18012 1562
rect 17960 1498 18012 1504
rect 17972 1426 18000 1498
rect 17960 1420 18012 1426
rect 17960 1362 18012 1368
rect 17868 1352 17920 1358
rect 17868 1294 17920 1300
rect 18064 1290 18092 1838
rect 18156 1426 18184 1838
rect 18524 1562 18552 16730
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18800 15706 18828 15982
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18708 15162 18736 15506
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18616 14958 18644 15098
rect 18800 15026 18828 15642
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18788 14068 18840 14074
rect 18708 14028 18788 14056
rect 18708 13394 18736 14028
rect 18788 14010 18840 14016
rect 18788 13728 18840 13734
rect 18788 13670 18840 13676
rect 18800 13462 18828 13670
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18616 12986 18644 13330
rect 18708 13190 18736 13330
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18602 12336 18658 12345
rect 18658 12280 18828 12288
rect 18602 12271 18604 12280
rect 18656 12260 18828 12280
rect 18604 12242 18656 12248
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18616 10810 18644 11154
rect 18800 11150 18828 12260
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18892 10470 18920 15574
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19076 14278 19104 14894
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 19064 10532 19116 10538
rect 19064 10474 19116 10480
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 19076 10266 19104 10474
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 19076 10169 19104 10202
rect 18602 10160 18658 10169
rect 19062 10160 19118 10169
rect 18602 10095 18604 10104
rect 18656 10095 18658 10104
rect 18880 10124 18932 10130
rect 18604 10066 18656 10072
rect 19062 10095 19064 10104
rect 18880 10066 18932 10072
rect 19116 10095 19118 10104
rect 19064 10066 19116 10072
rect 18892 9926 18920 10066
rect 18880 9920 18932 9926
rect 18880 9862 18932 9868
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18616 7954 18644 8230
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18708 7818 18736 8910
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18800 8090 18828 8298
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18708 6338 18736 7754
rect 18984 7546 19012 9454
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19076 9178 19104 9318
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 19168 7562 19196 16730
rect 19536 16658 19564 17002
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 19616 16720 19668 16726
rect 19616 16662 19668 16668
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19352 15094 19380 15846
rect 19444 15638 19472 15846
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 19430 14920 19486 14929
rect 19430 14855 19486 14864
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19246 13560 19302 13569
rect 19246 13495 19302 13504
rect 19260 13394 19288 13495
rect 19352 13394 19380 14758
rect 19444 13802 19472 14855
rect 19536 14618 19564 14962
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 19260 12238 19288 12854
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19260 11218 19288 12174
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 18972 7540 19024 7546
rect 19168 7534 19288 7562
rect 18972 7482 19024 7488
rect 18616 6310 18736 6338
rect 18616 6254 18644 6310
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18616 4214 18644 4558
rect 18604 4208 18656 4214
rect 18604 4150 18656 4156
rect 19064 1964 19116 1970
rect 19064 1906 19116 1912
rect 19076 1562 19104 1906
rect 19168 1902 19196 4966
rect 19156 1896 19208 1902
rect 19156 1838 19208 1844
rect 18512 1556 18564 1562
rect 18512 1498 18564 1504
rect 19064 1556 19116 1562
rect 19064 1498 19116 1504
rect 19260 1465 19288 7534
rect 19352 7410 19380 10066
rect 19444 9654 19472 13262
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19536 11354 19564 12242
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19628 10146 19656 16662
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 19720 13734 19748 13806
rect 19708 13728 19760 13734
rect 19708 13670 19760 13676
rect 19812 12434 19840 16934
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 19892 15564 19944 15570
rect 19892 15506 19944 15512
rect 19904 14958 19932 15506
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19904 13530 19932 14350
rect 19892 13524 19944 13530
rect 19892 13466 19944 13472
rect 19996 13410 20024 16730
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20088 14618 20116 15982
rect 20272 15706 20300 15982
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20168 15564 20220 15570
rect 20168 15506 20220 15512
rect 20180 14618 20208 15506
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20168 14476 20220 14482
rect 20272 14464 20300 14894
rect 20220 14436 20300 14464
rect 20168 14418 20220 14424
rect 20180 13870 20208 14418
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20364 13433 20392 16934
rect 20546 16892 20854 16901
rect 20546 16890 20552 16892
rect 20608 16890 20632 16892
rect 20688 16890 20712 16892
rect 20768 16890 20792 16892
rect 20848 16890 20854 16892
rect 20608 16838 20610 16890
rect 20790 16838 20792 16890
rect 20546 16836 20552 16838
rect 20608 16836 20632 16838
rect 20688 16836 20712 16838
rect 20768 16836 20792 16838
rect 20848 16836 20854 16838
rect 20546 16827 20854 16836
rect 21468 16522 21496 16934
rect 21548 16788 21600 16794
rect 21548 16730 21600 16736
rect 21456 16516 21508 16522
rect 21456 16458 21508 16464
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 20546 15804 20854 15813
rect 20546 15802 20552 15804
rect 20608 15802 20632 15804
rect 20688 15802 20712 15804
rect 20768 15802 20792 15804
rect 20848 15802 20854 15804
rect 20608 15750 20610 15802
rect 20790 15750 20792 15802
rect 20546 15748 20552 15750
rect 20608 15748 20632 15750
rect 20688 15748 20712 15750
rect 20768 15748 20792 15750
rect 20848 15748 20854 15750
rect 20546 15739 20854 15748
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 20456 14482 20484 15438
rect 20916 15026 20944 15846
rect 21100 15570 21128 15846
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20812 14952 20864 14958
rect 20810 14920 20812 14929
rect 20864 14920 20866 14929
rect 20810 14855 20866 14864
rect 20546 14716 20854 14725
rect 20546 14714 20552 14716
rect 20608 14714 20632 14716
rect 20688 14714 20712 14716
rect 20768 14714 20792 14716
rect 20848 14714 20854 14716
rect 20608 14662 20610 14714
rect 20790 14662 20792 14714
rect 20546 14660 20552 14662
rect 20608 14660 20632 14662
rect 20688 14660 20712 14662
rect 20768 14660 20792 14662
rect 20848 14660 20854 14662
rect 20546 14651 20854 14660
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20732 14482 20760 14554
rect 20916 14550 20944 14962
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 21192 14550 21220 14826
rect 21560 14600 21588 16730
rect 21744 16590 21772 16934
rect 21732 16584 21784 16590
rect 21732 16526 21784 16532
rect 22756 16522 22784 16934
rect 22744 16516 22796 16522
rect 22744 16458 22796 16464
rect 24044 16454 24072 16934
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 23904 16348 24212 16357
rect 23904 16346 23910 16348
rect 23966 16346 23990 16348
rect 24046 16346 24070 16348
rect 24126 16346 24150 16348
rect 24206 16346 24212 16348
rect 23966 16294 23968 16346
rect 24148 16294 24150 16346
rect 23904 16292 23910 16294
rect 23966 16292 23990 16294
rect 24046 16292 24070 16294
rect 24126 16292 24150 16294
rect 24206 16292 24212 16294
rect 23904 16283 24212 16292
rect 24688 16250 24716 16934
rect 24872 16658 24900 16934
rect 25792 16794 25820 17070
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24780 16538 24808 16594
rect 25320 16584 25372 16590
rect 24780 16510 24992 16538
rect 25320 16526 25372 16532
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 23940 16108 23992 16114
rect 23940 16050 23992 16056
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21744 15366 21772 15982
rect 22836 15700 22888 15706
rect 22836 15642 22888 15648
rect 22652 15632 22704 15638
rect 22848 15609 22876 15642
rect 22652 15574 22704 15580
rect 22834 15600 22890 15609
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 21732 15360 21784 15366
rect 21784 15320 21864 15348
rect 21732 15302 21784 15308
rect 21468 14572 21588 14600
rect 20904 14544 20956 14550
rect 20904 14486 20956 14492
rect 21180 14544 21232 14550
rect 21180 14486 21232 14492
rect 20444 14476 20496 14482
rect 20444 14418 20496 14424
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 21008 13802 21036 14418
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20546 13628 20854 13637
rect 20546 13626 20552 13628
rect 20608 13626 20632 13628
rect 20688 13626 20712 13628
rect 20768 13626 20792 13628
rect 20848 13626 20854 13628
rect 20608 13574 20610 13626
rect 20790 13574 20792 13626
rect 20546 13572 20552 13574
rect 20608 13572 20632 13574
rect 20688 13572 20712 13574
rect 20768 13572 20792 13574
rect 20848 13572 20854 13574
rect 20546 13563 20854 13572
rect 20916 13462 20944 13670
rect 20904 13456 20956 13462
rect 19536 10118 19656 10146
rect 19720 12406 19840 12434
rect 19904 13382 20024 13410
rect 20350 13424 20406 13433
rect 20076 13388 20128 13394
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19536 9160 19564 10118
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 19444 9132 19564 9160
rect 19444 8537 19472 9132
rect 19524 9036 19576 9042
rect 19524 8978 19576 8984
rect 19430 8528 19486 8537
rect 19430 8463 19486 8472
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19352 6866 19380 7346
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19352 6662 19380 6802
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19444 5658 19472 8463
rect 19536 8294 19564 8978
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19536 7954 19564 8230
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19628 7342 19656 9862
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19628 6934 19656 7278
rect 19616 6928 19668 6934
rect 19536 6876 19616 6882
rect 19536 6870 19668 6876
rect 19536 6854 19656 6870
rect 19536 5778 19564 6854
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19628 6458 19656 6734
rect 19720 6662 19748 12406
rect 19800 12368 19852 12374
rect 19800 12310 19852 12316
rect 19812 11218 19840 12310
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19800 10464 19852 10470
rect 19800 10406 19852 10412
rect 19812 9926 19840 10406
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19800 8968 19852 8974
rect 19800 8910 19852 8916
rect 19812 7886 19840 8910
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19904 7562 19932 13382
rect 20076 13330 20128 13336
rect 20168 13388 20220 13394
rect 20220 13348 20300 13376
rect 20904 13398 20956 13404
rect 20350 13359 20406 13368
rect 20628 13388 20680 13394
rect 20168 13330 20220 13336
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19996 11218 20024 13126
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19996 10130 20024 10610
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 20088 9654 20116 13330
rect 20166 12880 20222 12889
rect 20166 12815 20222 12824
rect 20180 11098 20208 12815
rect 20272 12714 20300 13348
rect 20628 13330 20680 13336
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20260 12708 20312 12714
rect 20260 12650 20312 12656
rect 20272 11200 20300 12650
rect 20364 11898 20392 12922
rect 20640 12889 20668 13330
rect 21008 13258 21036 13738
rect 21100 13530 21128 13806
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 20626 12880 20682 12889
rect 20626 12815 20682 12824
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20456 12306 20484 12650
rect 20546 12540 20854 12549
rect 20546 12538 20552 12540
rect 20608 12538 20632 12540
rect 20688 12538 20712 12540
rect 20768 12538 20792 12540
rect 20848 12538 20854 12540
rect 20608 12486 20610 12538
rect 20790 12486 20792 12538
rect 20546 12484 20552 12486
rect 20608 12484 20632 12486
rect 20688 12484 20712 12486
rect 20768 12484 20792 12486
rect 20848 12484 20854 12486
rect 20546 12475 20854 12484
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20272 11172 20392 11200
rect 20180 11070 20300 11098
rect 20364 11082 20392 11172
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 20180 10742 20208 10950
rect 20168 10736 20220 10742
rect 20168 10678 20220 10684
rect 20168 10600 20220 10606
rect 20272 10588 20300 11070
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20220 10560 20300 10588
rect 20352 10600 20404 10606
rect 20168 10542 20220 10548
rect 20352 10542 20404 10548
rect 20180 10130 20208 10542
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20168 10124 20220 10130
rect 20168 10066 20220 10072
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 20076 9104 20128 9110
rect 20076 9046 20128 9052
rect 20088 8634 20116 9046
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 20088 7954 20116 8570
rect 20180 8498 20208 10066
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20180 8090 20208 8434
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 19800 7540 19852 7546
rect 19904 7534 20208 7562
rect 19800 7482 19852 7488
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19444 5630 19748 5658
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19524 4548 19576 4554
rect 19524 4490 19576 4496
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19352 4078 19380 4422
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19444 2990 19472 3878
rect 19536 3738 19564 4490
rect 19628 4282 19656 4762
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19246 1456 19302 1465
rect 18144 1420 18196 1426
rect 19536 1442 19564 3674
rect 19720 2774 19748 5630
rect 19812 3602 19840 7482
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 20088 6866 20116 7142
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 19892 5908 19944 5914
rect 19892 5850 19944 5856
rect 19904 5166 19932 5850
rect 19996 5778 20024 6326
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19892 5160 19944 5166
rect 19892 5102 19944 5108
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19892 3664 19944 3670
rect 19892 3606 19944 3612
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 19720 2746 19840 2774
rect 19812 2666 19840 2746
rect 19720 2638 19840 2666
rect 19720 1902 19748 2638
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 19708 1896 19760 1902
rect 19708 1838 19760 1844
rect 19352 1426 19564 1442
rect 19246 1391 19248 1400
rect 18144 1362 18196 1368
rect 19300 1391 19302 1400
rect 19340 1420 19564 1426
rect 19248 1362 19300 1368
rect 19392 1414 19564 1420
rect 19340 1362 19392 1368
rect 18052 1284 18104 1290
rect 18052 1226 18104 1232
rect 18328 1216 18380 1222
rect 18328 1158 18380 1164
rect 17188 1116 17496 1125
rect 17188 1114 17194 1116
rect 17250 1114 17274 1116
rect 17330 1114 17354 1116
rect 17410 1114 17434 1116
rect 17490 1114 17496 1116
rect 17250 1062 17252 1114
rect 17432 1062 17434 1114
rect 17188 1060 17194 1062
rect 17250 1060 17274 1062
rect 17330 1060 17354 1062
rect 17410 1060 17434 1062
rect 17490 1060 17496 1062
rect 17188 1051 17496 1060
rect 18340 400 18368 1158
rect 19720 678 19748 1838
rect 19812 1834 19840 2450
rect 19800 1828 19852 1834
rect 19800 1770 19852 1776
rect 19812 1426 19840 1770
rect 19904 1426 19932 3606
rect 19996 2514 20024 4218
rect 20088 2650 20116 6598
rect 20180 2774 20208 7534
rect 20272 7002 20300 10406
rect 20364 10130 20392 10542
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20456 9722 20484 12242
rect 20546 11452 20854 11461
rect 20546 11450 20552 11452
rect 20608 11450 20632 11452
rect 20688 11450 20712 11452
rect 20768 11450 20792 11452
rect 20848 11450 20854 11452
rect 20608 11398 20610 11450
rect 20790 11398 20792 11450
rect 20546 11396 20552 11398
rect 20608 11396 20632 11398
rect 20688 11396 20712 11398
rect 20768 11396 20792 11398
rect 20848 11396 20854 11398
rect 20546 11387 20854 11396
rect 21008 11354 21036 13194
rect 21192 12646 21220 13262
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 21100 11218 21128 11834
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 21088 11212 21140 11218
rect 21088 11154 21140 11160
rect 20548 11082 20576 11154
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20548 10674 20576 11018
rect 20824 10810 20852 11086
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 21192 10690 21220 12582
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21284 11218 21312 11698
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 21008 10662 21220 10690
rect 21008 10606 21036 10662
rect 20996 10600 21048 10606
rect 20996 10542 21048 10548
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 20546 10364 20854 10373
rect 20546 10362 20552 10364
rect 20608 10362 20632 10364
rect 20688 10362 20712 10364
rect 20768 10362 20792 10364
rect 20848 10362 20854 10364
rect 20608 10310 20610 10362
rect 20790 10310 20792 10362
rect 20546 10308 20552 10310
rect 20608 10308 20632 10310
rect 20688 10308 20712 10310
rect 20768 10308 20792 10310
rect 20848 10308 20854 10310
rect 20546 10299 20854 10308
rect 21100 10266 21128 10542
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20364 8634 20392 9318
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20352 7268 20404 7274
rect 20352 7210 20404 7216
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20272 5778 20300 6598
rect 20364 5914 20392 7210
rect 20456 6798 20484 9658
rect 20824 9382 20852 10066
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20546 9276 20854 9285
rect 20546 9274 20552 9276
rect 20608 9274 20632 9276
rect 20688 9274 20712 9276
rect 20768 9274 20792 9276
rect 20848 9274 20854 9276
rect 20608 9222 20610 9274
rect 20790 9222 20792 9274
rect 20546 9220 20552 9222
rect 20608 9220 20632 9222
rect 20688 9220 20712 9222
rect 20768 9220 20792 9222
rect 20848 9220 20854 9222
rect 20546 9211 20854 9220
rect 20916 9178 20944 9318
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20546 8188 20854 8197
rect 20546 8186 20552 8188
rect 20608 8186 20632 8188
rect 20688 8186 20712 8188
rect 20768 8186 20792 8188
rect 20848 8186 20854 8188
rect 20608 8134 20610 8186
rect 20790 8134 20792 8186
rect 20546 8132 20552 8134
rect 20608 8132 20632 8134
rect 20688 8132 20712 8134
rect 20768 8132 20792 8134
rect 20848 8132 20854 8134
rect 20546 8123 20854 8132
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20548 7206 20576 8026
rect 20812 8016 20864 8022
rect 20916 8004 20944 9114
rect 20864 7976 20944 8004
rect 20812 7958 20864 7964
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 20640 7721 20668 7754
rect 20626 7712 20682 7721
rect 20626 7647 20682 7656
rect 20536 7200 20588 7206
rect 20536 7142 20588 7148
rect 20546 7100 20854 7109
rect 20546 7098 20552 7100
rect 20608 7098 20632 7100
rect 20688 7098 20712 7100
rect 20768 7098 20792 7100
rect 20848 7098 20854 7100
rect 20608 7046 20610 7098
rect 20790 7046 20792 7098
rect 20546 7044 20552 7046
rect 20608 7044 20632 7046
rect 20688 7044 20712 7046
rect 20768 7044 20792 7046
rect 20848 7044 20854 7046
rect 20546 7035 20854 7044
rect 21008 7018 21036 10202
rect 21088 8356 21140 8362
rect 21088 8298 21140 8304
rect 21100 7886 21128 8298
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 21192 7546 21220 10662
rect 21364 10192 21416 10198
rect 21364 10134 21416 10140
rect 21376 9518 21404 10134
rect 21364 9512 21416 9518
rect 21364 9454 21416 9460
rect 21468 9466 21496 14572
rect 21836 14482 21864 15320
rect 21914 14920 21970 14929
rect 21914 14855 21970 14864
rect 22008 14884 22060 14890
rect 21928 14482 21956 14855
rect 22008 14826 22060 14832
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 21916 14476 21968 14482
rect 21916 14418 21968 14424
rect 21560 14006 21588 14418
rect 22020 14414 22048 14826
rect 22572 14618 22600 15506
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 21652 14074 21680 14350
rect 22296 14074 22324 14350
rect 21640 14068 21692 14074
rect 21640 14010 21692 14016
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 21548 14000 21600 14006
rect 21548 13942 21600 13948
rect 21560 13530 21588 13942
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 22204 13462 22232 13670
rect 22192 13456 22244 13462
rect 22192 13398 22244 13404
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22100 12776 22152 12782
rect 21836 12736 22100 12764
rect 21836 12646 21864 12736
rect 22100 12718 22152 12724
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 21928 12238 21956 12582
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 21640 11620 21692 11626
rect 21640 11562 21692 11568
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21560 10810 21588 11154
rect 21652 10810 21680 11562
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21640 10804 21692 10810
rect 21640 10746 21692 10752
rect 22204 10674 22232 11222
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 22112 10470 22140 10610
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22296 10266 22324 12718
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 22388 10606 22416 10950
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21732 10124 21784 10130
rect 21732 10066 21784 10072
rect 21468 9438 21588 9466
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21468 9042 21496 9318
rect 21456 9036 21508 9042
rect 21456 8978 21508 8984
rect 21362 8936 21418 8945
rect 21362 8871 21418 8880
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20916 6990 21220 7018
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20456 6254 20484 6734
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20640 6118 20668 6938
rect 20916 6866 20944 6990
rect 20996 6928 21048 6934
rect 20996 6870 21048 6876
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20824 6254 20852 6802
rect 20904 6384 20956 6390
rect 20904 6326 20956 6332
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20546 6012 20854 6021
rect 20546 6010 20552 6012
rect 20608 6010 20632 6012
rect 20688 6010 20712 6012
rect 20768 6010 20792 6012
rect 20848 6010 20854 6012
rect 20608 5958 20610 6010
rect 20790 5958 20792 6010
rect 20546 5956 20552 5958
rect 20608 5956 20632 5958
rect 20688 5956 20712 5958
rect 20768 5956 20792 5958
rect 20848 5956 20854 5958
rect 20546 5947 20854 5956
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20916 5386 20944 6326
rect 21008 6202 21036 6870
rect 21008 6186 21128 6202
rect 21008 6180 21140 6186
rect 21008 6174 21088 6180
rect 21008 5642 21036 6174
rect 21088 6122 21140 6128
rect 21192 5914 21220 6990
rect 21284 6458 21312 8774
rect 21376 8294 21404 8871
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21376 7954 21404 8230
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 21376 6474 21404 7142
rect 21272 6452 21324 6458
rect 21376 6446 21496 6474
rect 21272 6394 21324 6400
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21284 6186 21312 6258
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 21272 6180 21324 6186
rect 21272 6122 21324 6128
rect 21376 5914 21404 6190
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21192 5710 21220 5850
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 20996 5636 21048 5642
rect 20996 5578 21048 5584
rect 21468 5574 21496 6446
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 20824 5370 20944 5386
rect 20812 5364 20944 5370
rect 20864 5358 20944 5364
rect 20812 5306 20864 5312
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 20546 4924 20854 4933
rect 20546 4922 20552 4924
rect 20608 4922 20632 4924
rect 20688 4922 20712 4924
rect 20768 4922 20792 4924
rect 20848 4922 20854 4924
rect 20608 4870 20610 4922
rect 20790 4870 20792 4922
rect 20546 4868 20552 4870
rect 20608 4868 20632 4870
rect 20688 4868 20712 4870
rect 20768 4868 20792 4870
rect 20848 4868 20854 4870
rect 20546 4859 20854 4868
rect 21008 4146 21036 5102
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20546 3836 20854 3845
rect 20546 3834 20552 3836
rect 20608 3834 20632 3836
rect 20688 3834 20712 3836
rect 20768 3834 20792 3836
rect 20848 3834 20854 3836
rect 20608 3782 20610 3834
rect 20790 3782 20792 3834
rect 20546 3780 20552 3782
rect 20608 3780 20632 3782
rect 20688 3780 20712 3782
rect 20768 3780 20792 3782
rect 20848 3780 20854 3782
rect 20546 3771 20854 3780
rect 21008 3602 21036 4082
rect 20444 3596 20496 3602
rect 20444 3538 20496 3544
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 20456 3194 20484 3538
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20364 3040 20392 3130
rect 20364 3012 20484 3040
rect 20180 2746 20392 2774
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20088 2514 20116 2586
rect 20364 2553 20392 2746
rect 20350 2544 20406 2553
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 20076 2508 20128 2514
rect 20350 2479 20406 2488
rect 20076 2450 20128 2456
rect 20456 1902 20484 3012
rect 21560 2774 21588 9438
rect 21652 9178 21680 10066
rect 21744 9994 21772 10066
rect 21732 9988 21784 9994
rect 21732 9930 21784 9936
rect 22480 9674 22508 13126
rect 22664 11354 22692 15574
rect 23952 15570 23980 16050
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 22834 15535 22890 15544
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 22744 15360 22796 15366
rect 22744 15302 22796 15308
rect 22756 13870 22784 15302
rect 22940 14521 22968 15506
rect 23124 14550 23152 15506
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 23112 14544 23164 14550
rect 22926 14512 22982 14521
rect 23112 14486 23164 14492
rect 23216 14482 23244 14758
rect 23400 14482 23428 15506
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23492 15026 23520 15438
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 22926 14447 22928 14456
rect 22980 14447 22982 14456
rect 23020 14476 23072 14482
rect 22928 14418 22980 14424
rect 23020 14418 23072 14424
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22848 13938 22876 14214
rect 22836 13932 22888 13938
rect 22836 13874 22888 13880
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22928 13524 22980 13530
rect 22928 13466 22980 13472
rect 22940 13394 22968 13466
rect 22928 13388 22980 13394
rect 22928 13330 22980 13336
rect 22940 12434 22968 13330
rect 23032 12986 23060 14418
rect 23216 14074 23244 14418
rect 23400 14074 23428 14418
rect 23204 14068 23256 14074
rect 23204 14010 23256 14016
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23032 12782 23060 12922
rect 23400 12782 23428 14010
rect 23584 13530 23612 15506
rect 23904 15260 24212 15269
rect 23904 15258 23910 15260
rect 23966 15258 23990 15260
rect 24046 15258 24070 15260
rect 24126 15258 24150 15260
rect 24206 15258 24212 15260
rect 23966 15206 23968 15258
rect 24148 15206 24150 15258
rect 23904 15204 23910 15206
rect 23966 15204 23990 15206
rect 24046 15204 24070 15206
rect 24126 15204 24150 15206
rect 24206 15204 24212 15206
rect 23904 15195 24212 15204
rect 24032 15088 24084 15094
rect 24032 15030 24084 15036
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23676 14346 23704 14486
rect 24044 14482 24072 15030
rect 24412 14482 24440 15846
rect 24504 15706 24532 15982
rect 24964 15910 24992 16510
rect 25228 16448 25280 16454
rect 25228 16390 25280 16396
rect 24952 15904 25004 15910
rect 24952 15846 25004 15852
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 24504 15162 24532 15642
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24676 15360 24728 15366
rect 24676 15302 24728 15308
rect 24492 15156 24544 15162
rect 24492 15098 24544 15104
rect 24688 14958 24716 15302
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 23756 14476 23808 14482
rect 23756 14418 23808 14424
rect 24032 14476 24084 14482
rect 24032 14418 24084 14424
rect 24400 14476 24452 14482
rect 24400 14418 24452 14424
rect 23664 14340 23716 14346
rect 23664 14282 23716 14288
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23676 12850 23704 14282
rect 23768 13870 23796 14418
rect 24584 14272 24636 14278
rect 24584 14214 24636 14220
rect 23904 14172 24212 14181
rect 23904 14170 23910 14172
rect 23966 14170 23990 14172
rect 24046 14170 24070 14172
rect 24126 14170 24150 14172
rect 24206 14170 24212 14172
rect 23966 14118 23968 14170
rect 24148 14118 24150 14170
rect 23904 14116 23910 14118
rect 23966 14116 23990 14118
rect 24046 14116 24070 14118
rect 24126 14116 24150 14118
rect 24206 14116 24212 14118
rect 23904 14107 24212 14116
rect 24596 14006 24624 14214
rect 24584 14000 24636 14006
rect 24584 13942 24636 13948
rect 24688 13870 24716 14894
rect 24872 14618 24900 15506
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24964 14482 24992 15846
rect 25240 15638 25268 16390
rect 25332 16046 25360 16526
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25320 16040 25372 16046
rect 25320 15982 25372 15988
rect 25228 15632 25280 15638
rect 25228 15574 25280 15580
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 24768 14408 24820 14414
rect 24964 14362 24992 14418
rect 24820 14356 24992 14362
rect 24768 14350 24992 14356
rect 24780 14334 24992 14350
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 24584 13864 24636 13870
rect 24584 13806 24636 13812
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 23860 13394 23888 13670
rect 24596 13530 24624 13806
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24688 13394 24716 13806
rect 24872 13462 24900 13874
rect 24860 13456 24912 13462
rect 24860 13398 24912 13404
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24688 13274 24716 13330
rect 24964 13274 24992 14334
rect 24688 13246 24808 13274
rect 23904 13084 24212 13093
rect 23904 13082 23910 13084
rect 23966 13082 23990 13084
rect 24046 13082 24070 13084
rect 24126 13082 24150 13084
rect 24206 13082 24212 13084
rect 23966 13030 23968 13082
rect 24148 13030 24150 13082
rect 23904 13028 23910 13030
rect 23966 13028 23990 13030
rect 24046 13028 24070 13030
rect 24126 13028 24150 13030
rect 24206 13028 24212 13030
rect 23904 13019 24212 13028
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 23388 12776 23440 12782
rect 24308 12776 24360 12782
rect 23388 12718 23440 12724
rect 24306 12744 24308 12753
rect 24492 12776 24544 12782
rect 24360 12744 24362 12753
rect 24492 12718 24544 12724
rect 24676 12776 24728 12782
rect 24676 12718 24728 12724
rect 24306 12679 24362 12688
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 22940 12406 23060 12434
rect 23032 12102 23060 12406
rect 24412 12238 24440 12582
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22928 10600 22980 10606
rect 22928 10542 22980 10548
rect 22836 10532 22888 10538
rect 22836 10474 22888 10480
rect 22848 10130 22876 10474
rect 22940 10266 22968 10542
rect 22928 10260 22980 10266
rect 22928 10202 22980 10208
rect 22836 10124 22888 10130
rect 22836 10066 22888 10072
rect 22296 9646 22508 9674
rect 21732 9444 21784 9450
rect 21732 9386 21784 9392
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21652 7993 21680 8910
rect 21744 8634 21772 9386
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21744 8498 21772 8570
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21638 7984 21694 7993
rect 21638 7919 21640 7928
rect 21692 7919 21694 7928
rect 21640 7890 21692 7896
rect 21836 7274 21864 8366
rect 22008 8356 22060 8362
rect 22008 8298 22060 8304
rect 22020 8022 22048 8298
rect 22008 8016 22060 8022
rect 22008 7958 22060 7964
rect 22008 7744 22060 7750
rect 22296 7721 22324 9646
rect 22928 9376 22980 9382
rect 22928 9318 22980 9324
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22480 8498 22508 8774
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22468 8356 22520 8362
rect 22468 8298 22520 8304
rect 22480 7818 22508 8298
rect 22572 7954 22600 8570
rect 22652 8424 22704 8430
rect 22652 8366 22704 8372
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22664 7886 22692 8366
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22008 7686 22060 7692
rect 22282 7712 22338 7721
rect 22020 7342 22048 7686
rect 22282 7647 22338 7656
rect 22834 7712 22890 7721
rect 22834 7647 22890 7656
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 21824 7268 21876 7274
rect 21824 7210 21876 7216
rect 21836 6254 21864 7210
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 22388 6254 22416 6598
rect 21824 6248 21876 6254
rect 21824 6190 21876 6196
rect 22376 6248 22428 6254
rect 22376 6190 22428 6196
rect 21836 5166 21864 6190
rect 22848 6186 22876 7647
rect 22940 7342 22968 9318
rect 22928 7336 22980 7342
rect 22928 7278 22980 7284
rect 22008 6180 22060 6186
rect 22008 6122 22060 6128
rect 22744 6180 22796 6186
rect 22744 6122 22796 6128
rect 22836 6180 22888 6186
rect 22836 6122 22888 6128
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 22020 5658 22048 6122
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22572 5710 22600 6054
rect 22756 5914 22784 6122
rect 22744 5908 22796 5914
rect 22744 5850 22796 5856
rect 22376 5704 22428 5710
rect 22020 5652 22376 5658
rect 22020 5646 22428 5652
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 21928 5522 21956 5646
rect 22020 5630 22416 5646
rect 22100 5568 22152 5574
rect 21928 5516 22100 5522
rect 21928 5510 22152 5516
rect 21928 5494 22140 5510
rect 21928 5370 21956 5494
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 23032 4010 23060 12038
rect 23492 10606 23520 12038
rect 23768 11762 23796 12174
rect 23904 11996 24212 12005
rect 23904 11994 23910 11996
rect 23966 11994 23990 11996
rect 24046 11994 24070 11996
rect 24126 11994 24150 11996
rect 24206 11994 24212 11996
rect 23966 11942 23968 11994
rect 24148 11942 24150 11994
rect 23904 11940 23910 11942
rect 23966 11940 23990 11942
rect 24046 11940 24070 11942
rect 24126 11940 24150 11942
rect 24206 11940 24212 11942
rect 23904 11931 24212 11940
rect 24412 11898 24440 12174
rect 24400 11892 24452 11898
rect 24400 11834 24452 11840
rect 23756 11756 23808 11762
rect 23756 11698 23808 11704
rect 23768 11150 23796 11698
rect 24400 11688 24452 11694
rect 24400 11630 24452 11636
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23664 10192 23716 10198
rect 23664 10134 23716 10140
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 23204 9444 23256 9450
rect 23204 9386 23256 9392
rect 23216 9178 23244 9386
rect 23204 9172 23256 9178
rect 23204 9114 23256 9120
rect 23492 9110 23520 9862
rect 23676 9722 23704 10134
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23768 9586 23796 11086
rect 23904 10908 24212 10917
rect 23904 10906 23910 10908
rect 23966 10906 23990 10908
rect 24046 10906 24070 10908
rect 24126 10906 24150 10908
rect 24206 10906 24212 10908
rect 23966 10854 23968 10906
rect 24148 10854 24150 10906
rect 23904 10852 23910 10854
rect 23966 10852 23990 10854
rect 24046 10852 24070 10854
rect 24126 10852 24150 10854
rect 24206 10852 24212 10854
rect 23904 10843 24212 10852
rect 24412 10810 24440 11630
rect 24504 11014 24532 12718
rect 24492 11008 24544 11014
rect 24492 10950 24544 10956
rect 24400 10804 24452 10810
rect 24400 10746 24452 10752
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24504 10266 24532 10542
rect 24400 10260 24452 10266
rect 24400 10202 24452 10208
rect 24492 10260 24544 10266
rect 24492 10202 24544 10208
rect 24308 10124 24360 10130
rect 24308 10066 24360 10072
rect 23904 9820 24212 9829
rect 23904 9818 23910 9820
rect 23966 9818 23990 9820
rect 24046 9818 24070 9820
rect 24126 9818 24150 9820
rect 24206 9818 24212 9820
rect 23966 9766 23968 9818
rect 24148 9766 24150 9818
rect 23904 9764 23910 9766
rect 23966 9764 23990 9766
rect 24046 9764 24070 9766
rect 24126 9764 24150 9766
rect 24206 9764 24212 9766
rect 23904 9755 24212 9764
rect 23756 9580 23808 9586
rect 23756 9522 23808 9528
rect 23848 9512 23900 9518
rect 23848 9454 23900 9460
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23480 9104 23532 9110
rect 23480 9046 23532 9052
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23664 9036 23716 9042
rect 23664 8978 23716 8984
rect 23400 8566 23428 8978
rect 23480 8900 23532 8906
rect 23480 8842 23532 8848
rect 23492 8786 23520 8842
rect 23492 8758 23612 8786
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23400 8022 23428 8230
rect 23388 8016 23440 8022
rect 23388 7958 23440 7964
rect 23492 7818 23520 8366
rect 23584 7954 23612 8758
rect 23676 8634 23704 8978
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23768 8498 23796 9318
rect 23860 9178 23888 9454
rect 24320 9450 24348 10066
rect 24124 9444 24176 9450
rect 24124 9386 24176 9392
rect 24308 9444 24360 9450
rect 24308 9386 24360 9392
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 24136 9042 24164 9386
rect 24412 9217 24440 10202
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24504 9926 24532 10066
rect 24492 9920 24544 9926
rect 24492 9862 24544 9868
rect 24688 9654 24716 12718
rect 24780 12238 24808 13246
rect 24872 13246 24992 13274
rect 24872 12918 24900 13246
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 24860 12912 24912 12918
rect 24860 12854 24912 12860
rect 24964 12782 24992 13126
rect 25056 12986 25084 14418
rect 25148 14414 25176 14758
rect 25332 14482 25360 15982
rect 25320 14476 25372 14482
rect 25320 14418 25372 14424
rect 25136 14408 25188 14414
rect 25136 14350 25188 14356
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25332 12782 25360 14418
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24952 12776 25004 12782
rect 24952 12718 25004 12724
rect 25320 12776 25372 12782
rect 25320 12718 25372 12724
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24780 11762 24808 12174
rect 24768 11756 24820 11762
rect 24768 11698 24820 11704
rect 24768 11008 24820 11014
rect 24768 10950 24820 10956
rect 24780 10674 24808 10950
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24780 10130 24808 10610
rect 24872 10538 24900 12718
rect 25228 12640 25280 12646
rect 25228 12582 25280 12588
rect 25240 12374 25268 12582
rect 25228 12368 25280 12374
rect 25228 12310 25280 12316
rect 25424 11665 25452 16390
rect 25504 16040 25556 16046
rect 25504 15982 25556 15988
rect 25516 14618 25544 15982
rect 25792 15706 25820 16730
rect 25884 16658 25912 17600
rect 26528 17134 26556 17600
rect 26516 17128 26568 17134
rect 26516 17070 26568 17076
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 25976 16182 26004 16934
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 26700 16652 26752 16658
rect 26700 16594 26752 16600
rect 26240 16584 26292 16590
rect 26240 16526 26292 16532
rect 25964 16176 26016 16182
rect 25964 16118 26016 16124
rect 26056 15904 26108 15910
rect 26056 15846 26108 15852
rect 25780 15700 25832 15706
rect 25780 15642 25832 15648
rect 25780 15360 25832 15366
rect 25780 15302 25832 15308
rect 25792 14890 25820 15302
rect 25964 14952 26016 14958
rect 25964 14894 26016 14900
rect 25780 14884 25832 14890
rect 25780 14826 25832 14832
rect 25872 14816 25924 14822
rect 25872 14758 25924 14764
rect 25504 14612 25556 14618
rect 25504 14554 25556 14560
rect 25502 14512 25558 14521
rect 25502 14447 25504 14456
rect 25556 14447 25558 14456
rect 25778 14512 25834 14521
rect 25778 14447 25834 14456
rect 25504 14418 25556 14424
rect 25688 13728 25740 13734
rect 25688 13670 25740 13676
rect 25700 12782 25728 13670
rect 25792 12782 25820 14447
rect 25884 14346 25912 14758
rect 25872 14340 25924 14346
rect 25872 14282 25924 14288
rect 25872 13796 25924 13802
rect 25872 13738 25924 13744
rect 25884 12918 25912 13738
rect 25976 13530 26004 14894
rect 26068 13870 26096 15846
rect 26252 14618 26280 16526
rect 26240 14612 26292 14618
rect 26240 14554 26292 14560
rect 26332 14544 26384 14550
rect 26332 14486 26384 14492
rect 26056 13864 26108 13870
rect 26238 13832 26294 13841
rect 26056 13806 26108 13812
rect 26160 13790 26238 13818
rect 25964 13524 26016 13530
rect 25964 13466 26016 13472
rect 25872 12912 25924 12918
rect 25872 12854 25924 12860
rect 25688 12776 25740 12782
rect 25780 12776 25832 12782
rect 25688 12718 25740 12724
rect 25778 12744 25780 12753
rect 25832 12744 25834 12753
rect 25778 12679 25834 12688
rect 26160 12345 26188 13790
rect 26238 13767 26294 13776
rect 26344 13410 26372 14486
rect 26436 14482 26464 16594
rect 26608 16040 26660 16046
rect 26608 15982 26660 15988
rect 26620 14482 26648 15982
rect 26712 14482 26740 16594
rect 26804 16114 26832 16934
rect 27068 16720 27120 16726
rect 27068 16662 27120 16668
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 26792 16108 26844 16114
rect 26792 16050 26844 16056
rect 26896 14521 26924 16594
rect 26976 16448 27028 16454
rect 26976 16390 27028 16396
rect 26988 15162 27016 16390
rect 26976 15156 27028 15162
rect 26976 15098 27028 15104
rect 26882 14512 26938 14521
rect 26424 14476 26476 14482
rect 26424 14418 26476 14424
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 26700 14476 26752 14482
rect 26700 14418 26752 14424
rect 26792 14476 26844 14482
rect 26882 14447 26884 14456
rect 26792 14418 26844 14424
rect 26936 14447 26938 14456
rect 26884 14418 26936 14424
rect 26436 14074 26464 14418
rect 26516 14272 26568 14278
rect 26516 14214 26568 14220
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26252 13382 26372 13410
rect 26146 12336 26202 12345
rect 26252 12306 26280 13382
rect 26436 12850 26464 14010
rect 26424 12844 26476 12850
rect 26424 12786 26476 12792
rect 26332 12708 26384 12714
rect 26332 12650 26384 12656
rect 26424 12708 26476 12714
rect 26528 12696 26556 14214
rect 26620 14074 26648 14418
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26476 12668 26556 12696
rect 26424 12650 26476 12656
rect 26146 12271 26202 12280
rect 26240 12300 26292 12306
rect 26240 12242 26292 12248
rect 25410 11656 25466 11665
rect 25410 11591 25466 11600
rect 25596 11620 25648 11626
rect 25596 11562 25648 11568
rect 24952 11212 25004 11218
rect 24952 11154 25004 11160
rect 24964 10810 24992 11154
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 25136 11076 25188 11082
rect 25136 11018 25188 11024
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 25148 10606 25176 11018
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 24860 10532 24912 10538
rect 24860 10474 24912 10480
rect 25136 10464 25188 10470
rect 25136 10406 25188 10412
rect 25228 10464 25280 10470
rect 25228 10406 25280 10412
rect 25148 10130 25176 10406
rect 25240 10130 25268 10406
rect 25332 10198 25360 11086
rect 25608 10266 25636 11562
rect 26344 11506 26372 12650
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 26436 11898 26464 12174
rect 26424 11892 26476 11898
rect 26424 11834 26476 11840
rect 26252 11478 26372 11506
rect 26252 11354 26280 11478
rect 26240 11348 26292 11354
rect 26240 11290 26292 11296
rect 26252 11218 26280 11290
rect 26240 11212 26292 11218
rect 26240 11154 26292 11160
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25792 10538 25820 10950
rect 26804 10674 26832 14418
rect 27080 13394 27108 16662
rect 27172 13841 27200 17600
rect 27262 16892 27570 16901
rect 27262 16890 27268 16892
rect 27324 16890 27348 16892
rect 27404 16890 27428 16892
rect 27484 16890 27508 16892
rect 27564 16890 27570 16892
rect 27324 16838 27326 16890
rect 27506 16838 27508 16890
rect 27262 16836 27268 16838
rect 27324 16836 27348 16838
rect 27404 16836 27428 16838
rect 27484 16836 27508 16838
rect 27564 16836 27570 16838
rect 27262 16827 27570 16836
rect 27262 15804 27570 15813
rect 27262 15802 27268 15804
rect 27324 15802 27348 15804
rect 27404 15802 27428 15804
rect 27484 15802 27508 15804
rect 27564 15802 27570 15804
rect 27324 15750 27326 15802
rect 27506 15750 27508 15802
rect 27262 15748 27268 15750
rect 27324 15748 27348 15750
rect 27404 15748 27428 15750
rect 27484 15748 27508 15750
rect 27564 15748 27570 15750
rect 27262 15739 27570 15748
rect 27262 14716 27570 14725
rect 27262 14714 27268 14716
rect 27324 14714 27348 14716
rect 27404 14714 27428 14716
rect 27484 14714 27508 14716
rect 27564 14714 27570 14716
rect 27324 14662 27326 14714
rect 27506 14662 27508 14714
rect 27262 14660 27268 14662
rect 27324 14660 27348 14662
rect 27404 14660 27428 14662
rect 27484 14660 27508 14662
rect 27564 14660 27570 14662
rect 27262 14651 27570 14660
rect 27158 13832 27214 13841
rect 27158 13767 27214 13776
rect 27262 13628 27570 13637
rect 27262 13626 27268 13628
rect 27324 13626 27348 13628
rect 27404 13626 27428 13628
rect 27484 13626 27508 13628
rect 27564 13626 27570 13628
rect 27324 13574 27326 13626
rect 27506 13574 27508 13626
rect 27262 13572 27268 13574
rect 27324 13572 27348 13574
rect 27404 13572 27428 13574
rect 27484 13572 27508 13574
rect 27564 13572 27570 13574
rect 27262 13563 27570 13572
rect 27068 13388 27120 13394
rect 27068 13330 27120 13336
rect 27080 12442 27108 13330
rect 27262 12540 27570 12549
rect 27262 12538 27268 12540
rect 27324 12538 27348 12540
rect 27404 12538 27428 12540
rect 27484 12538 27508 12540
rect 27564 12538 27570 12540
rect 27324 12486 27326 12538
rect 27506 12486 27508 12538
rect 27262 12484 27268 12486
rect 27324 12484 27348 12486
rect 27404 12484 27428 12486
rect 27484 12484 27508 12486
rect 27564 12484 27570 12486
rect 27262 12475 27570 12484
rect 27068 12436 27120 12442
rect 27068 12378 27120 12384
rect 26884 12300 26936 12306
rect 26884 12242 26936 12248
rect 26896 11218 26924 12242
rect 27262 11452 27570 11461
rect 27262 11450 27268 11452
rect 27324 11450 27348 11452
rect 27404 11450 27428 11452
rect 27484 11450 27508 11452
rect 27564 11450 27570 11452
rect 27324 11398 27326 11450
rect 27506 11398 27508 11450
rect 27262 11396 27268 11398
rect 27324 11396 27348 11398
rect 27404 11396 27428 11398
rect 27484 11396 27508 11398
rect 27564 11396 27570 11398
rect 27262 11387 27570 11396
rect 26884 11212 26936 11218
rect 26884 11154 26936 11160
rect 27068 11008 27120 11014
rect 27068 10950 27120 10956
rect 26792 10668 26844 10674
rect 26792 10610 26844 10616
rect 25780 10532 25832 10538
rect 25780 10474 25832 10480
rect 25596 10260 25648 10266
rect 25596 10202 25648 10208
rect 25320 10192 25372 10198
rect 25320 10134 25372 10140
rect 24768 10124 24820 10130
rect 24768 10066 24820 10072
rect 25136 10124 25188 10130
rect 25136 10066 25188 10072
rect 25228 10124 25280 10130
rect 25228 10066 25280 10072
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 24676 9648 24728 9654
rect 24676 9590 24728 9596
rect 24872 9518 24900 9930
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25780 9920 25832 9926
rect 25780 9862 25832 9868
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 24584 9376 24636 9382
rect 24584 9318 24636 9324
rect 24398 9208 24454 9217
rect 24398 9143 24454 9152
rect 24596 9058 24624 9318
rect 24124 9036 24176 9042
rect 24124 8978 24176 8984
rect 24320 9030 24624 9058
rect 24320 8974 24348 9030
rect 24308 8968 24360 8974
rect 24122 8936 24178 8945
rect 24308 8910 24360 8916
rect 24400 8968 24452 8974
rect 24400 8910 24452 8916
rect 24122 8871 24124 8880
rect 24176 8871 24178 8880
rect 24124 8842 24176 8848
rect 23904 8732 24212 8741
rect 23904 8730 23910 8732
rect 23966 8730 23990 8732
rect 24046 8730 24070 8732
rect 24126 8730 24150 8732
rect 24206 8730 24212 8732
rect 23966 8678 23968 8730
rect 24148 8678 24150 8730
rect 23904 8676 23910 8678
rect 23966 8676 23990 8678
rect 24046 8676 24070 8678
rect 24126 8676 24150 8678
rect 24206 8676 24212 8678
rect 23904 8667 24212 8676
rect 23848 8560 23900 8566
rect 23848 8502 23900 8508
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 23480 7812 23532 7818
rect 23480 7754 23532 7760
rect 23112 7744 23164 7750
rect 23112 7686 23164 7692
rect 23124 7342 23152 7686
rect 23492 7546 23520 7754
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23584 7478 23612 7890
rect 23768 7886 23796 8434
rect 23860 7954 23888 8502
rect 24412 8129 24440 8910
rect 24492 8628 24544 8634
rect 24492 8570 24544 8576
rect 24030 8120 24086 8129
rect 24030 8055 24032 8064
rect 24084 8055 24086 8064
rect 24398 8120 24454 8129
rect 24504 8090 24532 8570
rect 24398 8055 24454 8064
rect 24492 8084 24544 8090
rect 24032 8026 24084 8032
rect 24492 8026 24544 8032
rect 24596 7993 24624 9030
rect 24768 8900 24820 8906
rect 24768 8842 24820 8848
rect 24676 8560 24728 8566
rect 24674 8528 24676 8537
rect 24728 8528 24730 8537
rect 24674 8463 24730 8472
rect 24780 8362 24808 8842
rect 24872 8838 24900 9454
rect 25042 9208 25098 9217
rect 25042 9143 25098 9152
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 24860 8832 24912 8838
rect 24860 8774 24912 8780
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24674 8256 24730 8265
rect 24674 8191 24730 8200
rect 24214 7984 24270 7993
rect 23848 7948 23900 7954
rect 24214 7919 24216 7928
rect 23848 7890 23900 7896
rect 24268 7919 24270 7928
rect 24582 7984 24638 7993
rect 24688 7954 24716 8191
rect 24780 8022 24808 8298
rect 24768 8016 24820 8022
rect 24768 7958 24820 7964
rect 24582 7919 24638 7928
rect 24676 7948 24728 7954
rect 24216 7890 24268 7896
rect 24676 7890 24728 7896
rect 23756 7880 23808 7886
rect 24872 7868 24900 8298
rect 24964 8090 24992 8978
rect 24952 8084 25004 8090
rect 24952 8026 25004 8032
rect 24780 7840 24900 7868
rect 24780 7834 24808 7840
rect 23756 7822 23808 7828
rect 24688 7806 24808 7834
rect 24308 7744 24360 7750
rect 24308 7686 24360 7692
rect 23904 7644 24212 7653
rect 23904 7642 23910 7644
rect 23966 7642 23990 7644
rect 24046 7642 24070 7644
rect 24126 7642 24150 7644
rect 24206 7642 24212 7644
rect 23966 7590 23968 7642
rect 24148 7590 24150 7642
rect 23904 7588 23910 7590
rect 23966 7588 23990 7590
rect 24046 7588 24070 7590
rect 24126 7588 24150 7590
rect 24206 7588 24212 7590
rect 23904 7579 24212 7588
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 23572 7472 23624 7478
rect 23572 7414 23624 7420
rect 23112 7336 23164 7342
rect 23112 7278 23164 7284
rect 23480 7336 23532 7342
rect 23480 7278 23532 7284
rect 23492 6458 23520 7278
rect 23664 7268 23716 7274
rect 23664 7210 23716 7216
rect 23572 6860 23624 6866
rect 23572 6802 23624 6808
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23400 5234 23428 6258
rect 23480 6248 23532 6254
rect 23480 6190 23532 6196
rect 23492 5234 23520 6190
rect 23584 5778 23612 6802
rect 23676 6254 23704 7210
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 23768 6458 23796 7142
rect 24136 6866 24164 7482
rect 24216 7336 24268 7342
rect 24320 7324 24348 7686
rect 24584 7472 24636 7478
rect 24584 7414 24636 7420
rect 24268 7296 24348 7324
rect 24216 7278 24268 7284
rect 24320 6934 24348 7296
rect 24400 7268 24452 7274
rect 24400 7210 24452 7216
rect 24492 7268 24544 7274
rect 24492 7210 24544 7216
rect 24412 7002 24440 7210
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 24308 6928 24360 6934
rect 24308 6870 24360 6876
rect 24124 6860 24176 6866
rect 24124 6802 24176 6808
rect 24504 6746 24532 7210
rect 24596 6866 24624 7414
rect 24584 6860 24636 6866
rect 24584 6802 24636 6808
rect 24412 6730 24532 6746
rect 24400 6724 24532 6730
rect 24452 6718 24532 6724
rect 24400 6666 24452 6672
rect 24308 6656 24360 6662
rect 24308 6598 24360 6604
rect 23904 6556 24212 6565
rect 23904 6554 23910 6556
rect 23966 6554 23990 6556
rect 24046 6554 24070 6556
rect 24126 6554 24150 6556
rect 24206 6554 24212 6556
rect 23966 6502 23968 6554
rect 24148 6502 24150 6554
rect 23904 6500 23910 6502
rect 23966 6500 23990 6502
rect 24046 6500 24070 6502
rect 24126 6500 24150 6502
rect 24206 6500 24212 6502
rect 23904 6491 24212 6500
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 24320 6254 24348 6598
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 24308 6248 24360 6254
rect 24308 6190 24360 6196
rect 24216 6180 24268 6186
rect 24216 6122 24268 6128
rect 24228 5778 24256 6122
rect 23572 5772 23624 5778
rect 23572 5714 23624 5720
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 23584 5370 23612 5714
rect 24216 5636 24268 5642
rect 24412 5624 24440 6666
rect 24492 6316 24544 6322
rect 24596 6304 24624 6802
rect 24544 6276 24624 6304
rect 24492 6258 24544 6264
rect 24584 6180 24636 6186
rect 24584 6122 24636 6128
rect 24596 5846 24624 6122
rect 24584 5840 24636 5846
rect 24584 5782 24636 5788
rect 24688 5794 24716 7806
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 24780 7562 24808 7686
rect 24780 7534 24900 7562
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 24780 6866 24808 7346
rect 24872 7342 24900 7534
rect 24860 7336 24912 7342
rect 24860 7278 24912 7284
rect 25056 7274 25084 9143
rect 25148 7954 25176 9862
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25240 7954 25268 9658
rect 25792 9518 25820 9862
rect 26804 9722 26832 10610
rect 27080 10130 27108 10950
rect 27262 10364 27570 10373
rect 27262 10362 27268 10364
rect 27324 10362 27348 10364
rect 27404 10362 27428 10364
rect 27484 10362 27508 10364
rect 27564 10362 27570 10364
rect 27324 10310 27326 10362
rect 27506 10310 27508 10362
rect 27262 10308 27268 10310
rect 27324 10308 27348 10310
rect 27404 10308 27428 10310
rect 27484 10308 27508 10310
rect 27564 10308 27570 10310
rect 27262 10299 27570 10308
rect 27068 10124 27120 10130
rect 27068 10066 27120 10072
rect 26884 10056 26936 10062
rect 26884 9998 26936 10004
rect 26792 9716 26844 9722
rect 26792 9658 26844 9664
rect 25412 9512 25464 9518
rect 25412 9454 25464 9460
rect 25780 9512 25832 9518
rect 25780 9454 25832 9460
rect 25320 9104 25372 9110
rect 25320 9046 25372 9052
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 25228 7948 25280 7954
rect 25228 7890 25280 7896
rect 25044 7268 25096 7274
rect 25044 7210 25096 7216
rect 24768 6860 24820 6866
rect 24768 6802 24820 6808
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 24780 5914 24808 6122
rect 25148 5914 25176 7890
rect 25240 6458 25268 7890
rect 25332 7478 25360 9046
rect 25424 9042 25452 9454
rect 26896 9178 26924 9998
rect 27262 9276 27570 9285
rect 27262 9274 27268 9276
rect 27324 9274 27348 9276
rect 27404 9274 27428 9276
rect 27484 9274 27508 9276
rect 27564 9274 27570 9276
rect 27324 9222 27326 9274
rect 27506 9222 27508 9274
rect 27262 9220 27268 9222
rect 27324 9220 27348 9222
rect 27404 9220 27428 9222
rect 27484 9220 27508 9222
rect 27564 9220 27570 9222
rect 27262 9211 27570 9220
rect 26884 9172 26936 9178
rect 26884 9114 26936 9120
rect 25872 9104 25924 9110
rect 25872 9046 25924 9052
rect 25412 9036 25464 9042
rect 25412 8978 25464 8984
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25424 8362 25452 8434
rect 25412 8356 25464 8362
rect 25412 8298 25464 8304
rect 25596 8356 25648 8362
rect 25596 8298 25648 8304
rect 25608 7993 25636 8298
rect 25780 8288 25832 8294
rect 25780 8230 25832 8236
rect 25594 7984 25650 7993
rect 25594 7919 25650 7928
rect 25320 7472 25372 7478
rect 25320 7414 25372 7420
rect 25792 7342 25820 8230
rect 25780 7336 25832 7342
rect 25780 7278 25832 7284
rect 25884 7274 25912 9046
rect 26884 8356 26936 8362
rect 26884 8298 26936 8304
rect 26896 7546 26924 8298
rect 27262 8188 27570 8197
rect 27262 8186 27268 8188
rect 27324 8186 27348 8188
rect 27404 8186 27428 8188
rect 27484 8186 27508 8188
rect 27564 8186 27570 8188
rect 27324 8134 27326 8186
rect 27506 8134 27508 8186
rect 27262 8132 27268 8134
rect 27324 8132 27348 8134
rect 27404 8132 27428 8134
rect 27484 8132 27508 8134
rect 27564 8132 27570 8134
rect 27262 8123 27570 8132
rect 26884 7540 26936 7546
rect 26884 7482 26936 7488
rect 25872 7268 25924 7274
rect 25872 7210 25924 7216
rect 25884 7002 25912 7210
rect 27262 7100 27570 7109
rect 27262 7098 27268 7100
rect 27324 7098 27348 7100
rect 27404 7098 27428 7100
rect 27484 7098 27508 7100
rect 27564 7098 27570 7100
rect 27324 7046 27326 7098
rect 27506 7046 27508 7098
rect 27262 7044 27268 7046
rect 27324 7044 27348 7046
rect 27404 7044 27428 7046
rect 27484 7044 27508 7046
rect 27564 7044 27570 7046
rect 27262 7035 27570 7044
rect 25872 6996 25924 7002
rect 25872 6938 25924 6944
rect 25872 6792 25924 6798
rect 25872 6734 25924 6740
rect 25884 6458 25912 6734
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 25872 6452 25924 6458
rect 25872 6394 25924 6400
rect 27262 6012 27570 6021
rect 27262 6010 27268 6012
rect 27324 6010 27348 6012
rect 27404 6010 27428 6012
rect 27484 6010 27508 6012
rect 27564 6010 27570 6012
rect 27324 5958 27326 6010
rect 27506 5958 27508 6010
rect 27262 5956 27268 5958
rect 27324 5956 27348 5958
rect 27404 5956 27428 5958
rect 27484 5956 27508 5958
rect 27564 5956 27570 5958
rect 27262 5947 27570 5956
rect 24768 5908 24820 5914
rect 24768 5850 24820 5856
rect 25136 5908 25188 5914
rect 25136 5850 25188 5856
rect 24268 5596 24440 5624
rect 24216 5578 24268 5584
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 23572 5364 23624 5370
rect 23572 5306 23624 5312
rect 23768 5302 23796 5510
rect 23904 5468 24212 5477
rect 23904 5466 23910 5468
rect 23966 5466 23990 5468
rect 24046 5466 24070 5468
rect 24126 5466 24150 5468
rect 24206 5466 24212 5468
rect 23966 5414 23968 5466
rect 24148 5414 24150 5466
rect 23904 5412 23910 5414
rect 23966 5412 23990 5414
rect 24046 5412 24070 5414
rect 24126 5412 24150 5414
rect 24206 5412 24212 5414
rect 23904 5403 24212 5412
rect 24412 5352 24440 5596
rect 24492 5364 24544 5370
rect 24412 5324 24492 5352
rect 23756 5296 23808 5302
rect 23756 5238 23808 5244
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23480 5228 23532 5234
rect 23480 5170 23532 5176
rect 23756 5160 23808 5166
rect 23756 5102 23808 5108
rect 23768 4826 23796 5102
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 24412 4690 24440 5324
rect 24492 5306 24544 5312
rect 24596 4842 24624 5782
rect 24688 5766 24808 5794
rect 25148 5778 25176 5850
rect 24596 4826 24716 4842
rect 24596 4820 24728 4826
rect 24596 4814 24676 4820
rect 24676 4762 24728 4768
rect 24584 4752 24636 4758
rect 24780 4706 24808 5766
rect 25136 5772 25188 5778
rect 25136 5714 25188 5720
rect 26056 5772 26108 5778
rect 26056 5714 26108 5720
rect 25136 5568 25188 5574
rect 25136 5510 25188 5516
rect 24636 4700 24808 4706
rect 24584 4694 24808 4700
rect 24400 4684 24452 4690
rect 24400 4626 24452 4632
rect 24596 4678 24808 4694
rect 23904 4380 24212 4389
rect 23904 4378 23910 4380
rect 23966 4378 23990 4380
rect 24046 4378 24070 4380
rect 24126 4378 24150 4380
rect 24206 4378 24212 4380
rect 23966 4326 23968 4378
rect 24148 4326 24150 4378
rect 23904 4324 23910 4326
rect 23966 4324 23990 4326
rect 24046 4324 24070 4326
rect 24126 4324 24150 4326
rect 24206 4324 24212 4326
rect 23904 4315 24212 4324
rect 24596 4078 24624 4678
rect 25148 4486 25176 5510
rect 26068 5370 26096 5714
rect 26056 5364 26108 5370
rect 26056 5306 26108 5312
rect 25412 5092 25464 5098
rect 25412 5034 25464 5040
rect 25424 4826 25452 5034
rect 27262 4924 27570 4933
rect 27262 4922 27268 4924
rect 27324 4922 27348 4924
rect 27404 4922 27428 4924
rect 27484 4922 27508 4924
rect 27564 4922 27570 4924
rect 27324 4870 27326 4922
rect 27506 4870 27508 4922
rect 27262 4868 27268 4870
rect 27324 4868 27348 4870
rect 27404 4868 27428 4870
rect 27484 4868 27508 4870
rect 27564 4868 27570 4870
rect 27262 4859 27570 4868
rect 25412 4820 25464 4826
rect 25412 4762 25464 4768
rect 25136 4480 25188 4486
rect 25136 4422 25188 4428
rect 24584 4072 24636 4078
rect 24584 4014 24636 4020
rect 23020 4004 23072 4010
rect 23020 3946 23072 3952
rect 27262 3836 27570 3845
rect 27262 3834 27268 3836
rect 27324 3834 27348 3836
rect 27404 3834 27428 3836
rect 27484 3834 27508 3836
rect 27564 3834 27570 3836
rect 27324 3782 27326 3834
rect 27506 3782 27508 3834
rect 27262 3780 27268 3782
rect 27324 3780 27348 3782
rect 27404 3780 27428 3782
rect 27484 3780 27508 3782
rect 27564 3780 27570 3782
rect 27262 3771 27570 3780
rect 23904 3292 24212 3301
rect 23904 3290 23910 3292
rect 23966 3290 23990 3292
rect 24046 3290 24070 3292
rect 24126 3290 24150 3292
rect 24206 3290 24212 3292
rect 23966 3238 23968 3290
rect 24148 3238 24150 3290
rect 23904 3236 23910 3238
rect 23966 3236 23990 3238
rect 24046 3236 24070 3238
rect 24126 3236 24150 3238
rect 24206 3236 24212 3238
rect 23904 3227 24212 3236
rect 20546 2748 20854 2757
rect 20546 2746 20552 2748
rect 20608 2746 20632 2748
rect 20688 2746 20712 2748
rect 20768 2746 20792 2748
rect 20848 2746 20854 2748
rect 20608 2694 20610 2746
rect 20790 2694 20792 2746
rect 20546 2692 20552 2694
rect 20608 2692 20632 2694
rect 20688 2692 20712 2694
rect 20768 2692 20792 2694
rect 20848 2692 20854 2694
rect 20546 2683 20854 2692
rect 21468 2746 21588 2774
rect 27262 2748 27570 2757
rect 27262 2746 27268 2748
rect 27324 2746 27348 2748
rect 27404 2746 27428 2748
rect 27484 2746 27508 2748
rect 27564 2746 27570 2748
rect 20626 2544 20682 2553
rect 20626 2479 20682 2488
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 20548 1970 20576 2382
rect 20536 1964 20588 1970
rect 20536 1906 20588 1912
rect 20640 1902 20668 2479
rect 21468 2378 21496 2746
rect 27324 2694 27326 2746
rect 27506 2694 27508 2746
rect 27262 2692 27268 2694
rect 27324 2692 27348 2694
rect 27404 2692 27428 2694
rect 27484 2692 27508 2694
rect 27564 2692 27570 2694
rect 27262 2683 27570 2692
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 20444 1896 20496 1902
rect 20444 1838 20496 1844
rect 20628 1896 20680 1902
rect 20628 1838 20680 1844
rect 20546 1660 20854 1669
rect 20546 1658 20552 1660
rect 20608 1658 20632 1660
rect 20688 1658 20712 1660
rect 20768 1658 20792 1660
rect 20848 1658 20854 1660
rect 20608 1606 20610 1658
rect 20790 1606 20792 1658
rect 20546 1604 20552 1606
rect 20608 1604 20632 1606
rect 20688 1604 20712 1606
rect 20768 1604 20792 1606
rect 20848 1604 20854 1606
rect 20546 1595 20854 1604
rect 21468 1494 21496 2314
rect 21456 1488 21508 1494
rect 21456 1430 21508 1436
rect 19800 1420 19852 1426
rect 19800 1362 19852 1368
rect 19892 1420 19944 1426
rect 19892 1362 19944 1368
rect 20076 1216 20128 1222
rect 20076 1158 20128 1164
rect 19708 672 19760 678
rect 19708 614 19760 620
rect 20088 400 20116 1158
rect 20546 572 20854 581
rect 20546 570 20552 572
rect 20608 570 20632 572
rect 20688 570 20712 572
rect 20768 570 20792 572
rect 20848 570 20854 572
rect 20608 518 20610 570
rect 20790 518 20792 570
rect 20546 516 20552 518
rect 20608 516 20632 518
rect 20688 516 20712 518
rect 20768 516 20792 518
rect 20848 516 20854 518
rect 20546 507 20854 516
rect 21836 400 21864 2382
rect 23904 2204 24212 2213
rect 23904 2202 23910 2204
rect 23966 2202 23990 2204
rect 24046 2202 24070 2204
rect 24126 2202 24150 2204
rect 24206 2202 24212 2204
rect 23966 2150 23968 2202
rect 24148 2150 24150 2202
rect 23904 2148 23910 2150
rect 23966 2148 23990 2150
rect 24046 2148 24070 2150
rect 24126 2148 24150 2150
rect 24206 2148 24212 2150
rect 23904 2139 24212 2148
rect 27068 1828 27120 1834
rect 27068 1770 27120 1776
rect 25320 1760 25372 1766
rect 25320 1702 25372 1708
rect 23572 1420 23624 1426
rect 23572 1362 23624 1368
rect 23584 400 23612 1362
rect 23904 1116 24212 1125
rect 23904 1114 23910 1116
rect 23966 1114 23990 1116
rect 24046 1114 24070 1116
rect 24126 1114 24150 1116
rect 24206 1114 24212 1116
rect 23966 1062 23968 1114
rect 24148 1062 24150 1114
rect 23904 1060 23910 1062
rect 23966 1060 23990 1062
rect 24046 1060 24070 1062
rect 24126 1060 24150 1062
rect 24206 1060 24212 1062
rect 23904 1051 24212 1060
rect 25332 400 25360 1702
rect 27080 400 27108 1770
rect 27262 1660 27570 1669
rect 27262 1658 27268 1660
rect 27324 1658 27348 1660
rect 27404 1658 27428 1660
rect 27484 1658 27508 1660
rect 27564 1658 27570 1660
rect 27324 1606 27326 1658
rect 27506 1606 27508 1658
rect 27262 1604 27268 1606
rect 27324 1604 27348 1606
rect 27404 1604 27428 1606
rect 27484 1604 27508 1606
rect 27564 1604 27570 1606
rect 27262 1595 27570 1604
rect 27262 572 27570 581
rect 27262 570 27268 572
rect 27324 570 27348 572
rect 27404 570 27428 572
rect 27484 570 27508 572
rect 27564 570 27570 572
rect 27324 518 27326 570
rect 27506 518 27508 570
rect 27262 516 27268 518
rect 27324 516 27348 518
rect 27404 516 27428 518
rect 27484 516 27508 518
rect 27564 516 27570 518
rect 27262 507 27570 516
rect 846 0 902 400
rect 2594 0 2650 400
rect 4342 0 4398 400
rect 6090 0 6146 400
rect 7838 0 7894 400
rect 9586 0 9642 400
rect 11334 0 11390 400
rect 13082 0 13138 400
rect 14830 0 14886 400
rect 16578 0 16634 400
rect 18326 0 18382 400
rect 20074 0 20130 400
rect 21822 0 21878 400
rect 23570 0 23626 400
rect 25318 0 25374 400
rect 27066 0 27122 400
<< via2 >>
rect 3762 17434 3818 17436
rect 3842 17434 3898 17436
rect 3922 17434 3978 17436
rect 4002 17434 4058 17436
rect 3762 17382 3808 17434
rect 3808 17382 3818 17434
rect 3842 17382 3872 17434
rect 3872 17382 3884 17434
rect 3884 17382 3898 17434
rect 3922 17382 3936 17434
rect 3936 17382 3948 17434
rect 3948 17382 3978 17434
rect 4002 17382 4012 17434
rect 4012 17382 4058 17434
rect 3762 17380 3818 17382
rect 3842 17380 3898 17382
rect 3922 17380 3978 17382
rect 4002 17380 4058 17382
rect 3762 16346 3818 16348
rect 3842 16346 3898 16348
rect 3922 16346 3978 16348
rect 4002 16346 4058 16348
rect 3762 16294 3808 16346
rect 3808 16294 3818 16346
rect 3842 16294 3872 16346
rect 3872 16294 3884 16346
rect 3884 16294 3898 16346
rect 3922 16294 3936 16346
rect 3936 16294 3948 16346
rect 3948 16294 3978 16346
rect 4002 16294 4012 16346
rect 4012 16294 4058 16346
rect 3762 16292 3818 16294
rect 3842 16292 3898 16294
rect 3922 16292 3978 16294
rect 4002 16292 4058 16294
rect 3762 15258 3818 15260
rect 3842 15258 3898 15260
rect 3922 15258 3978 15260
rect 4002 15258 4058 15260
rect 3762 15206 3808 15258
rect 3808 15206 3818 15258
rect 3842 15206 3872 15258
rect 3872 15206 3884 15258
rect 3884 15206 3898 15258
rect 3922 15206 3936 15258
rect 3936 15206 3948 15258
rect 3948 15206 3978 15258
rect 4002 15206 4012 15258
rect 4012 15206 4058 15258
rect 3762 15204 3818 15206
rect 3842 15204 3898 15206
rect 3922 15204 3978 15206
rect 4002 15204 4058 15206
rect 3762 14170 3818 14172
rect 3842 14170 3898 14172
rect 3922 14170 3978 14172
rect 4002 14170 4058 14172
rect 3762 14118 3808 14170
rect 3808 14118 3818 14170
rect 3842 14118 3872 14170
rect 3872 14118 3884 14170
rect 3884 14118 3898 14170
rect 3922 14118 3936 14170
rect 3936 14118 3948 14170
rect 3948 14118 3978 14170
rect 4002 14118 4012 14170
rect 4012 14118 4058 14170
rect 3762 14116 3818 14118
rect 3842 14116 3898 14118
rect 3922 14116 3978 14118
rect 4002 14116 4058 14118
rect 3606 13504 3662 13560
rect 3790 13388 3846 13424
rect 3790 13368 3792 13388
rect 3792 13368 3844 13388
rect 3844 13368 3846 13388
rect 4342 13504 4398 13560
rect 3762 13082 3818 13084
rect 3842 13082 3898 13084
rect 3922 13082 3978 13084
rect 4002 13082 4058 13084
rect 3762 13030 3808 13082
rect 3808 13030 3818 13082
rect 3842 13030 3872 13082
rect 3872 13030 3884 13082
rect 3884 13030 3898 13082
rect 3922 13030 3936 13082
rect 3936 13030 3948 13082
rect 3948 13030 3978 13082
rect 4002 13030 4012 13082
rect 4012 13030 4058 13082
rect 3762 13028 3818 13030
rect 3842 13028 3898 13030
rect 3922 13028 3978 13030
rect 4002 13028 4058 13030
rect 4526 13368 4582 13424
rect 3762 11994 3818 11996
rect 3842 11994 3898 11996
rect 3922 11994 3978 11996
rect 4002 11994 4058 11996
rect 3762 11942 3808 11994
rect 3808 11942 3818 11994
rect 3842 11942 3872 11994
rect 3872 11942 3884 11994
rect 3884 11942 3898 11994
rect 3922 11942 3936 11994
rect 3936 11942 3948 11994
rect 3948 11942 3978 11994
rect 4002 11942 4012 11994
rect 4012 11942 4058 11994
rect 3762 11940 3818 11942
rect 3842 11940 3898 11942
rect 3922 11940 3978 11942
rect 4002 11940 4058 11942
rect 4802 13404 4804 13424
rect 4804 13404 4856 13424
rect 4856 13404 4858 13424
rect 4802 13368 4858 13404
rect 3762 10906 3818 10908
rect 3842 10906 3898 10908
rect 3922 10906 3978 10908
rect 4002 10906 4058 10908
rect 3762 10854 3808 10906
rect 3808 10854 3818 10906
rect 3842 10854 3872 10906
rect 3872 10854 3884 10906
rect 3884 10854 3898 10906
rect 3922 10854 3936 10906
rect 3936 10854 3948 10906
rect 3948 10854 3978 10906
rect 4002 10854 4012 10906
rect 4012 10854 4058 10906
rect 3762 10852 3818 10854
rect 3842 10852 3898 10854
rect 3922 10852 3978 10854
rect 4002 10852 4058 10854
rect 3762 9818 3818 9820
rect 3842 9818 3898 9820
rect 3922 9818 3978 9820
rect 4002 9818 4058 9820
rect 3762 9766 3808 9818
rect 3808 9766 3818 9818
rect 3842 9766 3872 9818
rect 3872 9766 3884 9818
rect 3884 9766 3898 9818
rect 3922 9766 3936 9818
rect 3936 9766 3948 9818
rect 3948 9766 3978 9818
rect 4002 9766 4012 9818
rect 4012 9766 4058 9818
rect 3762 9764 3818 9766
rect 3842 9764 3898 9766
rect 3922 9764 3978 9766
rect 4002 9764 4058 9766
rect 3762 8730 3818 8732
rect 3842 8730 3898 8732
rect 3922 8730 3978 8732
rect 4002 8730 4058 8732
rect 3762 8678 3808 8730
rect 3808 8678 3818 8730
rect 3842 8678 3872 8730
rect 3872 8678 3884 8730
rect 3884 8678 3898 8730
rect 3922 8678 3936 8730
rect 3936 8678 3948 8730
rect 3948 8678 3978 8730
rect 4002 8678 4012 8730
rect 4012 8678 4058 8730
rect 3762 8676 3818 8678
rect 3842 8676 3898 8678
rect 3922 8676 3978 8678
rect 4002 8676 4058 8678
rect 3762 7642 3818 7644
rect 3842 7642 3898 7644
rect 3922 7642 3978 7644
rect 4002 7642 4058 7644
rect 3762 7590 3808 7642
rect 3808 7590 3818 7642
rect 3842 7590 3872 7642
rect 3872 7590 3884 7642
rect 3884 7590 3898 7642
rect 3922 7590 3936 7642
rect 3936 7590 3948 7642
rect 3948 7590 3978 7642
rect 4002 7590 4012 7642
rect 4012 7590 4058 7642
rect 3762 7588 3818 7590
rect 3842 7588 3898 7590
rect 3922 7588 3978 7590
rect 4002 7588 4058 7590
rect 3762 6554 3818 6556
rect 3842 6554 3898 6556
rect 3922 6554 3978 6556
rect 4002 6554 4058 6556
rect 3762 6502 3808 6554
rect 3808 6502 3818 6554
rect 3842 6502 3872 6554
rect 3872 6502 3884 6554
rect 3884 6502 3898 6554
rect 3922 6502 3936 6554
rect 3936 6502 3948 6554
rect 3948 6502 3978 6554
rect 4002 6502 4012 6554
rect 4012 6502 4058 6554
rect 3762 6500 3818 6502
rect 3842 6500 3898 6502
rect 3922 6500 3978 6502
rect 4002 6500 4058 6502
rect 3762 5466 3818 5468
rect 3842 5466 3898 5468
rect 3922 5466 3978 5468
rect 4002 5466 4058 5468
rect 3762 5414 3808 5466
rect 3808 5414 3818 5466
rect 3842 5414 3872 5466
rect 3872 5414 3884 5466
rect 3884 5414 3898 5466
rect 3922 5414 3936 5466
rect 3936 5414 3948 5466
rect 3948 5414 3978 5466
rect 4002 5414 4012 5466
rect 4012 5414 4058 5466
rect 3762 5412 3818 5414
rect 3842 5412 3898 5414
rect 3922 5412 3978 5414
rect 4002 5412 4058 5414
rect 4434 9016 4490 9072
rect 3762 4378 3818 4380
rect 3842 4378 3898 4380
rect 3922 4378 3978 4380
rect 4002 4378 4058 4380
rect 3762 4326 3808 4378
rect 3808 4326 3818 4378
rect 3842 4326 3872 4378
rect 3872 4326 3884 4378
rect 3884 4326 3898 4378
rect 3922 4326 3936 4378
rect 3936 4326 3948 4378
rect 3948 4326 3978 4378
rect 4002 4326 4012 4378
rect 4012 4326 4058 4378
rect 3762 4324 3818 4326
rect 3842 4324 3898 4326
rect 3922 4324 3978 4326
rect 4002 4324 4058 4326
rect 5814 13368 5870 13424
rect 7120 16890 7176 16892
rect 7200 16890 7256 16892
rect 7280 16890 7336 16892
rect 7360 16890 7416 16892
rect 7120 16838 7166 16890
rect 7166 16838 7176 16890
rect 7200 16838 7230 16890
rect 7230 16838 7242 16890
rect 7242 16838 7256 16890
rect 7280 16838 7294 16890
rect 7294 16838 7306 16890
rect 7306 16838 7336 16890
rect 7360 16838 7370 16890
rect 7370 16838 7416 16890
rect 7120 16836 7176 16838
rect 7200 16836 7256 16838
rect 7280 16836 7336 16838
rect 7360 16836 7416 16838
rect 7120 15802 7176 15804
rect 7200 15802 7256 15804
rect 7280 15802 7336 15804
rect 7360 15802 7416 15804
rect 7120 15750 7166 15802
rect 7166 15750 7176 15802
rect 7200 15750 7230 15802
rect 7230 15750 7242 15802
rect 7242 15750 7256 15802
rect 7280 15750 7294 15802
rect 7294 15750 7306 15802
rect 7306 15750 7336 15802
rect 7360 15750 7370 15802
rect 7370 15750 7416 15802
rect 7120 15748 7176 15750
rect 7200 15748 7256 15750
rect 7280 15748 7336 15750
rect 7360 15748 7416 15750
rect 7120 14714 7176 14716
rect 7200 14714 7256 14716
rect 7280 14714 7336 14716
rect 7360 14714 7416 14716
rect 7120 14662 7166 14714
rect 7166 14662 7176 14714
rect 7200 14662 7230 14714
rect 7230 14662 7242 14714
rect 7242 14662 7256 14714
rect 7280 14662 7294 14714
rect 7294 14662 7306 14714
rect 7306 14662 7336 14714
rect 7360 14662 7370 14714
rect 7370 14662 7416 14714
rect 7120 14660 7176 14662
rect 7200 14660 7256 14662
rect 7280 14660 7336 14662
rect 7360 14660 7416 14662
rect 7120 13626 7176 13628
rect 7200 13626 7256 13628
rect 7280 13626 7336 13628
rect 7360 13626 7416 13628
rect 7120 13574 7166 13626
rect 7166 13574 7176 13626
rect 7200 13574 7230 13626
rect 7230 13574 7242 13626
rect 7242 13574 7256 13626
rect 7280 13574 7294 13626
rect 7294 13574 7306 13626
rect 7306 13574 7336 13626
rect 7360 13574 7370 13626
rect 7370 13574 7416 13626
rect 7120 13572 7176 13574
rect 7200 13572 7256 13574
rect 7280 13572 7336 13574
rect 7360 13572 7416 13574
rect 6642 12300 6698 12336
rect 6642 12280 6644 12300
rect 6644 12280 6696 12300
rect 6696 12280 6698 12300
rect 7562 12824 7618 12880
rect 7120 12538 7176 12540
rect 7200 12538 7256 12540
rect 7280 12538 7336 12540
rect 7360 12538 7416 12540
rect 7120 12486 7166 12538
rect 7166 12486 7176 12538
rect 7200 12486 7230 12538
rect 7230 12486 7242 12538
rect 7242 12486 7256 12538
rect 7280 12486 7294 12538
rect 7294 12486 7306 12538
rect 7306 12486 7336 12538
rect 7360 12486 7370 12538
rect 7370 12486 7416 12538
rect 7120 12484 7176 12486
rect 7200 12484 7256 12486
rect 7280 12484 7336 12486
rect 7360 12484 7416 12486
rect 7120 11450 7176 11452
rect 7200 11450 7256 11452
rect 7280 11450 7336 11452
rect 7360 11450 7416 11452
rect 7120 11398 7166 11450
rect 7166 11398 7176 11450
rect 7200 11398 7230 11450
rect 7230 11398 7242 11450
rect 7242 11398 7256 11450
rect 7280 11398 7294 11450
rect 7294 11398 7306 11450
rect 7306 11398 7336 11450
rect 7360 11398 7370 11450
rect 7370 11398 7416 11450
rect 7120 11396 7176 11398
rect 7200 11396 7256 11398
rect 7280 11396 7336 11398
rect 7360 11396 7416 11398
rect 3762 3290 3818 3292
rect 3842 3290 3898 3292
rect 3922 3290 3978 3292
rect 4002 3290 4058 3292
rect 3762 3238 3808 3290
rect 3808 3238 3818 3290
rect 3842 3238 3872 3290
rect 3872 3238 3884 3290
rect 3884 3238 3898 3290
rect 3922 3238 3936 3290
rect 3936 3238 3948 3290
rect 3948 3238 3978 3290
rect 4002 3238 4012 3290
rect 4012 3238 4058 3290
rect 3762 3236 3818 3238
rect 3842 3236 3898 3238
rect 3922 3236 3978 3238
rect 4002 3236 4058 3238
rect 5078 3576 5134 3632
rect 3762 2202 3818 2204
rect 3842 2202 3898 2204
rect 3922 2202 3978 2204
rect 4002 2202 4058 2204
rect 3762 2150 3808 2202
rect 3808 2150 3818 2202
rect 3842 2150 3872 2202
rect 3872 2150 3884 2202
rect 3884 2150 3898 2202
rect 3922 2150 3936 2202
rect 3936 2150 3948 2202
rect 3948 2150 3978 2202
rect 4002 2150 4012 2202
rect 4012 2150 4058 2202
rect 3762 2148 3818 2150
rect 3842 2148 3898 2150
rect 3922 2148 3978 2150
rect 4002 2148 4058 2150
rect 3762 1114 3818 1116
rect 3842 1114 3898 1116
rect 3922 1114 3978 1116
rect 4002 1114 4058 1116
rect 3762 1062 3808 1114
rect 3808 1062 3818 1114
rect 3842 1062 3872 1114
rect 3872 1062 3884 1114
rect 3884 1062 3898 1114
rect 3922 1062 3936 1114
rect 3936 1062 3948 1114
rect 3948 1062 3978 1114
rect 4002 1062 4012 1114
rect 4012 1062 4058 1114
rect 3762 1060 3818 1062
rect 3842 1060 3898 1062
rect 3922 1060 3978 1062
rect 4002 1060 4058 1062
rect 7120 10362 7176 10364
rect 7200 10362 7256 10364
rect 7280 10362 7336 10364
rect 7360 10362 7416 10364
rect 7120 10310 7166 10362
rect 7166 10310 7176 10362
rect 7200 10310 7230 10362
rect 7230 10310 7242 10362
rect 7242 10310 7256 10362
rect 7280 10310 7294 10362
rect 7294 10310 7306 10362
rect 7306 10310 7336 10362
rect 7360 10310 7370 10362
rect 7370 10310 7416 10362
rect 7120 10308 7176 10310
rect 7200 10308 7256 10310
rect 7280 10308 7336 10310
rect 7360 10308 7416 10310
rect 8482 15564 8538 15600
rect 8482 15544 8484 15564
rect 8484 15544 8536 15564
rect 8536 15544 8538 15564
rect 9770 15952 9826 16008
rect 8850 13388 8906 13424
rect 8850 13368 8852 13388
rect 8852 13368 8904 13388
rect 8904 13368 8906 13388
rect 10478 17434 10534 17436
rect 10558 17434 10614 17436
rect 10638 17434 10694 17436
rect 10718 17434 10774 17436
rect 10478 17382 10524 17434
rect 10524 17382 10534 17434
rect 10558 17382 10588 17434
rect 10588 17382 10600 17434
rect 10600 17382 10614 17434
rect 10638 17382 10652 17434
rect 10652 17382 10664 17434
rect 10664 17382 10694 17434
rect 10718 17382 10728 17434
rect 10728 17382 10774 17434
rect 10478 17380 10534 17382
rect 10558 17380 10614 17382
rect 10638 17380 10694 17382
rect 10718 17380 10774 17382
rect 10478 16346 10534 16348
rect 10558 16346 10614 16348
rect 10638 16346 10694 16348
rect 10718 16346 10774 16348
rect 10478 16294 10524 16346
rect 10524 16294 10534 16346
rect 10558 16294 10588 16346
rect 10588 16294 10600 16346
rect 10600 16294 10614 16346
rect 10638 16294 10652 16346
rect 10652 16294 10664 16346
rect 10664 16294 10694 16346
rect 10718 16294 10728 16346
rect 10728 16294 10774 16346
rect 10478 16292 10534 16294
rect 10558 16292 10614 16294
rect 10638 16292 10694 16294
rect 10718 16292 10774 16294
rect 10478 15258 10534 15260
rect 10558 15258 10614 15260
rect 10638 15258 10694 15260
rect 10718 15258 10774 15260
rect 10478 15206 10524 15258
rect 10524 15206 10534 15258
rect 10558 15206 10588 15258
rect 10588 15206 10600 15258
rect 10600 15206 10614 15258
rect 10638 15206 10652 15258
rect 10652 15206 10664 15258
rect 10664 15206 10694 15258
rect 10718 15206 10728 15258
rect 10728 15206 10774 15258
rect 10478 15204 10534 15206
rect 10558 15204 10614 15206
rect 10638 15204 10694 15206
rect 10718 15204 10774 15206
rect 7120 9274 7176 9276
rect 7200 9274 7256 9276
rect 7280 9274 7336 9276
rect 7360 9274 7416 9276
rect 7120 9222 7166 9274
rect 7166 9222 7176 9274
rect 7200 9222 7230 9274
rect 7230 9222 7242 9274
rect 7242 9222 7256 9274
rect 7280 9222 7294 9274
rect 7294 9222 7306 9274
rect 7306 9222 7336 9274
rect 7360 9222 7370 9274
rect 7370 9222 7416 9274
rect 7120 9220 7176 9222
rect 7200 9220 7256 9222
rect 7280 9220 7336 9222
rect 7360 9220 7416 9222
rect 10478 14170 10534 14172
rect 10558 14170 10614 14172
rect 10638 14170 10694 14172
rect 10718 14170 10774 14172
rect 10478 14118 10524 14170
rect 10524 14118 10534 14170
rect 10558 14118 10588 14170
rect 10588 14118 10600 14170
rect 10600 14118 10614 14170
rect 10638 14118 10652 14170
rect 10652 14118 10664 14170
rect 10664 14118 10694 14170
rect 10718 14118 10728 14170
rect 10728 14118 10774 14170
rect 10478 14116 10534 14118
rect 10558 14116 10614 14118
rect 10638 14116 10694 14118
rect 10718 14116 10774 14118
rect 10966 13368 11022 13424
rect 10478 13082 10534 13084
rect 10558 13082 10614 13084
rect 10638 13082 10694 13084
rect 10718 13082 10774 13084
rect 10478 13030 10524 13082
rect 10524 13030 10534 13082
rect 10558 13030 10588 13082
rect 10588 13030 10600 13082
rect 10600 13030 10614 13082
rect 10638 13030 10652 13082
rect 10652 13030 10664 13082
rect 10664 13030 10694 13082
rect 10718 13030 10728 13082
rect 10728 13030 10774 13082
rect 10478 13028 10534 13030
rect 10558 13028 10614 13030
rect 10638 13028 10694 13030
rect 10718 13028 10774 13030
rect 10478 11994 10534 11996
rect 10558 11994 10614 11996
rect 10638 11994 10694 11996
rect 10718 11994 10774 11996
rect 10478 11942 10524 11994
rect 10524 11942 10534 11994
rect 10558 11942 10588 11994
rect 10588 11942 10600 11994
rect 10600 11942 10614 11994
rect 10638 11942 10652 11994
rect 10652 11942 10664 11994
rect 10664 11942 10694 11994
rect 10718 11942 10728 11994
rect 10728 11942 10774 11994
rect 10478 11940 10534 11942
rect 10558 11940 10614 11942
rect 10638 11940 10694 11942
rect 10718 11940 10774 11942
rect 10046 11600 10102 11656
rect 7120 8186 7176 8188
rect 7200 8186 7256 8188
rect 7280 8186 7336 8188
rect 7360 8186 7416 8188
rect 7120 8134 7166 8186
rect 7166 8134 7176 8186
rect 7200 8134 7230 8186
rect 7230 8134 7242 8186
rect 7242 8134 7256 8186
rect 7280 8134 7294 8186
rect 7294 8134 7306 8186
rect 7306 8134 7336 8186
rect 7360 8134 7370 8186
rect 7370 8134 7416 8186
rect 7120 8132 7176 8134
rect 7200 8132 7256 8134
rect 7280 8132 7336 8134
rect 7360 8132 7416 8134
rect 7120 7098 7176 7100
rect 7200 7098 7256 7100
rect 7280 7098 7336 7100
rect 7360 7098 7416 7100
rect 7120 7046 7166 7098
rect 7166 7046 7176 7098
rect 7200 7046 7230 7098
rect 7230 7046 7242 7098
rect 7242 7046 7256 7098
rect 7280 7046 7294 7098
rect 7294 7046 7306 7098
rect 7306 7046 7336 7098
rect 7360 7046 7370 7098
rect 7370 7046 7416 7098
rect 7120 7044 7176 7046
rect 7200 7044 7256 7046
rect 7280 7044 7336 7046
rect 7360 7044 7416 7046
rect 8298 8880 8354 8936
rect 7838 6860 7894 6896
rect 7838 6840 7840 6860
rect 7840 6840 7892 6860
rect 7892 6840 7894 6860
rect 7838 6704 7894 6760
rect 7120 6010 7176 6012
rect 7200 6010 7256 6012
rect 7280 6010 7336 6012
rect 7360 6010 7416 6012
rect 7120 5958 7166 6010
rect 7166 5958 7176 6010
rect 7200 5958 7230 6010
rect 7230 5958 7242 6010
rect 7242 5958 7256 6010
rect 7280 5958 7294 6010
rect 7294 5958 7306 6010
rect 7306 5958 7336 6010
rect 7360 5958 7370 6010
rect 7370 5958 7416 6010
rect 7120 5956 7176 5958
rect 7200 5956 7256 5958
rect 7280 5956 7336 5958
rect 7360 5956 7416 5958
rect 7930 5480 7986 5536
rect 7120 4922 7176 4924
rect 7200 4922 7256 4924
rect 7280 4922 7336 4924
rect 7360 4922 7416 4924
rect 7120 4870 7166 4922
rect 7166 4870 7176 4922
rect 7200 4870 7230 4922
rect 7230 4870 7242 4922
rect 7242 4870 7256 4922
rect 7280 4870 7294 4922
rect 7294 4870 7306 4922
rect 7306 4870 7336 4922
rect 7360 4870 7370 4922
rect 7370 4870 7416 4922
rect 7120 4868 7176 4870
rect 7200 4868 7256 4870
rect 7280 4868 7336 4870
rect 7360 4868 7416 4870
rect 9310 8880 9366 8936
rect 9494 8336 9550 8392
rect 9678 9152 9734 9208
rect 7120 3834 7176 3836
rect 7200 3834 7256 3836
rect 7280 3834 7336 3836
rect 7360 3834 7416 3836
rect 7120 3782 7166 3834
rect 7166 3782 7176 3834
rect 7200 3782 7230 3834
rect 7230 3782 7242 3834
rect 7242 3782 7256 3834
rect 7280 3782 7294 3834
rect 7294 3782 7306 3834
rect 7306 3782 7336 3834
rect 7360 3782 7370 3834
rect 7370 3782 7416 3834
rect 7120 3780 7176 3782
rect 7200 3780 7256 3782
rect 7280 3780 7336 3782
rect 7360 3780 7416 3782
rect 8758 3576 8814 3632
rect 7562 2932 7564 2952
rect 7564 2932 7616 2952
rect 7616 2932 7618 2952
rect 7562 2896 7618 2932
rect 7120 2746 7176 2748
rect 7200 2746 7256 2748
rect 7280 2746 7336 2748
rect 7360 2746 7416 2748
rect 7120 2694 7166 2746
rect 7166 2694 7176 2746
rect 7200 2694 7230 2746
rect 7230 2694 7242 2746
rect 7242 2694 7256 2746
rect 7280 2694 7294 2746
rect 7294 2694 7306 2746
rect 7306 2694 7336 2746
rect 7360 2694 7370 2746
rect 7370 2694 7416 2746
rect 7120 2692 7176 2694
rect 7200 2692 7256 2694
rect 7280 2692 7336 2694
rect 7360 2692 7416 2694
rect 8114 2896 8170 2952
rect 7120 1658 7176 1660
rect 7200 1658 7256 1660
rect 7280 1658 7336 1660
rect 7360 1658 7416 1660
rect 7120 1606 7166 1658
rect 7166 1606 7176 1658
rect 7200 1606 7230 1658
rect 7230 1606 7242 1658
rect 7242 1606 7256 1658
rect 7280 1606 7294 1658
rect 7294 1606 7306 1658
rect 7306 1606 7336 1658
rect 7360 1606 7370 1658
rect 7370 1606 7416 1658
rect 7120 1604 7176 1606
rect 7200 1604 7256 1606
rect 7280 1604 7336 1606
rect 7360 1604 7416 1606
rect 7562 1944 7618 2000
rect 7654 1808 7710 1864
rect 8390 2524 8392 2544
rect 8392 2524 8444 2544
rect 8444 2524 8446 2544
rect 8390 2488 8446 2524
rect 7120 570 7176 572
rect 7200 570 7256 572
rect 7280 570 7336 572
rect 7360 570 7416 572
rect 7120 518 7166 570
rect 7166 518 7176 570
rect 7200 518 7230 570
rect 7230 518 7242 570
rect 7242 518 7256 570
rect 7280 518 7294 570
rect 7294 518 7306 570
rect 7306 518 7336 570
rect 7360 518 7370 570
rect 7370 518 7416 570
rect 7120 516 7176 518
rect 7200 516 7256 518
rect 7280 516 7336 518
rect 7360 516 7416 518
rect 8850 3068 8852 3088
rect 8852 3068 8904 3088
rect 8904 3068 8906 3088
rect 8850 3032 8906 3068
rect 9310 3068 9312 3088
rect 9312 3068 9364 3088
rect 9364 3068 9366 3088
rect 9310 3032 9366 3068
rect 9678 3032 9734 3088
rect 9862 10104 9918 10160
rect 10966 12300 11022 12336
rect 10966 12280 10968 12300
rect 10968 12280 11020 12300
rect 11020 12280 11022 12300
rect 10478 10906 10534 10908
rect 10558 10906 10614 10908
rect 10638 10906 10694 10908
rect 10718 10906 10774 10908
rect 10478 10854 10524 10906
rect 10524 10854 10534 10906
rect 10558 10854 10588 10906
rect 10588 10854 10600 10906
rect 10600 10854 10614 10906
rect 10638 10854 10652 10906
rect 10652 10854 10664 10906
rect 10664 10854 10694 10906
rect 10718 10854 10728 10906
rect 10728 10854 10774 10906
rect 10478 10852 10534 10854
rect 10558 10852 10614 10854
rect 10638 10852 10694 10854
rect 10718 10852 10774 10854
rect 10478 9818 10534 9820
rect 10558 9818 10614 9820
rect 10638 9818 10694 9820
rect 10718 9818 10774 9820
rect 10478 9766 10524 9818
rect 10524 9766 10534 9818
rect 10558 9766 10588 9818
rect 10588 9766 10600 9818
rect 10600 9766 10614 9818
rect 10638 9766 10652 9818
rect 10652 9766 10664 9818
rect 10664 9766 10694 9818
rect 10718 9766 10728 9818
rect 10728 9766 10774 9818
rect 10478 9764 10534 9766
rect 10558 9764 10614 9766
rect 10638 9764 10694 9766
rect 10718 9764 10774 9766
rect 10478 8730 10534 8732
rect 10558 8730 10614 8732
rect 10638 8730 10694 8732
rect 10718 8730 10774 8732
rect 10478 8678 10524 8730
rect 10524 8678 10534 8730
rect 10558 8678 10588 8730
rect 10588 8678 10600 8730
rect 10600 8678 10614 8730
rect 10638 8678 10652 8730
rect 10652 8678 10664 8730
rect 10664 8678 10694 8730
rect 10718 8678 10728 8730
rect 10728 8678 10774 8730
rect 10478 8676 10534 8678
rect 10558 8676 10614 8678
rect 10638 8676 10694 8678
rect 10718 8676 10774 8678
rect 11242 8472 11298 8528
rect 10322 8336 10378 8392
rect 10478 7642 10534 7644
rect 10558 7642 10614 7644
rect 10638 7642 10694 7644
rect 10718 7642 10774 7644
rect 10478 7590 10524 7642
rect 10524 7590 10534 7642
rect 10558 7590 10588 7642
rect 10588 7590 10600 7642
rect 10600 7590 10614 7642
rect 10638 7590 10652 7642
rect 10652 7590 10664 7642
rect 10664 7590 10694 7642
rect 10718 7590 10728 7642
rect 10728 7590 10774 7642
rect 10478 7588 10534 7590
rect 10558 7588 10614 7590
rect 10638 7588 10694 7590
rect 10718 7588 10774 7590
rect 10874 6840 10930 6896
rect 10414 6740 10416 6760
rect 10416 6740 10468 6760
rect 10468 6740 10470 6760
rect 10414 6704 10470 6740
rect 10478 6554 10534 6556
rect 10558 6554 10614 6556
rect 10638 6554 10694 6556
rect 10718 6554 10774 6556
rect 10478 6502 10524 6554
rect 10524 6502 10534 6554
rect 10558 6502 10588 6554
rect 10588 6502 10600 6554
rect 10600 6502 10614 6554
rect 10638 6502 10652 6554
rect 10652 6502 10664 6554
rect 10664 6502 10694 6554
rect 10718 6502 10728 6554
rect 10728 6502 10774 6554
rect 10478 6500 10534 6502
rect 10558 6500 10614 6502
rect 10638 6500 10694 6502
rect 10718 6500 10774 6502
rect 9862 3984 9918 4040
rect 10478 5466 10534 5468
rect 10558 5466 10614 5468
rect 10638 5466 10694 5468
rect 10718 5466 10774 5468
rect 10478 5414 10524 5466
rect 10524 5414 10534 5466
rect 10558 5414 10588 5466
rect 10588 5414 10600 5466
rect 10600 5414 10614 5466
rect 10638 5414 10652 5466
rect 10652 5414 10664 5466
rect 10664 5414 10694 5466
rect 10718 5414 10728 5466
rect 10728 5414 10774 5466
rect 10478 5412 10534 5414
rect 10558 5412 10614 5414
rect 10638 5412 10694 5414
rect 10718 5412 10774 5414
rect 10478 4378 10534 4380
rect 10558 4378 10614 4380
rect 10638 4378 10694 4380
rect 10718 4378 10774 4380
rect 10478 4326 10524 4378
rect 10524 4326 10534 4378
rect 10558 4326 10588 4378
rect 10588 4326 10600 4378
rect 10600 4326 10614 4378
rect 10638 4326 10652 4378
rect 10652 4326 10664 4378
rect 10664 4326 10694 4378
rect 10718 4326 10728 4378
rect 10728 4326 10774 4378
rect 10478 4324 10534 4326
rect 10558 4324 10614 4326
rect 10638 4324 10694 4326
rect 10718 4324 10774 4326
rect 11058 4020 11060 4040
rect 11060 4020 11112 4040
rect 11112 4020 11114 4040
rect 11058 3984 11114 4020
rect 10478 3290 10534 3292
rect 10558 3290 10614 3292
rect 10638 3290 10694 3292
rect 10718 3290 10774 3292
rect 10478 3238 10524 3290
rect 10524 3238 10534 3290
rect 10558 3238 10588 3290
rect 10588 3238 10600 3290
rect 10600 3238 10614 3290
rect 10638 3238 10652 3290
rect 10652 3238 10664 3290
rect 10664 3238 10694 3290
rect 10718 3238 10728 3290
rect 10728 3238 10774 3290
rect 10478 3236 10534 3238
rect 10558 3236 10614 3238
rect 10638 3236 10694 3238
rect 10718 3236 10774 3238
rect 11610 8200 11666 8256
rect 12438 16652 12494 16688
rect 12438 16632 12440 16652
rect 12440 16632 12492 16652
rect 12492 16632 12494 16652
rect 12162 16124 12164 16144
rect 12164 16124 12216 16144
rect 12216 16124 12218 16144
rect 12162 16088 12218 16124
rect 11978 15988 11980 16008
rect 11980 15988 12032 16008
rect 12032 15988 12034 16008
rect 11978 15952 12034 15988
rect 12714 15988 12716 16008
rect 12716 15988 12768 16008
rect 12768 15988 12770 16008
rect 12714 15952 12770 15988
rect 12438 9152 12494 9208
rect 13836 16890 13892 16892
rect 13916 16890 13972 16892
rect 13996 16890 14052 16892
rect 14076 16890 14132 16892
rect 13836 16838 13882 16890
rect 13882 16838 13892 16890
rect 13916 16838 13946 16890
rect 13946 16838 13958 16890
rect 13958 16838 13972 16890
rect 13996 16838 14010 16890
rect 14010 16838 14022 16890
rect 14022 16838 14052 16890
rect 14076 16838 14086 16890
rect 14086 16838 14132 16890
rect 13836 16836 13892 16838
rect 13916 16836 13972 16838
rect 13996 16836 14052 16838
rect 14076 16836 14132 16838
rect 14646 16088 14702 16144
rect 14186 15988 14188 16008
rect 14188 15988 14240 16008
rect 14240 15988 14242 16008
rect 14186 15952 14242 15988
rect 13836 15802 13892 15804
rect 13916 15802 13972 15804
rect 13996 15802 14052 15804
rect 14076 15802 14132 15804
rect 13836 15750 13882 15802
rect 13882 15750 13892 15802
rect 13916 15750 13946 15802
rect 13946 15750 13958 15802
rect 13958 15750 13972 15802
rect 13996 15750 14010 15802
rect 14010 15750 14022 15802
rect 14022 15750 14052 15802
rect 14076 15750 14086 15802
rect 14086 15750 14132 15802
rect 13836 15748 13892 15750
rect 13916 15748 13972 15750
rect 13996 15748 14052 15750
rect 14076 15748 14132 15750
rect 12254 5908 12310 5944
rect 12254 5888 12256 5908
rect 12256 5888 12308 5908
rect 12308 5888 12310 5908
rect 11794 4020 11796 4040
rect 11796 4020 11848 4040
rect 11848 4020 11850 4040
rect 11794 3984 11850 4020
rect 13450 12144 13506 12200
rect 13174 9152 13230 9208
rect 13266 8200 13322 8256
rect 11150 2488 11206 2544
rect 10478 2202 10534 2204
rect 10558 2202 10614 2204
rect 10638 2202 10694 2204
rect 10718 2202 10774 2204
rect 10478 2150 10524 2202
rect 10524 2150 10534 2202
rect 10558 2150 10588 2202
rect 10588 2150 10600 2202
rect 10600 2150 10614 2202
rect 10638 2150 10652 2202
rect 10652 2150 10664 2202
rect 10664 2150 10694 2202
rect 10718 2150 10728 2202
rect 10728 2150 10774 2202
rect 10478 2148 10534 2150
rect 10558 2148 10614 2150
rect 10638 2148 10694 2150
rect 10718 2148 10774 2150
rect 10478 1114 10534 1116
rect 10558 1114 10614 1116
rect 10638 1114 10694 1116
rect 10718 1114 10774 1116
rect 10478 1062 10524 1114
rect 10524 1062 10534 1114
rect 10558 1062 10588 1114
rect 10588 1062 10600 1114
rect 10600 1062 10614 1114
rect 10638 1062 10652 1114
rect 10652 1062 10664 1114
rect 10664 1062 10694 1114
rect 10718 1062 10728 1114
rect 10728 1062 10774 1114
rect 10478 1060 10534 1062
rect 10558 1060 10614 1062
rect 10638 1060 10694 1062
rect 10718 1060 10774 1062
rect 13836 14714 13892 14716
rect 13916 14714 13972 14716
rect 13996 14714 14052 14716
rect 14076 14714 14132 14716
rect 13836 14662 13882 14714
rect 13882 14662 13892 14714
rect 13916 14662 13946 14714
rect 13946 14662 13958 14714
rect 13958 14662 13972 14714
rect 13996 14662 14010 14714
rect 14010 14662 14022 14714
rect 14022 14662 14052 14714
rect 14076 14662 14086 14714
rect 14086 14662 14132 14714
rect 13836 14660 13892 14662
rect 13916 14660 13972 14662
rect 13996 14660 14052 14662
rect 14076 14660 14132 14662
rect 13836 13626 13892 13628
rect 13916 13626 13972 13628
rect 13996 13626 14052 13628
rect 14076 13626 14132 13628
rect 13836 13574 13882 13626
rect 13882 13574 13892 13626
rect 13916 13574 13946 13626
rect 13946 13574 13958 13626
rect 13958 13574 13972 13626
rect 13996 13574 14010 13626
rect 14010 13574 14022 13626
rect 14022 13574 14052 13626
rect 14076 13574 14086 13626
rect 14086 13574 14132 13626
rect 13836 13572 13892 13574
rect 13916 13572 13972 13574
rect 13996 13572 14052 13574
rect 14076 13572 14132 13574
rect 13836 12538 13892 12540
rect 13916 12538 13972 12540
rect 13996 12538 14052 12540
rect 14076 12538 14132 12540
rect 13836 12486 13882 12538
rect 13882 12486 13892 12538
rect 13916 12486 13946 12538
rect 13946 12486 13958 12538
rect 13958 12486 13972 12538
rect 13996 12486 14010 12538
rect 14010 12486 14022 12538
rect 14022 12486 14052 12538
rect 14076 12486 14086 12538
rect 14086 12486 14132 12538
rect 13836 12484 13892 12486
rect 13916 12484 13972 12486
rect 13996 12484 14052 12486
rect 14076 12484 14132 12486
rect 15014 12144 15070 12200
rect 13836 11450 13892 11452
rect 13916 11450 13972 11452
rect 13996 11450 14052 11452
rect 14076 11450 14132 11452
rect 13836 11398 13882 11450
rect 13882 11398 13892 11450
rect 13916 11398 13946 11450
rect 13946 11398 13958 11450
rect 13958 11398 13972 11450
rect 13996 11398 14010 11450
rect 14010 11398 14022 11450
rect 14022 11398 14052 11450
rect 14076 11398 14086 11450
rect 14086 11398 14132 11450
rect 13836 11396 13892 11398
rect 13916 11396 13972 11398
rect 13996 11396 14052 11398
rect 14076 11396 14132 11398
rect 13836 10362 13892 10364
rect 13916 10362 13972 10364
rect 13996 10362 14052 10364
rect 14076 10362 14132 10364
rect 13836 10310 13882 10362
rect 13882 10310 13892 10362
rect 13916 10310 13946 10362
rect 13946 10310 13958 10362
rect 13958 10310 13972 10362
rect 13996 10310 14010 10362
rect 14010 10310 14022 10362
rect 14022 10310 14052 10362
rect 14076 10310 14086 10362
rect 14086 10310 14132 10362
rect 13836 10308 13892 10310
rect 13916 10308 13972 10310
rect 13996 10308 14052 10310
rect 14076 10308 14132 10310
rect 14278 9580 14334 9616
rect 14278 9560 14280 9580
rect 14280 9560 14332 9580
rect 14332 9560 14334 9580
rect 13836 9274 13892 9276
rect 13916 9274 13972 9276
rect 13996 9274 14052 9276
rect 14076 9274 14132 9276
rect 13836 9222 13882 9274
rect 13882 9222 13892 9274
rect 13916 9222 13946 9274
rect 13946 9222 13958 9274
rect 13958 9222 13972 9274
rect 13996 9222 14010 9274
rect 14010 9222 14022 9274
rect 14022 9222 14052 9274
rect 14076 9222 14086 9274
rect 14086 9222 14132 9274
rect 13836 9220 13892 9222
rect 13916 9220 13972 9222
rect 13996 9220 14052 9222
rect 14076 9220 14132 9222
rect 13836 8186 13892 8188
rect 13916 8186 13972 8188
rect 13996 8186 14052 8188
rect 14076 8186 14132 8188
rect 13836 8134 13882 8186
rect 13882 8134 13892 8186
rect 13916 8134 13946 8186
rect 13946 8134 13958 8186
rect 13958 8134 13972 8186
rect 13996 8134 14010 8186
rect 14010 8134 14022 8186
rect 14022 8134 14052 8186
rect 14076 8134 14086 8186
rect 14086 8134 14132 8186
rect 13836 8132 13892 8134
rect 13916 8132 13972 8134
rect 13996 8132 14052 8134
rect 14076 8132 14132 8134
rect 15106 8336 15162 8392
rect 13836 7098 13892 7100
rect 13916 7098 13972 7100
rect 13996 7098 14052 7100
rect 14076 7098 14132 7100
rect 13836 7046 13882 7098
rect 13882 7046 13892 7098
rect 13916 7046 13946 7098
rect 13946 7046 13958 7098
rect 13958 7046 13972 7098
rect 13996 7046 14010 7098
rect 14010 7046 14022 7098
rect 14022 7046 14052 7098
rect 14076 7046 14086 7098
rect 14086 7046 14132 7098
rect 13836 7044 13892 7046
rect 13916 7044 13972 7046
rect 13996 7044 14052 7046
rect 14076 7044 14132 7046
rect 13836 6010 13892 6012
rect 13916 6010 13972 6012
rect 13996 6010 14052 6012
rect 14076 6010 14132 6012
rect 13836 5958 13882 6010
rect 13882 5958 13892 6010
rect 13916 5958 13946 6010
rect 13946 5958 13958 6010
rect 13958 5958 13972 6010
rect 13996 5958 14010 6010
rect 14010 5958 14022 6010
rect 14022 5958 14052 6010
rect 14076 5958 14086 6010
rect 14086 5958 14132 6010
rect 13836 5956 13892 5958
rect 13916 5956 13972 5958
rect 13996 5956 14052 5958
rect 14076 5956 14132 5958
rect 13450 5208 13506 5264
rect 13836 4922 13892 4924
rect 13916 4922 13972 4924
rect 13996 4922 14052 4924
rect 14076 4922 14132 4924
rect 13836 4870 13882 4922
rect 13882 4870 13892 4922
rect 13916 4870 13946 4922
rect 13946 4870 13958 4922
rect 13958 4870 13972 4922
rect 13996 4870 14010 4922
rect 14010 4870 14022 4922
rect 14022 4870 14052 4922
rect 14076 4870 14086 4922
rect 14086 4870 14132 4922
rect 13836 4868 13892 4870
rect 13916 4868 13972 4870
rect 13996 4868 14052 4870
rect 14076 4868 14132 4870
rect 13836 3834 13892 3836
rect 13916 3834 13972 3836
rect 13996 3834 14052 3836
rect 14076 3834 14132 3836
rect 13836 3782 13882 3834
rect 13882 3782 13892 3834
rect 13916 3782 13946 3834
rect 13946 3782 13958 3834
rect 13958 3782 13972 3834
rect 13996 3782 14010 3834
rect 14010 3782 14022 3834
rect 14022 3782 14052 3834
rect 14076 3782 14086 3834
rect 14086 3782 14132 3834
rect 13836 3780 13892 3782
rect 13916 3780 13972 3782
rect 13996 3780 14052 3782
rect 14076 3780 14132 3782
rect 14278 3576 14334 3632
rect 13910 3440 13966 3496
rect 13836 2746 13892 2748
rect 13916 2746 13972 2748
rect 13996 2746 14052 2748
rect 14076 2746 14132 2748
rect 13836 2694 13882 2746
rect 13882 2694 13892 2746
rect 13916 2694 13946 2746
rect 13946 2694 13958 2746
rect 13958 2694 13972 2746
rect 13996 2694 14010 2746
rect 14010 2694 14022 2746
rect 14022 2694 14052 2746
rect 14076 2694 14086 2746
rect 14086 2694 14132 2746
rect 13836 2692 13892 2694
rect 13916 2692 13972 2694
rect 13996 2692 14052 2694
rect 14076 2692 14132 2694
rect 13836 1658 13892 1660
rect 13916 1658 13972 1660
rect 13996 1658 14052 1660
rect 14076 1658 14132 1660
rect 13836 1606 13882 1658
rect 13882 1606 13892 1658
rect 13916 1606 13946 1658
rect 13946 1606 13958 1658
rect 13958 1606 13972 1658
rect 13996 1606 14010 1658
rect 14010 1606 14022 1658
rect 14022 1606 14052 1658
rect 14076 1606 14086 1658
rect 14086 1606 14132 1658
rect 13836 1604 13892 1606
rect 13916 1604 13972 1606
rect 13996 1604 14052 1606
rect 14076 1604 14132 1606
rect 15750 12280 15806 12336
rect 17194 17434 17250 17436
rect 17274 17434 17330 17436
rect 17354 17434 17410 17436
rect 17434 17434 17490 17436
rect 17194 17382 17240 17434
rect 17240 17382 17250 17434
rect 17274 17382 17304 17434
rect 17304 17382 17316 17434
rect 17316 17382 17330 17434
rect 17354 17382 17368 17434
rect 17368 17382 17380 17434
rect 17380 17382 17410 17434
rect 17434 17382 17444 17434
rect 17444 17382 17490 17434
rect 17194 17380 17250 17382
rect 17274 17380 17330 17382
rect 17354 17380 17410 17382
rect 17434 17380 17490 17382
rect 23910 17434 23966 17436
rect 23990 17434 24046 17436
rect 24070 17434 24126 17436
rect 24150 17434 24206 17436
rect 23910 17382 23956 17434
rect 23956 17382 23966 17434
rect 23990 17382 24020 17434
rect 24020 17382 24032 17434
rect 24032 17382 24046 17434
rect 24070 17382 24084 17434
rect 24084 17382 24096 17434
rect 24096 17382 24126 17434
rect 24150 17382 24160 17434
rect 24160 17382 24206 17434
rect 23910 17380 23966 17382
rect 23990 17380 24046 17382
rect 24070 17380 24126 17382
rect 24150 17380 24206 17382
rect 16026 9444 16082 9480
rect 16026 9424 16028 9444
rect 16028 9424 16080 9444
rect 16080 9424 16082 9444
rect 17130 16632 17186 16688
rect 17194 16346 17250 16348
rect 17274 16346 17330 16348
rect 17354 16346 17410 16348
rect 17434 16346 17490 16348
rect 17194 16294 17240 16346
rect 17240 16294 17250 16346
rect 17274 16294 17304 16346
rect 17304 16294 17316 16346
rect 17316 16294 17330 16346
rect 17354 16294 17368 16346
rect 17368 16294 17380 16346
rect 17380 16294 17410 16346
rect 17434 16294 17444 16346
rect 17444 16294 17490 16346
rect 17194 16292 17250 16294
rect 17274 16292 17330 16294
rect 17354 16292 17410 16294
rect 17434 16292 17490 16294
rect 17958 15544 18014 15600
rect 17194 15258 17250 15260
rect 17274 15258 17330 15260
rect 17354 15258 17410 15260
rect 17434 15258 17490 15260
rect 17194 15206 17240 15258
rect 17240 15206 17250 15258
rect 17274 15206 17304 15258
rect 17304 15206 17316 15258
rect 17316 15206 17330 15258
rect 17354 15206 17368 15258
rect 17368 15206 17380 15258
rect 17380 15206 17410 15258
rect 17434 15206 17444 15258
rect 17444 15206 17490 15258
rect 17194 15204 17250 15206
rect 17274 15204 17330 15206
rect 17354 15204 17410 15206
rect 17434 15204 17490 15206
rect 17194 14170 17250 14172
rect 17274 14170 17330 14172
rect 17354 14170 17410 14172
rect 17434 14170 17490 14172
rect 17194 14118 17240 14170
rect 17240 14118 17250 14170
rect 17274 14118 17304 14170
rect 17304 14118 17316 14170
rect 17316 14118 17330 14170
rect 17354 14118 17368 14170
rect 17368 14118 17380 14170
rect 17380 14118 17410 14170
rect 17434 14118 17444 14170
rect 17444 14118 17490 14170
rect 17194 14116 17250 14118
rect 17274 14116 17330 14118
rect 17354 14116 17410 14118
rect 17434 14116 17490 14118
rect 17774 13524 17830 13560
rect 17774 13504 17776 13524
rect 17776 13504 17828 13524
rect 17828 13504 17830 13524
rect 17194 13082 17250 13084
rect 17274 13082 17330 13084
rect 17354 13082 17410 13084
rect 17434 13082 17490 13084
rect 17194 13030 17240 13082
rect 17240 13030 17250 13082
rect 17274 13030 17304 13082
rect 17304 13030 17316 13082
rect 17316 13030 17330 13082
rect 17354 13030 17368 13082
rect 17368 13030 17380 13082
rect 17380 13030 17410 13082
rect 17434 13030 17444 13082
rect 17444 13030 17490 13082
rect 17194 13028 17250 13030
rect 17274 13028 17330 13030
rect 17354 13028 17410 13030
rect 17434 13028 17490 13030
rect 17194 11994 17250 11996
rect 17274 11994 17330 11996
rect 17354 11994 17410 11996
rect 17434 11994 17490 11996
rect 17194 11942 17240 11994
rect 17240 11942 17250 11994
rect 17274 11942 17304 11994
rect 17304 11942 17316 11994
rect 17316 11942 17330 11994
rect 17354 11942 17368 11994
rect 17368 11942 17380 11994
rect 17380 11942 17410 11994
rect 17434 11942 17444 11994
rect 17444 11942 17490 11994
rect 17194 11940 17250 11942
rect 17274 11940 17330 11942
rect 17354 11940 17410 11942
rect 17434 11940 17490 11942
rect 17194 10906 17250 10908
rect 17274 10906 17330 10908
rect 17354 10906 17410 10908
rect 17434 10906 17490 10908
rect 17194 10854 17240 10906
rect 17240 10854 17250 10906
rect 17274 10854 17304 10906
rect 17304 10854 17316 10906
rect 17316 10854 17330 10906
rect 17354 10854 17368 10906
rect 17368 10854 17380 10906
rect 17380 10854 17410 10906
rect 17434 10854 17444 10906
rect 17444 10854 17490 10906
rect 17194 10852 17250 10854
rect 17274 10852 17330 10854
rect 17354 10852 17410 10854
rect 17434 10852 17490 10854
rect 17194 9818 17250 9820
rect 17274 9818 17330 9820
rect 17354 9818 17410 9820
rect 17434 9818 17490 9820
rect 17194 9766 17240 9818
rect 17240 9766 17250 9818
rect 17274 9766 17304 9818
rect 17304 9766 17316 9818
rect 17316 9766 17330 9818
rect 17354 9766 17368 9818
rect 17368 9766 17380 9818
rect 17380 9766 17410 9818
rect 17434 9766 17444 9818
rect 17444 9766 17490 9818
rect 17194 9764 17250 9766
rect 17274 9764 17330 9766
rect 17354 9764 17410 9766
rect 17434 9764 17490 9766
rect 17194 8730 17250 8732
rect 17274 8730 17330 8732
rect 17354 8730 17410 8732
rect 17434 8730 17490 8732
rect 17194 8678 17240 8730
rect 17240 8678 17250 8730
rect 17274 8678 17304 8730
rect 17304 8678 17316 8730
rect 17316 8678 17330 8730
rect 17354 8678 17368 8730
rect 17368 8678 17380 8730
rect 17380 8678 17410 8730
rect 17434 8678 17444 8730
rect 17444 8678 17490 8730
rect 17194 8676 17250 8678
rect 17274 8676 17330 8678
rect 17354 8676 17410 8678
rect 17434 8676 17490 8678
rect 17194 7642 17250 7644
rect 17274 7642 17330 7644
rect 17354 7642 17410 7644
rect 17434 7642 17490 7644
rect 17194 7590 17240 7642
rect 17240 7590 17250 7642
rect 17274 7590 17304 7642
rect 17304 7590 17316 7642
rect 17316 7590 17330 7642
rect 17354 7590 17368 7642
rect 17368 7590 17380 7642
rect 17380 7590 17410 7642
rect 17434 7590 17444 7642
rect 17444 7590 17490 7642
rect 17194 7588 17250 7590
rect 17274 7588 17330 7590
rect 17354 7588 17410 7590
rect 17434 7588 17490 7590
rect 18050 9016 18106 9072
rect 17194 6554 17250 6556
rect 17274 6554 17330 6556
rect 17354 6554 17410 6556
rect 17434 6554 17490 6556
rect 17194 6502 17240 6554
rect 17240 6502 17250 6554
rect 17274 6502 17304 6554
rect 17304 6502 17316 6554
rect 17316 6502 17330 6554
rect 17354 6502 17368 6554
rect 17368 6502 17380 6554
rect 17380 6502 17410 6554
rect 17434 6502 17444 6554
rect 17444 6502 17490 6554
rect 17194 6500 17250 6502
rect 17274 6500 17330 6502
rect 17354 6500 17410 6502
rect 17434 6500 17490 6502
rect 16394 4700 16396 4720
rect 16396 4700 16448 4720
rect 16448 4700 16450 4720
rect 16394 4664 16450 4700
rect 17194 5466 17250 5468
rect 17274 5466 17330 5468
rect 17354 5466 17410 5468
rect 17434 5466 17490 5468
rect 17194 5414 17240 5466
rect 17240 5414 17250 5466
rect 17274 5414 17304 5466
rect 17304 5414 17316 5466
rect 17316 5414 17330 5466
rect 17354 5414 17368 5466
rect 17368 5414 17380 5466
rect 17380 5414 17410 5466
rect 17434 5414 17444 5466
rect 17444 5414 17490 5466
rect 17194 5412 17250 5414
rect 17274 5412 17330 5414
rect 17354 5412 17410 5414
rect 17434 5412 17490 5414
rect 17130 5208 17186 5264
rect 17038 4700 17040 4720
rect 17040 4700 17092 4720
rect 17092 4700 17094 4720
rect 17038 4664 17094 4700
rect 17194 4378 17250 4380
rect 17274 4378 17330 4380
rect 17354 4378 17410 4380
rect 17434 4378 17490 4380
rect 17194 4326 17240 4378
rect 17240 4326 17250 4378
rect 17274 4326 17304 4378
rect 17304 4326 17316 4378
rect 17316 4326 17330 4378
rect 17354 4326 17368 4378
rect 17368 4326 17380 4378
rect 17380 4326 17410 4378
rect 17434 4326 17444 4378
rect 17444 4326 17490 4378
rect 17194 4324 17250 4326
rect 17274 4324 17330 4326
rect 17354 4324 17410 4326
rect 17434 4324 17490 4326
rect 16946 3440 17002 3496
rect 15934 1944 15990 2000
rect 17194 3290 17250 3292
rect 17274 3290 17330 3292
rect 17354 3290 17410 3292
rect 17434 3290 17490 3292
rect 17194 3238 17240 3290
rect 17240 3238 17250 3290
rect 17274 3238 17304 3290
rect 17304 3238 17316 3290
rect 17316 3238 17330 3290
rect 17354 3238 17368 3290
rect 17368 3238 17380 3290
rect 17380 3238 17410 3290
rect 17434 3238 17444 3290
rect 17444 3238 17490 3290
rect 17194 3236 17250 3238
rect 17274 3236 17330 3238
rect 17354 3236 17410 3238
rect 17434 3236 17490 3238
rect 17958 3032 18014 3088
rect 17194 2202 17250 2204
rect 17274 2202 17330 2204
rect 17354 2202 17410 2204
rect 17434 2202 17490 2204
rect 17194 2150 17240 2202
rect 17240 2150 17250 2202
rect 17274 2150 17304 2202
rect 17304 2150 17316 2202
rect 17316 2150 17330 2202
rect 17354 2150 17368 2202
rect 17368 2150 17380 2202
rect 17380 2150 17410 2202
rect 17434 2150 17444 2202
rect 17444 2150 17490 2202
rect 17194 2148 17250 2150
rect 17274 2148 17330 2150
rect 17354 2148 17410 2150
rect 17434 2148 17490 2150
rect 13836 570 13892 572
rect 13916 570 13972 572
rect 13996 570 14052 572
rect 14076 570 14132 572
rect 13836 518 13882 570
rect 13882 518 13892 570
rect 13916 518 13946 570
rect 13946 518 13958 570
rect 13958 518 13972 570
rect 13996 518 14010 570
rect 14010 518 14022 570
rect 14022 518 14052 570
rect 14076 518 14086 570
rect 14086 518 14132 570
rect 13836 516 13892 518
rect 13916 516 13972 518
rect 13996 516 14052 518
rect 14076 516 14132 518
rect 17958 1944 18014 2000
rect 18602 12300 18658 12336
rect 18602 12280 18604 12300
rect 18604 12280 18656 12300
rect 18656 12280 18658 12300
rect 18602 10124 18658 10160
rect 18602 10104 18604 10124
rect 18604 10104 18656 10124
rect 18656 10104 18658 10124
rect 19062 10124 19118 10160
rect 19062 10104 19064 10124
rect 19064 10104 19116 10124
rect 19116 10104 19118 10124
rect 19430 14864 19486 14920
rect 19246 13504 19302 13560
rect 20552 16890 20608 16892
rect 20632 16890 20688 16892
rect 20712 16890 20768 16892
rect 20792 16890 20848 16892
rect 20552 16838 20598 16890
rect 20598 16838 20608 16890
rect 20632 16838 20662 16890
rect 20662 16838 20674 16890
rect 20674 16838 20688 16890
rect 20712 16838 20726 16890
rect 20726 16838 20738 16890
rect 20738 16838 20768 16890
rect 20792 16838 20802 16890
rect 20802 16838 20848 16890
rect 20552 16836 20608 16838
rect 20632 16836 20688 16838
rect 20712 16836 20768 16838
rect 20792 16836 20848 16838
rect 20552 15802 20608 15804
rect 20632 15802 20688 15804
rect 20712 15802 20768 15804
rect 20792 15802 20848 15804
rect 20552 15750 20598 15802
rect 20598 15750 20608 15802
rect 20632 15750 20662 15802
rect 20662 15750 20674 15802
rect 20674 15750 20688 15802
rect 20712 15750 20726 15802
rect 20726 15750 20738 15802
rect 20738 15750 20768 15802
rect 20792 15750 20802 15802
rect 20802 15750 20848 15802
rect 20552 15748 20608 15750
rect 20632 15748 20688 15750
rect 20712 15748 20768 15750
rect 20792 15748 20848 15750
rect 20810 14900 20812 14920
rect 20812 14900 20864 14920
rect 20864 14900 20866 14920
rect 20810 14864 20866 14900
rect 20552 14714 20608 14716
rect 20632 14714 20688 14716
rect 20712 14714 20768 14716
rect 20792 14714 20848 14716
rect 20552 14662 20598 14714
rect 20598 14662 20608 14714
rect 20632 14662 20662 14714
rect 20662 14662 20674 14714
rect 20674 14662 20688 14714
rect 20712 14662 20726 14714
rect 20726 14662 20738 14714
rect 20738 14662 20768 14714
rect 20792 14662 20802 14714
rect 20802 14662 20848 14714
rect 20552 14660 20608 14662
rect 20632 14660 20688 14662
rect 20712 14660 20768 14662
rect 20792 14660 20848 14662
rect 23910 16346 23966 16348
rect 23990 16346 24046 16348
rect 24070 16346 24126 16348
rect 24150 16346 24206 16348
rect 23910 16294 23956 16346
rect 23956 16294 23966 16346
rect 23990 16294 24020 16346
rect 24020 16294 24032 16346
rect 24032 16294 24046 16346
rect 24070 16294 24084 16346
rect 24084 16294 24096 16346
rect 24096 16294 24126 16346
rect 24150 16294 24160 16346
rect 24160 16294 24206 16346
rect 23910 16292 23966 16294
rect 23990 16292 24046 16294
rect 24070 16292 24126 16294
rect 24150 16292 24206 16294
rect 20552 13626 20608 13628
rect 20632 13626 20688 13628
rect 20712 13626 20768 13628
rect 20792 13626 20848 13628
rect 20552 13574 20598 13626
rect 20598 13574 20608 13626
rect 20632 13574 20662 13626
rect 20662 13574 20674 13626
rect 20674 13574 20688 13626
rect 20712 13574 20726 13626
rect 20726 13574 20738 13626
rect 20738 13574 20768 13626
rect 20792 13574 20802 13626
rect 20802 13574 20848 13626
rect 20552 13572 20608 13574
rect 20632 13572 20688 13574
rect 20712 13572 20768 13574
rect 20792 13572 20848 13574
rect 19430 8472 19486 8528
rect 20350 13368 20406 13424
rect 20166 12824 20222 12880
rect 20626 12824 20682 12880
rect 20552 12538 20608 12540
rect 20632 12538 20688 12540
rect 20712 12538 20768 12540
rect 20792 12538 20848 12540
rect 20552 12486 20598 12538
rect 20598 12486 20608 12538
rect 20632 12486 20662 12538
rect 20662 12486 20674 12538
rect 20674 12486 20688 12538
rect 20712 12486 20726 12538
rect 20726 12486 20738 12538
rect 20738 12486 20768 12538
rect 20792 12486 20802 12538
rect 20802 12486 20848 12538
rect 20552 12484 20608 12486
rect 20632 12484 20688 12486
rect 20712 12484 20768 12486
rect 20792 12484 20848 12486
rect 19246 1420 19302 1456
rect 19246 1400 19248 1420
rect 19248 1400 19300 1420
rect 19300 1400 19302 1420
rect 17194 1114 17250 1116
rect 17274 1114 17330 1116
rect 17354 1114 17410 1116
rect 17434 1114 17490 1116
rect 17194 1062 17240 1114
rect 17240 1062 17250 1114
rect 17274 1062 17304 1114
rect 17304 1062 17316 1114
rect 17316 1062 17330 1114
rect 17354 1062 17368 1114
rect 17368 1062 17380 1114
rect 17380 1062 17410 1114
rect 17434 1062 17444 1114
rect 17444 1062 17490 1114
rect 17194 1060 17250 1062
rect 17274 1060 17330 1062
rect 17354 1060 17410 1062
rect 17434 1060 17490 1062
rect 20552 11450 20608 11452
rect 20632 11450 20688 11452
rect 20712 11450 20768 11452
rect 20792 11450 20848 11452
rect 20552 11398 20598 11450
rect 20598 11398 20608 11450
rect 20632 11398 20662 11450
rect 20662 11398 20674 11450
rect 20674 11398 20688 11450
rect 20712 11398 20726 11450
rect 20726 11398 20738 11450
rect 20738 11398 20768 11450
rect 20792 11398 20802 11450
rect 20802 11398 20848 11450
rect 20552 11396 20608 11398
rect 20632 11396 20688 11398
rect 20712 11396 20768 11398
rect 20792 11396 20848 11398
rect 20552 10362 20608 10364
rect 20632 10362 20688 10364
rect 20712 10362 20768 10364
rect 20792 10362 20848 10364
rect 20552 10310 20598 10362
rect 20598 10310 20608 10362
rect 20632 10310 20662 10362
rect 20662 10310 20674 10362
rect 20674 10310 20688 10362
rect 20712 10310 20726 10362
rect 20726 10310 20738 10362
rect 20738 10310 20768 10362
rect 20792 10310 20802 10362
rect 20802 10310 20848 10362
rect 20552 10308 20608 10310
rect 20632 10308 20688 10310
rect 20712 10308 20768 10310
rect 20792 10308 20848 10310
rect 20552 9274 20608 9276
rect 20632 9274 20688 9276
rect 20712 9274 20768 9276
rect 20792 9274 20848 9276
rect 20552 9222 20598 9274
rect 20598 9222 20608 9274
rect 20632 9222 20662 9274
rect 20662 9222 20674 9274
rect 20674 9222 20688 9274
rect 20712 9222 20726 9274
rect 20726 9222 20738 9274
rect 20738 9222 20768 9274
rect 20792 9222 20802 9274
rect 20802 9222 20848 9274
rect 20552 9220 20608 9222
rect 20632 9220 20688 9222
rect 20712 9220 20768 9222
rect 20792 9220 20848 9222
rect 20552 8186 20608 8188
rect 20632 8186 20688 8188
rect 20712 8186 20768 8188
rect 20792 8186 20848 8188
rect 20552 8134 20598 8186
rect 20598 8134 20608 8186
rect 20632 8134 20662 8186
rect 20662 8134 20674 8186
rect 20674 8134 20688 8186
rect 20712 8134 20726 8186
rect 20726 8134 20738 8186
rect 20738 8134 20768 8186
rect 20792 8134 20802 8186
rect 20802 8134 20848 8186
rect 20552 8132 20608 8134
rect 20632 8132 20688 8134
rect 20712 8132 20768 8134
rect 20792 8132 20848 8134
rect 20626 7656 20682 7712
rect 20552 7098 20608 7100
rect 20632 7098 20688 7100
rect 20712 7098 20768 7100
rect 20792 7098 20848 7100
rect 20552 7046 20598 7098
rect 20598 7046 20608 7098
rect 20632 7046 20662 7098
rect 20662 7046 20674 7098
rect 20674 7046 20688 7098
rect 20712 7046 20726 7098
rect 20726 7046 20738 7098
rect 20738 7046 20768 7098
rect 20792 7046 20802 7098
rect 20802 7046 20848 7098
rect 20552 7044 20608 7046
rect 20632 7044 20688 7046
rect 20712 7044 20768 7046
rect 20792 7044 20848 7046
rect 21914 14864 21970 14920
rect 21362 8880 21418 8936
rect 20552 6010 20608 6012
rect 20632 6010 20688 6012
rect 20712 6010 20768 6012
rect 20792 6010 20848 6012
rect 20552 5958 20598 6010
rect 20598 5958 20608 6010
rect 20632 5958 20662 6010
rect 20662 5958 20674 6010
rect 20674 5958 20688 6010
rect 20712 5958 20726 6010
rect 20726 5958 20738 6010
rect 20738 5958 20768 6010
rect 20792 5958 20802 6010
rect 20802 5958 20848 6010
rect 20552 5956 20608 5958
rect 20632 5956 20688 5958
rect 20712 5956 20768 5958
rect 20792 5956 20848 5958
rect 20552 4922 20608 4924
rect 20632 4922 20688 4924
rect 20712 4922 20768 4924
rect 20792 4922 20848 4924
rect 20552 4870 20598 4922
rect 20598 4870 20608 4922
rect 20632 4870 20662 4922
rect 20662 4870 20674 4922
rect 20674 4870 20688 4922
rect 20712 4870 20726 4922
rect 20726 4870 20738 4922
rect 20738 4870 20768 4922
rect 20792 4870 20802 4922
rect 20802 4870 20848 4922
rect 20552 4868 20608 4870
rect 20632 4868 20688 4870
rect 20712 4868 20768 4870
rect 20792 4868 20848 4870
rect 20552 3834 20608 3836
rect 20632 3834 20688 3836
rect 20712 3834 20768 3836
rect 20792 3834 20848 3836
rect 20552 3782 20598 3834
rect 20598 3782 20608 3834
rect 20632 3782 20662 3834
rect 20662 3782 20674 3834
rect 20674 3782 20688 3834
rect 20712 3782 20726 3834
rect 20726 3782 20738 3834
rect 20738 3782 20768 3834
rect 20792 3782 20802 3834
rect 20802 3782 20848 3834
rect 20552 3780 20608 3782
rect 20632 3780 20688 3782
rect 20712 3780 20768 3782
rect 20792 3780 20848 3782
rect 20350 2488 20406 2544
rect 22834 15544 22890 15600
rect 22926 14476 22982 14512
rect 22926 14456 22928 14476
rect 22928 14456 22980 14476
rect 22980 14456 22982 14476
rect 23910 15258 23966 15260
rect 23990 15258 24046 15260
rect 24070 15258 24126 15260
rect 24150 15258 24206 15260
rect 23910 15206 23956 15258
rect 23956 15206 23966 15258
rect 23990 15206 24020 15258
rect 24020 15206 24032 15258
rect 24032 15206 24046 15258
rect 24070 15206 24084 15258
rect 24084 15206 24096 15258
rect 24096 15206 24126 15258
rect 24150 15206 24160 15258
rect 24160 15206 24206 15258
rect 23910 15204 23966 15206
rect 23990 15204 24046 15206
rect 24070 15204 24126 15206
rect 24150 15204 24206 15206
rect 23910 14170 23966 14172
rect 23990 14170 24046 14172
rect 24070 14170 24126 14172
rect 24150 14170 24206 14172
rect 23910 14118 23956 14170
rect 23956 14118 23966 14170
rect 23990 14118 24020 14170
rect 24020 14118 24032 14170
rect 24032 14118 24046 14170
rect 24070 14118 24084 14170
rect 24084 14118 24096 14170
rect 24096 14118 24126 14170
rect 24150 14118 24160 14170
rect 24160 14118 24206 14170
rect 23910 14116 23966 14118
rect 23990 14116 24046 14118
rect 24070 14116 24126 14118
rect 24150 14116 24206 14118
rect 23910 13082 23966 13084
rect 23990 13082 24046 13084
rect 24070 13082 24126 13084
rect 24150 13082 24206 13084
rect 23910 13030 23956 13082
rect 23956 13030 23966 13082
rect 23990 13030 24020 13082
rect 24020 13030 24032 13082
rect 24032 13030 24046 13082
rect 24070 13030 24084 13082
rect 24084 13030 24096 13082
rect 24096 13030 24126 13082
rect 24150 13030 24160 13082
rect 24160 13030 24206 13082
rect 23910 13028 23966 13030
rect 23990 13028 24046 13030
rect 24070 13028 24126 13030
rect 24150 13028 24206 13030
rect 24306 12724 24308 12744
rect 24308 12724 24360 12744
rect 24360 12724 24362 12744
rect 24306 12688 24362 12724
rect 21638 7948 21694 7984
rect 21638 7928 21640 7948
rect 21640 7928 21692 7948
rect 21692 7928 21694 7948
rect 22282 7656 22338 7712
rect 22834 7656 22890 7712
rect 23910 11994 23966 11996
rect 23990 11994 24046 11996
rect 24070 11994 24126 11996
rect 24150 11994 24206 11996
rect 23910 11942 23956 11994
rect 23956 11942 23966 11994
rect 23990 11942 24020 11994
rect 24020 11942 24032 11994
rect 24032 11942 24046 11994
rect 24070 11942 24084 11994
rect 24084 11942 24096 11994
rect 24096 11942 24126 11994
rect 24150 11942 24160 11994
rect 24160 11942 24206 11994
rect 23910 11940 23966 11942
rect 23990 11940 24046 11942
rect 24070 11940 24126 11942
rect 24150 11940 24206 11942
rect 23910 10906 23966 10908
rect 23990 10906 24046 10908
rect 24070 10906 24126 10908
rect 24150 10906 24206 10908
rect 23910 10854 23956 10906
rect 23956 10854 23966 10906
rect 23990 10854 24020 10906
rect 24020 10854 24032 10906
rect 24032 10854 24046 10906
rect 24070 10854 24084 10906
rect 24084 10854 24096 10906
rect 24096 10854 24126 10906
rect 24150 10854 24160 10906
rect 24160 10854 24206 10906
rect 23910 10852 23966 10854
rect 23990 10852 24046 10854
rect 24070 10852 24126 10854
rect 24150 10852 24206 10854
rect 23910 9818 23966 9820
rect 23990 9818 24046 9820
rect 24070 9818 24126 9820
rect 24150 9818 24206 9820
rect 23910 9766 23956 9818
rect 23956 9766 23966 9818
rect 23990 9766 24020 9818
rect 24020 9766 24032 9818
rect 24032 9766 24046 9818
rect 24070 9766 24084 9818
rect 24084 9766 24096 9818
rect 24096 9766 24126 9818
rect 24150 9766 24160 9818
rect 24160 9766 24206 9818
rect 23910 9764 23966 9766
rect 23990 9764 24046 9766
rect 24070 9764 24126 9766
rect 24150 9764 24206 9766
rect 25502 14476 25558 14512
rect 25502 14456 25504 14476
rect 25504 14456 25556 14476
rect 25556 14456 25558 14476
rect 25778 14456 25834 14512
rect 25778 12724 25780 12744
rect 25780 12724 25832 12744
rect 25832 12724 25834 12744
rect 25778 12688 25834 12724
rect 26238 13776 26294 13832
rect 26882 14476 26938 14512
rect 26882 14456 26884 14476
rect 26884 14456 26936 14476
rect 26936 14456 26938 14476
rect 26146 12280 26202 12336
rect 25410 11600 25466 11656
rect 27268 16890 27324 16892
rect 27348 16890 27404 16892
rect 27428 16890 27484 16892
rect 27508 16890 27564 16892
rect 27268 16838 27314 16890
rect 27314 16838 27324 16890
rect 27348 16838 27378 16890
rect 27378 16838 27390 16890
rect 27390 16838 27404 16890
rect 27428 16838 27442 16890
rect 27442 16838 27454 16890
rect 27454 16838 27484 16890
rect 27508 16838 27518 16890
rect 27518 16838 27564 16890
rect 27268 16836 27324 16838
rect 27348 16836 27404 16838
rect 27428 16836 27484 16838
rect 27508 16836 27564 16838
rect 27268 15802 27324 15804
rect 27348 15802 27404 15804
rect 27428 15802 27484 15804
rect 27508 15802 27564 15804
rect 27268 15750 27314 15802
rect 27314 15750 27324 15802
rect 27348 15750 27378 15802
rect 27378 15750 27390 15802
rect 27390 15750 27404 15802
rect 27428 15750 27442 15802
rect 27442 15750 27454 15802
rect 27454 15750 27484 15802
rect 27508 15750 27518 15802
rect 27518 15750 27564 15802
rect 27268 15748 27324 15750
rect 27348 15748 27404 15750
rect 27428 15748 27484 15750
rect 27508 15748 27564 15750
rect 27268 14714 27324 14716
rect 27348 14714 27404 14716
rect 27428 14714 27484 14716
rect 27508 14714 27564 14716
rect 27268 14662 27314 14714
rect 27314 14662 27324 14714
rect 27348 14662 27378 14714
rect 27378 14662 27390 14714
rect 27390 14662 27404 14714
rect 27428 14662 27442 14714
rect 27442 14662 27454 14714
rect 27454 14662 27484 14714
rect 27508 14662 27518 14714
rect 27518 14662 27564 14714
rect 27268 14660 27324 14662
rect 27348 14660 27404 14662
rect 27428 14660 27484 14662
rect 27508 14660 27564 14662
rect 27158 13776 27214 13832
rect 27268 13626 27324 13628
rect 27348 13626 27404 13628
rect 27428 13626 27484 13628
rect 27508 13626 27564 13628
rect 27268 13574 27314 13626
rect 27314 13574 27324 13626
rect 27348 13574 27378 13626
rect 27378 13574 27390 13626
rect 27390 13574 27404 13626
rect 27428 13574 27442 13626
rect 27442 13574 27454 13626
rect 27454 13574 27484 13626
rect 27508 13574 27518 13626
rect 27518 13574 27564 13626
rect 27268 13572 27324 13574
rect 27348 13572 27404 13574
rect 27428 13572 27484 13574
rect 27508 13572 27564 13574
rect 27268 12538 27324 12540
rect 27348 12538 27404 12540
rect 27428 12538 27484 12540
rect 27508 12538 27564 12540
rect 27268 12486 27314 12538
rect 27314 12486 27324 12538
rect 27348 12486 27378 12538
rect 27378 12486 27390 12538
rect 27390 12486 27404 12538
rect 27428 12486 27442 12538
rect 27442 12486 27454 12538
rect 27454 12486 27484 12538
rect 27508 12486 27518 12538
rect 27518 12486 27564 12538
rect 27268 12484 27324 12486
rect 27348 12484 27404 12486
rect 27428 12484 27484 12486
rect 27508 12484 27564 12486
rect 27268 11450 27324 11452
rect 27348 11450 27404 11452
rect 27428 11450 27484 11452
rect 27508 11450 27564 11452
rect 27268 11398 27314 11450
rect 27314 11398 27324 11450
rect 27348 11398 27378 11450
rect 27378 11398 27390 11450
rect 27390 11398 27404 11450
rect 27428 11398 27442 11450
rect 27442 11398 27454 11450
rect 27454 11398 27484 11450
rect 27508 11398 27518 11450
rect 27518 11398 27564 11450
rect 27268 11396 27324 11398
rect 27348 11396 27404 11398
rect 27428 11396 27484 11398
rect 27508 11396 27564 11398
rect 24398 9152 24454 9208
rect 24122 8900 24178 8936
rect 24122 8880 24124 8900
rect 24124 8880 24176 8900
rect 24176 8880 24178 8900
rect 23910 8730 23966 8732
rect 23990 8730 24046 8732
rect 24070 8730 24126 8732
rect 24150 8730 24206 8732
rect 23910 8678 23956 8730
rect 23956 8678 23966 8730
rect 23990 8678 24020 8730
rect 24020 8678 24032 8730
rect 24032 8678 24046 8730
rect 24070 8678 24084 8730
rect 24084 8678 24096 8730
rect 24096 8678 24126 8730
rect 24150 8678 24160 8730
rect 24160 8678 24206 8730
rect 23910 8676 23966 8678
rect 23990 8676 24046 8678
rect 24070 8676 24126 8678
rect 24150 8676 24206 8678
rect 24030 8084 24086 8120
rect 24030 8064 24032 8084
rect 24032 8064 24084 8084
rect 24084 8064 24086 8084
rect 24398 8064 24454 8120
rect 24674 8508 24676 8528
rect 24676 8508 24728 8528
rect 24728 8508 24730 8528
rect 24674 8472 24730 8508
rect 25042 9152 25098 9208
rect 24674 8200 24730 8256
rect 24214 7948 24270 7984
rect 24214 7928 24216 7948
rect 24216 7928 24268 7948
rect 24268 7928 24270 7948
rect 24582 7928 24638 7984
rect 23910 7642 23966 7644
rect 23990 7642 24046 7644
rect 24070 7642 24126 7644
rect 24150 7642 24206 7644
rect 23910 7590 23956 7642
rect 23956 7590 23966 7642
rect 23990 7590 24020 7642
rect 24020 7590 24032 7642
rect 24032 7590 24046 7642
rect 24070 7590 24084 7642
rect 24084 7590 24096 7642
rect 24096 7590 24126 7642
rect 24150 7590 24160 7642
rect 24160 7590 24206 7642
rect 23910 7588 23966 7590
rect 23990 7588 24046 7590
rect 24070 7588 24126 7590
rect 24150 7588 24206 7590
rect 23910 6554 23966 6556
rect 23990 6554 24046 6556
rect 24070 6554 24126 6556
rect 24150 6554 24206 6556
rect 23910 6502 23956 6554
rect 23956 6502 23966 6554
rect 23990 6502 24020 6554
rect 24020 6502 24032 6554
rect 24032 6502 24046 6554
rect 24070 6502 24084 6554
rect 24084 6502 24096 6554
rect 24096 6502 24126 6554
rect 24150 6502 24160 6554
rect 24160 6502 24206 6554
rect 23910 6500 23966 6502
rect 23990 6500 24046 6502
rect 24070 6500 24126 6502
rect 24150 6500 24206 6502
rect 27268 10362 27324 10364
rect 27348 10362 27404 10364
rect 27428 10362 27484 10364
rect 27508 10362 27564 10364
rect 27268 10310 27314 10362
rect 27314 10310 27324 10362
rect 27348 10310 27378 10362
rect 27378 10310 27390 10362
rect 27390 10310 27404 10362
rect 27428 10310 27442 10362
rect 27442 10310 27454 10362
rect 27454 10310 27484 10362
rect 27508 10310 27518 10362
rect 27518 10310 27564 10362
rect 27268 10308 27324 10310
rect 27348 10308 27404 10310
rect 27428 10308 27484 10310
rect 27508 10308 27564 10310
rect 27268 9274 27324 9276
rect 27348 9274 27404 9276
rect 27428 9274 27484 9276
rect 27508 9274 27564 9276
rect 27268 9222 27314 9274
rect 27314 9222 27324 9274
rect 27348 9222 27378 9274
rect 27378 9222 27390 9274
rect 27390 9222 27404 9274
rect 27428 9222 27442 9274
rect 27442 9222 27454 9274
rect 27454 9222 27484 9274
rect 27508 9222 27518 9274
rect 27518 9222 27564 9274
rect 27268 9220 27324 9222
rect 27348 9220 27404 9222
rect 27428 9220 27484 9222
rect 27508 9220 27564 9222
rect 25594 7928 25650 7984
rect 27268 8186 27324 8188
rect 27348 8186 27404 8188
rect 27428 8186 27484 8188
rect 27508 8186 27564 8188
rect 27268 8134 27314 8186
rect 27314 8134 27324 8186
rect 27348 8134 27378 8186
rect 27378 8134 27390 8186
rect 27390 8134 27404 8186
rect 27428 8134 27442 8186
rect 27442 8134 27454 8186
rect 27454 8134 27484 8186
rect 27508 8134 27518 8186
rect 27518 8134 27564 8186
rect 27268 8132 27324 8134
rect 27348 8132 27404 8134
rect 27428 8132 27484 8134
rect 27508 8132 27564 8134
rect 27268 7098 27324 7100
rect 27348 7098 27404 7100
rect 27428 7098 27484 7100
rect 27508 7098 27564 7100
rect 27268 7046 27314 7098
rect 27314 7046 27324 7098
rect 27348 7046 27378 7098
rect 27378 7046 27390 7098
rect 27390 7046 27404 7098
rect 27428 7046 27442 7098
rect 27442 7046 27454 7098
rect 27454 7046 27484 7098
rect 27508 7046 27518 7098
rect 27518 7046 27564 7098
rect 27268 7044 27324 7046
rect 27348 7044 27404 7046
rect 27428 7044 27484 7046
rect 27508 7044 27564 7046
rect 27268 6010 27324 6012
rect 27348 6010 27404 6012
rect 27428 6010 27484 6012
rect 27508 6010 27564 6012
rect 27268 5958 27314 6010
rect 27314 5958 27324 6010
rect 27348 5958 27378 6010
rect 27378 5958 27390 6010
rect 27390 5958 27404 6010
rect 27428 5958 27442 6010
rect 27442 5958 27454 6010
rect 27454 5958 27484 6010
rect 27508 5958 27518 6010
rect 27518 5958 27564 6010
rect 27268 5956 27324 5958
rect 27348 5956 27404 5958
rect 27428 5956 27484 5958
rect 27508 5956 27564 5958
rect 23910 5466 23966 5468
rect 23990 5466 24046 5468
rect 24070 5466 24126 5468
rect 24150 5466 24206 5468
rect 23910 5414 23956 5466
rect 23956 5414 23966 5466
rect 23990 5414 24020 5466
rect 24020 5414 24032 5466
rect 24032 5414 24046 5466
rect 24070 5414 24084 5466
rect 24084 5414 24096 5466
rect 24096 5414 24126 5466
rect 24150 5414 24160 5466
rect 24160 5414 24206 5466
rect 23910 5412 23966 5414
rect 23990 5412 24046 5414
rect 24070 5412 24126 5414
rect 24150 5412 24206 5414
rect 23910 4378 23966 4380
rect 23990 4378 24046 4380
rect 24070 4378 24126 4380
rect 24150 4378 24206 4380
rect 23910 4326 23956 4378
rect 23956 4326 23966 4378
rect 23990 4326 24020 4378
rect 24020 4326 24032 4378
rect 24032 4326 24046 4378
rect 24070 4326 24084 4378
rect 24084 4326 24096 4378
rect 24096 4326 24126 4378
rect 24150 4326 24160 4378
rect 24160 4326 24206 4378
rect 23910 4324 23966 4326
rect 23990 4324 24046 4326
rect 24070 4324 24126 4326
rect 24150 4324 24206 4326
rect 27268 4922 27324 4924
rect 27348 4922 27404 4924
rect 27428 4922 27484 4924
rect 27508 4922 27564 4924
rect 27268 4870 27314 4922
rect 27314 4870 27324 4922
rect 27348 4870 27378 4922
rect 27378 4870 27390 4922
rect 27390 4870 27404 4922
rect 27428 4870 27442 4922
rect 27442 4870 27454 4922
rect 27454 4870 27484 4922
rect 27508 4870 27518 4922
rect 27518 4870 27564 4922
rect 27268 4868 27324 4870
rect 27348 4868 27404 4870
rect 27428 4868 27484 4870
rect 27508 4868 27564 4870
rect 27268 3834 27324 3836
rect 27348 3834 27404 3836
rect 27428 3834 27484 3836
rect 27508 3834 27564 3836
rect 27268 3782 27314 3834
rect 27314 3782 27324 3834
rect 27348 3782 27378 3834
rect 27378 3782 27390 3834
rect 27390 3782 27404 3834
rect 27428 3782 27442 3834
rect 27442 3782 27454 3834
rect 27454 3782 27484 3834
rect 27508 3782 27518 3834
rect 27518 3782 27564 3834
rect 27268 3780 27324 3782
rect 27348 3780 27404 3782
rect 27428 3780 27484 3782
rect 27508 3780 27564 3782
rect 23910 3290 23966 3292
rect 23990 3290 24046 3292
rect 24070 3290 24126 3292
rect 24150 3290 24206 3292
rect 23910 3238 23956 3290
rect 23956 3238 23966 3290
rect 23990 3238 24020 3290
rect 24020 3238 24032 3290
rect 24032 3238 24046 3290
rect 24070 3238 24084 3290
rect 24084 3238 24096 3290
rect 24096 3238 24126 3290
rect 24150 3238 24160 3290
rect 24160 3238 24206 3290
rect 23910 3236 23966 3238
rect 23990 3236 24046 3238
rect 24070 3236 24126 3238
rect 24150 3236 24206 3238
rect 20552 2746 20608 2748
rect 20632 2746 20688 2748
rect 20712 2746 20768 2748
rect 20792 2746 20848 2748
rect 20552 2694 20598 2746
rect 20598 2694 20608 2746
rect 20632 2694 20662 2746
rect 20662 2694 20674 2746
rect 20674 2694 20688 2746
rect 20712 2694 20726 2746
rect 20726 2694 20738 2746
rect 20738 2694 20768 2746
rect 20792 2694 20802 2746
rect 20802 2694 20848 2746
rect 20552 2692 20608 2694
rect 20632 2692 20688 2694
rect 20712 2692 20768 2694
rect 20792 2692 20848 2694
rect 27268 2746 27324 2748
rect 27348 2746 27404 2748
rect 27428 2746 27484 2748
rect 27508 2746 27564 2748
rect 20626 2488 20682 2544
rect 27268 2694 27314 2746
rect 27314 2694 27324 2746
rect 27348 2694 27378 2746
rect 27378 2694 27390 2746
rect 27390 2694 27404 2746
rect 27428 2694 27442 2746
rect 27442 2694 27454 2746
rect 27454 2694 27484 2746
rect 27508 2694 27518 2746
rect 27518 2694 27564 2746
rect 27268 2692 27324 2694
rect 27348 2692 27404 2694
rect 27428 2692 27484 2694
rect 27508 2692 27564 2694
rect 20552 1658 20608 1660
rect 20632 1658 20688 1660
rect 20712 1658 20768 1660
rect 20792 1658 20848 1660
rect 20552 1606 20598 1658
rect 20598 1606 20608 1658
rect 20632 1606 20662 1658
rect 20662 1606 20674 1658
rect 20674 1606 20688 1658
rect 20712 1606 20726 1658
rect 20726 1606 20738 1658
rect 20738 1606 20768 1658
rect 20792 1606 20802 1658
rect 20802 1606 20848 1658
rect 20552 1604 20608 1606
rect 20632 1604 20688 1606
rect 20712 1604 20768 1606
rect 20792 1604 20848 1606
rect 20552 570 20608 572
rect 20632 570 20688 572
rect 20712 570 20768 572
rect 20792 570 20848 572
rect 20552 518 20598 570
rect 20598 518 20608 570
rect 20632 518 20662 570
rect 20662 518 20674 570
rect 20674 518 20688 570
rect 20712 518 20726 570
rect 20726 518 20738 570
rect 20738 518 20768 570
rect 20792 518 20802 570
rect 20802 518 20848 570
rect 20552 516 20608 518
rect 20632 516 20688 518
rect 20712 516 20768 518
rect 20792 516 20848 518
rect 23910 2202 23966 2204
rect 23990 2202 24046 2204
rect 24070 2202 24126 2204
rect 24150 2202 24206 2204
rect 23910 2150 23956 2202
rect 23956 2150 23966 2202
rect 23990 2150 24020 2202
rect 24020 2150 24032 2202
rect 24032 2150 24046 2202
rect 24070 2150 24084 2202
rect 24084 2150 24096 2202
rect 24096 2150 24126 2202
rect 24150 2150 24160 2202
rect 24160 2150 24206 2202
rect 23910 2148 23966 2150
rect 23990 2148 24046 2150
rect 24070 2148 24126 2150
rect 24150 2148 24206 2150
rect 23910 1114 23966 1116
rect 23990 1114 24046 1116
rect 24070 1114 24126 1116
rect 24150 1114 24206 1116
rect 23910 1062 23956 1114
rect 23956 1062 23966 1114
rect 23990 1062 24020 1114
rect 24020 1062 24032 1114
rect 24032 1062 24046 1114
rect 24070 1062 24084 1114
rect 24084 1062 24096 1114
rect 24096 1062 24126 1114
rect 24150 1062 24160 1114
rect 24160 1062 24206 1114
rect 23910 1060 23966 1062
rect 23990 1060 24046 1062
rect 24070 1060 24126 1062
rect 24150 1060 24206 1062
rect 27268 1658 27324 1660
rect 27348 1658 27404 1660
rect 27428 1658 27484 1660
rect 27508 1658 27564 1660
rect 27268 1606 27314 1658
rect 27314 1606 27324 1658
rect 27348 1606 27378 1658
rect 27378 1606 27390 1658
rect 27390 1606 27404 1658
rect 27428 1606 27442 1658
rect 27442 1606 27454 1658
rect 27454 1606 27484 1658
rect 27508 1606 27518 1658
rect 27518 1606 27564 1658
rect 27268 1604 27324 1606
rect 27348 1604 27404 1606
rect 27428 1604 27484 1606
rect 27508 1604 27564 1606
rect 27268 570 27324 572
rect 27348 570 27404 572
rect 27428 570 27484 572
rect 27508 570 27564 572
rect 27268 518 27314 570
rect 27314 518 27324 570
rect 27348 518 27378 570
rect 27378 518 27390 570
rect 27390 518 27404 570
rect 27428 518 27442 570
rect 27442 518 27454 570
rect 27454 518 27484 570
rect 27508 518 27518 570
rect 27518 518 27564 570
rect 27268 516 27324 518
rect 27348 516 27404 518
rect 27428 516 27484 518
rect 27508 516 27564 518
<< metal3 >>
rect 3752 17440 4068 17441
rect 3752 17376 3758 17440
rect 3822 17376 3838 17440
rect 3902 17376 3918 17440
rect 3982 17376 3998 17440
rect 4062 17376 4068 17440
rect 3752 17375 4068 17376
rect 10468 17440 10784 17441
rect 10468 17376 10474 17440
rect 10538 17376 10554 17440
rect 10618 17376 10634 17440
rect 10698 17376 10714 17440
rect 10778 17376 10784 17440
rect 10468 17375 10784 17376
rect 17184 17440 17500 17441
rect 17184 17376 17190 17440
rect 17254 17376 17270 17440
rect 17334 17376 17350 17440
rect 17414 17376 17430 17440
rect 17494 17376 17500 17440
rect 17184 17375 17500 17376
rect 23900 17440 24216 17441
rect 23900 17376 23906 17440
rect 23970 17376 23986 17440
rect 24050 17376 24066 17440
rect 24130 17376 24146 17440
rect 24210 17376 24216 17440
rect 23900 17375 24216 17376
rect 7110 16896 7426 16897
rect 7110 16832 7116 16896
rect 7180 16832 7196 16896
rect 7260 16832 7276 16896
rect 7340 16832 7356 16896
rect 7420 16832 7426 16896
rect 7110 16831 7426 16832
rect 13826 16896 14142 16897
rect 13826 16832 13832 16896
rect 13896 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14142 16896
rect 13826 16831 14142 16832
rect 20542 16896 20858 16897
rect 20542 16832 20548 16896
rect 20612 16832 20628 16896
rect 20692 16832 20708 16896
rect 20772 16832 20788 16896
rect 20852 16832 20858 16896
rect 20542 16831 20858 16832
rect 27258 16896 27574 16897
rect 27258 16832 27264 16896
rect 27328 16832 27344 16896
rect 27408 16832 27424 16896
rect 27488 16832 27504 16896
rect 27568 16832 27574 16896
rect 27258 16831 27574 16832
rect 12433 16690 12499 16693
rect 12566 16690 12572 16692
rect 12433 16688 12572 16690
rect 12433 16632 12438 16688
rect 12494 16632 12572 16688
rect 12433 16630 12572 16632
rect 12433 16627 12499 16630
rect 12566 16628 12572 16630
rect 12636 16628 12642 16692
rect 16798 16628 16804 16692
rect 16868 16690 16874 16692
rect 17125 16690 17191 16693
rect 16868 16688 17191 16690
rect 16868 16632 17130 16688
rect 17186 16632 17191 16688
rect 16868 16630 17191 16632
rect 16868 16628 16874 16630
rect 17125 16627 17191 16630
rect 3752 16352 4068 16353
rect 3752 16288 3758 16352
rect 3822 16288 3838 16352
rect 3902 16288 3918 16352
rect 3982 16288 3998 16352
rect 4062 16288 4068 16352
rect 3752 16287 4068 16288
rect 10468 16352 10784 16353
rect 10468 16288 10474 16352
rect 10538 16288 10554 16352
rect 10618 16288 10634 16352
rect 10698 16288 10714 16352
rect 10778 16288 10784 16352
rect 10468 16287 10784 16288
rect 17184 16352 17500 16353
rect 17184 16288 17190 16352
rect 17254 16288 17270 16352
rect 17334 16288 17350 16352
rect 17414 16288 17430 16352
rect 17494 16288 17500 16352
rect 17184 16287 17500 16288
rect 23900 16352 24216 16353
rect 23900 16288 23906 16352
rect 23970 16288 23986 16352
rect 24050 16288 24066 16352
rect 24130 16288 24146 16352
rect 24210 16288 24216 16352
rect 23900 16287 24216 16288
rect 12157 16146 12223 16149
rect 14641 16146 14707 16149
rect 12157 16144 14707 16146
rect 12157 16088 12162 16144
rect 12218 16088 14646 16144
rect 14702 16088 14707 16144
rect 12157 16086 14707 16088
rect 12157 16083 12223 16086
rect 14641 16083 14707 16086
rect 9765 16010 9831 16013
rect 11973 16010 12039 16013
rect 9765 16008 12039 16010
rect 9765 15952 9770 16008
rect 9826 15952 11978 16008
rect 12034 15952 12039 16008
rect 9765 15950 12039 15952
rect 9765 15947 9831 15950
rect 11973 15947 12039 15950
rect 12709 16010 12775 16013
rect 14181 16010 14247 16013
rect 12709 16008 14247 16010
rect 12709 15952 12714 16008
rect 12770 15952 14186 16008
rect 14242 15952 14247 16008
rect 12709 15950 14247 15952
rect 12709 15947 12775 15950
rect 14181 15947 14247 15950
rect 7110 15808 7426 15809
rect 7110 15744 7116 15808
rect 7180 15744 7196 15808
rect 7260 15744 7276 15808
rect 7340 15744 7356 15808
rect 7420 15744 7426 15808
rect 7110 15743 7426 15744
rect 13826 15808 14142 15809
rect 13826 15744 13832 15808
rect 13896 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14142 15808
rect 13826 15743 14142 15744
rect 20542 15808 20858 15809
rect 20542 15744 20548 15808
rect 20612 15744 20628 15808
rect 20692 15744 20708 15808
rect 20772 15744 20788 15808
rect 20852 15744 20858 15808
rect 20542 15743 20858 15744
rect 27258 15808 27574 15809
rect 27258 15744 27264 15808
rect 27328 15744 27344 15808
rect 27408 15744 27424 15808
rect 27488 15744 27504 15808
rect 27568 15744 27574 15808
rect 27258 15743 27574 15744
rect 8477 15602 8543 15605
rect 17953 15602 18019 15605
rect 22829 15602 22895 15605
rect 8477 15600 22895 15602
rect 8477 15544 8482 15600
rect 8538 15544 17958 15600
rect 18014 15544 22834 15600
rect 22890 15544 22895 15600
rect 8477 15542 22895 15544
rect 8477 15539 8543 15542
rect 17953 15539 18019 15542
rect 22829 15539 22895 15542
rect 3752 15264 4068 15265
rect 3752 15200 3758 15264
rect 3822 15200 3838 15264
rect 3902 15200 3918 15264
rect 3982 15200 3998 15264
rect 4062 15200 4068 15264
rect 3752 15199 4068 15200
rect 10468 15264 10784 15265
rect 10468 15200 10474 15264
rect 10538 15200 10554 15264
rect 10618 15200 10634 15264
rect 10698 15200 10714 15264
rect 10778 15200 10784 15264
rect 10468 15199 10784 15200
rect 17184 15264 17500 15265
rect 17184 15200 17190 15264
rect 17254 15200 17270 15264
rect 17334 15200 17350 15264
rect 17414 15200 17430 15264
rect 17494 15200 17500 15264
rect 17184 15199 17500 15200
rect 23900 15264 24216 15265
rect 23900 15200 23906 15264
rect 23970 15200 23986 15264
rect 24050 15200 24066 15264
rect 24130 15200 24146 15264
rect 24210 15200 24216 15264
rect 23900 15199 24216 15200
rect 19425 14922 19491 14925
rect 20805 14922 20871 14925
rect 21909 14922 21975 14925
rect 19425 14920 21975 14922
rect 19425 14864 19430 14920
rect 19486 14864 20810 14920
rect 20866 14864 21914 14920
rect 21970 14864 21975 14920
rect 19425 14862 21975 14864
rect 19425 14859 19491 14862
rect 20805 14859 20871 14862
rect 21909 14859 21975 14862
rect 7110 14720 7426 14721
rect 7110 14656 7116 14720
rect 7180 14656 7196 14720
rect 7260 14656 7276 14720
rect 7340 14656 7356 14720
rect 7420 14656 7426 14720
rect 7110 14655 7426 14656
rect 13826 14720 14142 14721
rect 13826 14656 13832 14720
rect 13896 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14142 14720
rect 13826 14655 14142 14656
rect 20542 14720 20858 14721
rect 20542 14656 20548 14720
rect 20612 14656 20628 14720
rect 20692 14656 20708 14720
rect 20772 14656 20788 14720
rect 20852 14656 20858 14720
rect 20542 14655 20858 14656
rect 27258 14720 27574 14721
rect 27258 14656 27264 14720
rect 27328 14656 27344 14720
rect 27408 14656 27424 14720
rect 27488 14656 27504 14720
rect 27568 14656 27574 14720
rect 27258 14655 27574 14656
rect 22921 14514 22987 14517
rect 25497 14514 25563 14517
rect 25773 14514 25839 14517
rect 26877 14514 26943 14517
rect 22921 14512 26943 14514
rect 22921 14456 22926 14512
rect 22982 14456 25502 14512
rect 25558 14456 25778 14512
rect 25834 14456 26882 14512
rect 26938 14456 26943 14512
rect 22921 14454 26943 14456
rect 22921 14451 22987 14454
rect 25497 14451 25563 14454
rect 25773 14451 25839 14454
rect 26877 14451 26943 14454
rect 3752 14176 4068 14177
rect 3752 14112 3758 14176
rect 3822 14112 3838 14176
rect 3902 14112 3918 14176
rect 3982 14112 3998 14176
rect 4062 14112 4068 14176
rect 3752 14111 4068 14112
rect 10468 14176 10784 14177
rect 10468 14112 10474 14176
rect 10538 14112 10554 14176
rect 10618 14112 10634 14176
rect 10698 14112 10714 14176
rect 10778 14112 10784 14176
rect 10468 14111 10784 14112
rect 17184 14176 17500 14177
rect 17184 14112 17190 14176
rect 17254 14112 17270 14176
rect 17334 14112 17350 14176
rect 17414 14112 17430 14176
rect 17494 14112 17500 14176
rect 17184 14111 17500 14112
rect 23900 14176 24216 14177
rect 23900 14112 23906 14176
rect 23970 14112 23986 14176
rect 24050 14112 24066 14176
rect 24130 14112 24146 14176
rect 24210 14112 24216 14176
rect 23900 14111 24216 14112
rect 26233 13834 26299 13837
rect 27153 13834 27219 13837
rect 26233 13832 27219 13834
rect 26233 13776 26238 13832
rect 26294 13776 27158 13832
rect 27214 13776 27219 13832
rect 26233 13774 27219 13776
rect 26233 13771 26299 13774
rect 27153 13771 27219 13774
rect 7110 13632 7426 13633
rect 7110 13568 7116 13632
rect 7180 13568 7196 13632
rect 7260 13568 7276 13632
rect 7340 13568 7356 13632
rect 7420 13568 7426 13632
rect 7110 13567 7426 13568
rect 13826 13632 14142 13633
rect 13826 13568 13832 13632
rect 13896 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14142 13632
rect 13826 13567 14142 13568
rect 20542 13632 20858 13633
rect 20542 13568 20548 13632
rect 20612 13568 20628 13632
rect 20692 13568 20708 13632
rect 20772 13568 20788 13632
rect 20852 13568 20858 13632
rect 20542 13567 20858 13568
rect 27258 13632 27574 13633
rect 27258 13568 27264 13632
rect 27328 13568 27344 13632
rect 27408 13568 27424 13632
rect 27488 13568 27504 13632
rect 27568 13568 27574 13632
rect 27258 13567 27574 13568
rect 3601 13562 3667 13565
rect 4337 13562 4403 13565
rect 3601 13560 4403 13562
rect 3601 13504 3606 13560
rect 3662 13504 4342 13560
rect 4398 13504 4403 13560
rect 3601 13502 4403 13504
rect 3601 13499 3667 13502
rect 4337 13499 4403 13502
rect 17769 13562 17835 13565
rect 19241 13562 19307 13565
rect 17769 13560 19307 13562
rect 17769 13504 17774 13560
rect 17830 13504 19246 13560
rect 19302 13504 19307 13560
rect 17769 13502 19307 13504
rect 17769 13499 17835 13502
rect 19241 13499 19307 13502
rect 3785 13426 3851 13429
rect 4521 13426 4587 13429
rect 4797 13426 4863 13429
rect 3785 13424 4863 13426
rect 3785 13368 3790 13424
rect 3846 13368 4526 13424
rect 4582 13368 4802 13424
rect 4858 13368 4863 13424
rect 3785 13366 4863 13368
rect 3785 13363 3851 13366
rect 4521 13363 4587 13366
rect 4797 13363 4863 13366
rect 5809 13426 5875 13429
rect 8845 13426 8911 13429
rect 5809 13424 8911 13426
rect 5809 13368 5814 13424
rect 5870 13368 8850 13424
rect 8906 13368 8911 13424
rect 5809 13366 8911 13368
rect 5809 13363 5875 13366
rect 8845 13363 8911 13366
rect 10961 13426 11027 13429
rect 20345 13426 20411 13429
rect 10961 13424 20411 13426
rect 10961 13368 10966 13424
rect 11022 13368 20350 13424
rect 20406 13368 20411 13424
rect 10961 13366 20411 13368
rect 10961 13363 11027 13366
rect 20345 13363 20411 13366
rect 3752 13088 4068 13089
rect 3752 13024 3758 13088
rect 3822 13024 3838 13088
rect 3902 13024 3918 13088
rect 3982 13024 3998 13088
rect 4062 13024 4068 13088
rect 3752 13023 4068 13024
rect 10468 13088 10784 13089
rect 10468 13024 10474 13088
rect 10538 13024 10554 13088
rect 10618 13024 10634 13088
rect 10698 13024 10714 13088
rect 10778 13024 10784 13088
rect 10468 13023 10784 13024
rect 17184 13088 17500 13089
rect 17184 13024 17190 13088
rect 17254 13024 17270 13088
rect 17334 13024 17350 13088
rect 17414 13024 17430 13088
rect 17494 13024 17500 13088
rect 17184 13023 17500 13024
rect 23900 13088 24216 13089
rect 23900 13024 23906 13088
rect 23970 13024 23986 13088
rect 24050 13024 24066 13088
rect 24130 13024 24146 13088
rect 24210 13024 24216 13088
rect 23900 13023 24216 13024
rect 7557 12882 7623 12885
rect 20161 12882 20227 12885
rect 20621 12882 20687 12885
rect 7557 12880 20687 12882
rect 7557 12824 7562 12880
rect 7618 12824 20166 12880
rect 20222 12824 20626 12880
rect 20682 12824 20687 12880
rect 7557 12822 20687 12824
rect 7557 12819 7623 12822
rect 20161 12819 20227 12822
rect 20621 12819 20687 12822
rect 24301 12746 24367 12749
rect 25773 12746 25839 12749
rect 24301 12744 25839 12746
rect 24301 12688 24306 12744
rect 24362 12688 25778 12744
rect 25834 12688 25839 12744
rect 24301 12686 25839 12688
rect 24301 12683 24367 12686
rect 25773 12683 25839 12686
rect 7110 12544 7426 12545
rect 7110 12480 7116 12544
rect 7180 12480 7196 12544
rect 7260 12480 7276 12544
rect 7340 12480 7356 12544
rect 7420 12480 7426 12544
rect 7110 12479 7426 12480
rect 13826 12544 14142 12545
rect 13826 12480 13832 12544
rect 13896 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14142 12544
rect 13826 12479 14142 12480
rect 20542 12544 20858 12545
rect 20542 12480 20548 12544
rect 20612 12480 20628 12544
rect 20692 12480 20708 12544
rect 20772 12480 20788 12544
rect 20852 12480 20858 12544
rect 20542 12479 20858 12480
rect 27258 12544 27574 12545
rect 27258 12480 27264 12544
rect 27328 12480 27344 12544
rect 27408 12480 27424 12544
rect 27488 12480 27504 12544
rect 27568 12480 27574 12544
rect 27258 12479 27574 12480
rect 6637 12338 6703 12341
rect 10961 12340 11027 12341
rect 10910 12338 10916 12340
rect 6637 12336 10916 12338
rect 10980 12336 11027 12340
rect 6637 12280 6642 12336
rect 6698 12280 10916 12336
rect 11022 12280 11027 12336
rect 6637 12278 10916 12280
rect 6637 12275 6703 12278
rect 10910 12276 10916 12278
rect 10980 12276 11027 12280
rect 10961 12275 11027 12276
rect 15745 12338 15811 12341
rect 18597 12338 18663 12341
rect 15745 12336 18663 12338
rect 15745 12280 15750 12336
rect 15806 12280 18602 12336
rect 18658 12280 18663 12336
rect 15745 12278 18663 12280
rect 15745 12275 15811 12278
rect 18597 12275 18663 12278
rect 26141 12340 26207 12341
rect 26141 12336 26188 12340
rect 26252 12338 26258 12340
rect 26141 12280 26146 12336
rect 26141 12276 26188 12280
rect 26252 12278 26298 12338
rect 26252 12276 26258 12278
rect 26141 12275 26207 12276
rect 13445 12202 13511 12205
rect 15009 12202 15075 12205
rect 13445 12200 15075 12202
rect 13445 12144 13450 12200
rect 13506 12144 15014 12200
rect 15070 12144 15075 12200
rect 13445 12142 15075 12144
rect 13445 12139 13511 12142
rect 15009 12139 15075 12142
rect 3752 12000 4068 12001
rect 3752 11936 3758 12000
rect 3822 11936 3838 12000
rect 3902 11936 3918 12000
rect 3982 11936 3998 12000
rect 4062 11936 4068 12000
rect 3752 11935 4068 11936
rect 10468 12000 10784 12001
rect 10468 11936 10474 12000
rect 10538 11936 10554 12000
rect 10618 11936 10634 12000
rect 10698 11936 10714 12000
rect 10778 11936 10784 12000
rect 10468 11935 10784 11936
rect 17184 12000 17500 12001
rect 17184 11936 17190 12000
rect 17254 11936 17270 12000
rect 17334 11936 17350 12000
rect 17414 11936 17430 12000
rect 17494 11936 17500 12000
rect 17184 11935 17500 11936
rect 23900 12000 24216 12001
rect 23900 11936 23906 12000
rect 23970 11936 23986 12000
rect 24050 11936 24066 12000
rect 24130 11936 24146 12000
rect 24210 11936 24216 12000
rect 23900 11935 24216 11936
rect 10041 11658 10107 11661
rect 25405 11658 25471 11661
rect 10041 11656 25471 11658
rect 10041 11600 10046 11656
rect 10102 11600 25410 11656
rect 25466 11600 25471 11656
rect 10041 11598 25471 11600
rect 10041 11595 10107 11598
rect 25405 11595 25471 11598
rect 7110 11456 7426 11457
rect 7110 11392 7116 11456
rect 7180 11392 7196 11456
rect 7260 11392 7276 11456
rect 7340 11392 7356 11456
rect 7420 11392 7426 11456
rect 7110 11391 7426 11392
rect 13826 11456 14142 11457
rect 13826 11392 13832 11456
rect 13896 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14142 11456
rect 13826 11391 14142 11392
rect 20542 11456 20858 11457
rect 20542 11392 20548 11456
rect 20612 11392 20628 11456
rect 20692 11392 20708 11456
rect 20772 11392 20788 11456
rect 20852 11392 20858 11456
rect 20542 11391 20858 11392
rect 27258 11456 27574 11457
rect 27258 11392 27264 11456
rect 27328 11392 27344 11456
rect 27408 11392 27424 11456
rect 27488 11392 27504 11456
rect 27568 11392 27574 11456
rect 27258 11391 27574 11392
rect 3752 10912 4068 10913
rect 3752 10848 3758 10912
rect 3822 10848 3838 10912
rect 3902 10848 3918 10912
rect 3982 10848 3998 10912
rect 4062 10848 4068 10912
rect 3752 10847 4068 10848
rect 10468 10912 10784 10913
rect 10468 10848 10474 10912
rect 10538 10848 10554 10912
rect 10618 10848 10634 10912
rect 10698 10848 10714 10912
rect 10778 10848 10784 10912
rect 10468 10847 10784 10848
rect 17184 10912 17500 10913
rect 17184 10848 17190 10912
rect 17254 10848 17270 10912
rect 17334 10848 17350 10912
rect 17414 10848 17430 10912
rect 17494 10848 17500 10912
rect 17184 10847 17500 10848
rect 23900 10912 24216 10913
rect 23900 10848 23906 10912
rect 23970 10848 23986 10912
rect 24050 10848 24066 10912
rect 24130 10848 24146 10912
rect 24210 10848 24216 10912
rect 23900 10847 24216 10848
rect 7110 10368 7426 10369
rect 7110 10304 7116 10368
rect 7180 10304 7196 10368
rect 7260 10304 7276 10368
rect 7340 10304 7356 10368
rect 7420 10304 7426 10368
rect 7110 10303 7426 10304
rect 13826 10368 14142 10369
rect 13826 10304 13832 10368
rect 13896 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14142 10368
rect 13826 10303 14142 10304
rect 20542 10368 20858 10369
rect 20542 10304 20548 10368
rect 20612 10304 20628 10368
rect 20692 10304 20708 10368
rect 20772 10304 20788 10368
rect 20852 10304 20858 10368
rect 20542 10303 20858 10304
rect 27258 10368 27574 10369
rect 27258 10304 27264 10368
rect 27328 10304 27344 10368
rect 27408 10304 27424 10368
rect 27488 10304 27504 10368
rect 27568 10304 27574 10368
rect 27258 10303 27574 10304
rect 9857 10162 9923 10165
rect 18597 10162 18663 10165
rect 19057 10162 19123 10165
rect 9857 10160 19123 10162
rect 9857 10104 9862 10160
rect 9918 10104 18602 10160
rect 18658 10104 19062 10160
rect 19118 10104 19123 10160
rect 9857 10102 19123 10104
rect 9857 10099 9923 10102
rect 18597 10099 18663 10102
rect 19057 10099 19123 10102
rect 3752 9824 4068 9825
rect 3752 9760 3758 9824
rect 3822 9760 3838 9824
rect 3902 9760 3918 9824
rect 3982 9760 3998 9824
rect 4062 9760 4068 9824
rect 3752 9759 4068 9760
rect 10468 9824 10784 9825
rect 10468 9760 10474 9824
rect 10538 9760 10554 9824
rect 10618 9760 10634 9824
rect 10698 9760 10714 9824
rect 10778 9760 10784 9824
rect 10468 9759 10784 9760
rect 17184 9824 17500 9825
rect 17184 9760 17190 9824
rect 17254 9760 17270 9824
rect 17334 9760 17350 9824
rect 17414 9760 17430 9824
rect 17494 9760 17500 9824
rect 17184 9759 17500 9760
rect 23900 9824 24216 9825
rect 23900 9760 23906 9824
rect 23970 9760 23986 9824
rect 24050 9760 24066 9824
rect 24130 9760 24146 9824
rect 24210 9760 24216 9824
rect 23900 9759 24216 9760
rect 10910 9556 10916 9620
rect 10980 9618 10986 9620
rect 14273 9618 14339 9621
rect 10980 9616 14339 9618
rect 10980 9560 14278 9616
rect 14334 9560 14339 9616
rect 10980 9558 14339 9560
rect 10980 9556 10986 9558
rect 14273 9555 14339 9558
rect 16021 9482 16087 9485
rect 26182 9482 26188 9484
rect 16021 9480 26188 9482
rect 16021 9424 16026 9480
rect 16082 9424 26188 9480
rect 16021 9422 26188 9424
rect 16021 9419 16087 9422
rect 26182 9420 26188 9422
rect 26252 9420 26258 9484
rect 7110 9280 7426 9281
rect 7110 9216 7116 9280
rect 7180 9216 7196 9280
rect 7260 9216 7276 9280
rect 7340 9216 7356 9280
rect 7420 9216 7426 9280
rect 7110 9215 7426 9216
rect 13826 9280 14142 9281
rect 13826 9216 13832 9280
rect 13896 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14142 9280
rect 13826 9215 14142 9216
rect 20542 9280 20858 9281
rect 20542 9216 20548 9280
rect 20612 9216 20628 9280
rect 20692 9216 20708 9280
rect 20772 9216 20788 9280
rect 20852 9216 20858 9280
rect 20542 9215 20858 9216
rect 27258 9280 27574 9281
rect 27258 9216 27264 9280
rect 27328 9216 27344 9280
rect 27408 9216 27424 9280
rect 27488 9216 27504 9280
rect 27568 9216 27574 9280
rect 27258 9215 27574 9216
rect 9673 9210 9739 9213
rect 12433 9210 12499 9213
rect 13169 9210 13235 9213
rect 9673 9208 13235 9210
rect 9673 9152 9678 9208
rect 9734 9152 12438 9208
rect 12494 9152 13174 9208
rect 13230 9152 13235 9208
rect 9673 9150 13235 9152
rect 9673 9147 9739 9150
rect 12433 9147 12499 9150
rect 13169 9147 13235 9150
rect 24393 9210 24459 9213
rect 25037 9210 25103 9213
rect 24393 9208 25103 9210
rect 24393 9152 24398 9208
rect 24454 9152 25042 9208
rect 25098 9152 25103 9208
rect 24393 9150 25103 9152
rect 24393 9147 24459 9150
rect 25037 9147 25103 9150
rect 4429 9074 4495 9077
rect 18045 9074 18111 9077
rect 4429 9072 18111 9074
rect 4429 9016 4434 9072
rect 4490 9016 18050 9072
rect 18106 9016 18111 9072
rect 4429 9014 18111 9016
rect 4429 9011 4495 9014
rect 18045 9011 18111 9014
rect 8293 8940 8359 8941
rect 8293 8938 8340 8940
rect 8248 8936 8340 8938
rect 8404 8938 8410 8940
rect 9305 8938 9371 8941
rect 8404 8936 9371 8938
rect 8248 8880 8298 8936
rect 8404 8880 9310 8936
rect 9366 8880 9371 8936
rect 8248 8878 8340 8880
rect 8293 8876 8340 8878
rect 8404 8878 9371 8880
rect 8404 8876 8410 8878
rect 8293 8875 8359 8876
rect 9305 8875 9371 8878
rect 21357 8938 21423 8941
rect 24117 8938 24183 8941
rect 21357 8936 24183 8938
rect 21357 8880 21362 8936
rect 21418 8880 24122 8936
rect 24178 8880 24183 8936
rect 21357 8878 24183 8880
rect 21357 8875 21423 8878
rect 24117 8875 24183 8878
rect 3752 8736 4068 8737
rect 3752 8672 3758 8736
rect 3822 8672 3838 8736
rect 3902 8672 3918 8736
rect 3982 8672 3998 8736
rect 4062 8672 4068 8736
rect 3752 8671 4068 8672
rect 10468 8736 10784 8737
rect 10468 8672 10474 8736
rect 10538 8672 10554 8736
rect 10618 8672 10634 8736
rect 10698 8672 10714 8736
rect 10778 8672 10784 8736
rect 10468 8671 10784 8672
rect 17184 8736 17500 8737
rect 17184 8672 17190 8736
rect 17254 8672 17270 8736
rect 17334 8672 17350 8736
rect 17414 8672 17430 8736
rect 17494 8672 17500 8736
rect 17184 8671 17500 8672
rect 23900 8736 24216 8737
rect 23900 8672 23906 8736
rect 23970 8672 23986 8736
rect 24050 8672 24066 8736
rect 24130 8672 24146 8736
rect 24210 8672 24216 8736
rect 23900 8671 24216 8672
rect 11237 8530 11303 8533
rect 19425 8530 19491 8533
rect 11237 8528 19491 8530
rect 11237 8472 11242 8528
rect 11298 8472 19430 8528
rect 19486 8472 19491 8528
rect 11237 8470 19491 8472
rect 11237 8467 11303 8470
rect 19425 8467 19491 8470
rect 24669 8530 24735 8533
rect 24669 8528 24778 8530
rect 24669 8472 24674 8528
rect 24730 8472 24778 8528
rect 24669 8467 24778 8472
rect 8518 8332 8524 8396
rect 8588 8394 8594 8396
rect 9489 8394 9555 8397
rect 8588 8392 9555 8394
rect 8588 8336 9494 8392
rect 9550 8336 9555 8392
rect 8588 8334 9555 8336
rect 8588 8332 8594 8334
rect 9489 8331 9555 8334
rect 10317 8394 10383 8397
rect 15101 8394 15167 8397
rect 10317 8392 15167 8394
rect 10317 8336 10322 8392
rect 10378 8336 15106 8392
rect 15162 8336 15167 8392
rect 10317 8334 15167 8336
rect 10317 8331 10383 8334
rect 15101 8331 15167 8334
rect 24718 8261 24778 8467
rect 11605 8258 11671 8261
rect 13261 8258 13327 8261
rect 11605 8256 13327 8258
rect 11605 8200 11610 8256
rect 11666 8200 13266 8256
rect 13322 8200 13327 8256
rect 11605 8198 13327 8200
rect 11605 8195 11671 8198
rect 13261 8195 13327 8198
rect 24669 8256 24778 8261
rect 24669 8200 24674 8256
rect 24730 8200 24778 8256
rect 24669 8198 24778 8200
rect 24669 8195 24735 8198
rect 7110 8192 7426 8193
rect 7110 8128 7116 8192
rect 7180 8128 7196 8192
rect 7260 8128 7276 8192
rect 7340 8128 7356 8192
rect 7420 8128 7426 8192
rect 7110 8127 7426 8128
rect 13826 8192 14142 8193
rect 13826 8128 13832 8192
rect 13896 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14142 8192
rect 13826 8127 14142 8128
rect 20542 8192 20858 8193
rect 20542 8128 20548 8192
rect 20612 8128 20628 8192
rect 20692 8128 20708 8192
rect 20772 8128 20788 8192
rect 20852 8128 20858 8192
rect 20542 8127 20858 8128
rect 27258 8192 27574 8193
rect 27258 8128 27264 8192
rect 27328 8128 27344 8192
rect 27408 8128 27424 8192
rect 27488 8128 27504 8192
rect 27568 8128 27574 8192
rect 27258 8127 27574 8128
rect 24025 8122 24091 8125
rect 24393 8122 24459 8125
rect 24025 8120 24459 8122
rect 24025 8064 24030 8120
rect 24086 8064 24398 8120
rect 24454 8064 24459 8120
rect 24025 8062 24459 8064
rect 24025 8059 24091 8062
rect 24393 8059 24459 8062
rect 21633 7986 21699 7989
rect 24209 7986 24275 7989
rect 24577 7986 24643 7989
rect 25589 7986 25655 7989
rect 21633 7984 25655 7986
rect 21633 7928 21638 7984
rect 21694 7928 24214 7984
rect 24270 7928 24582 7984
rect 24638 7928 25594 7984
rect 25650 7928 25655 7984
rect 21633 7926 25655 7928
rect 21633 7923 21699 7926
rect 24209 7923 24275 7926
rect 24577 7923 24643 7926
rect 25589 7923 25655 7926
rect 20621 7714 20687 7717
rect 22277 7714 22343 7717
rect 22829 7714 22895 7717
rect 20621 7712 22895 7714
rect 20621 7656 20626 7712
rect 20682 7656 22282 7712
rect 22338 7656 22834 7712
rect 22890 7656 22895 7712
rect 20621 7654 22895 7656
rect 20621 7651 20687 7654
rect 22277 7651 22343 7654
rect 22829 7651 22895 7654
rect 3752 7648 4068 7649
rect 3752 7584 3758 7648
rect 3822 7584 3838 7648
rect 3902 7584 3918 7648
rect 3982 7584 3998 7648
rect 4062 7584 4068 7648
rect 3752 7583 4068 7584
rect 10468 7648 10784 7649
rect 10468 7584 10474 7648
rect 10538 7584 10554 7648
rect 10618 7584 10634 7648
rect 10698 7584 10714 7648
rect 10778 7584 10784 7648
rect 10468 7583 10784 7584
rect 17184 7648 17500 7649
rect 17184 7584 17190 7648
rect 17254 7584 17270 7648
rect 17334 7584 17350 7648
rect 17414 7584 17430 7648
rect 17494 7584 17500 7648
rect 17184 7583 17500 7584
rect 23900 7648 24216 7649
rect 23900 7584 23906 7648
rect 23970 7584 23986 7648
rect 24050 7584 24066 7648
rect 24130 7584 24146 7648
rect 24210 7584 24216 7648
rect 23900 7583 24216 7584
rect 7110 7104 7426 7105
rect 7110 7040 7116 7104
rect 7180 7040 7196 7104
rect 7260 7040 7276 7104
rect 7340 7040 7356 7104
rect 7420 7040 7426 7104
rect 7110 7039 7426 7040
rect 13826 7104 14142 7105
rect 13826 7040 13832 7104
rect 13896 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14142 7104
rect 13826 7039 14142 7040
rect 20542 7104 20858 7105
rect 20542 7040 20548 7104
rect 20612 7040 20628 7104
rect 20692 7040 20708 7104
rect 20772 7040 20788 7104
rect 20852 7040 20858 7104
rect 20542 7039 20858 7040
rect 27258 7104 27574 7105
rect 27258 7040 27264 7104
rect 27328 7040 27344 7104
rect 27408 7040 27424 7104
rect 27488 7040 27504 7104
rect 27568 7040 27574 7104
rect 27258 7039 27574 7040
rect 7833 6898 7899 6901
rect 10869 6900 10935 6901
rect 10869 6898 10916 6900
rect 7833 6896 10916 6898
rect 7833 6840 7838 6896
rect 7894 6840 10874 6896
rect 7833 6838 10916 6840
rect 7833 6835 7899 6838
rect 10869 6836 10916 6838
rect 10980 6836 10986 6900
rect 10869 6835 10935 6836
rect 7833 6762 7899 6765
rect 10409 6762 10475 6765
rect 7833 6760 10475 6762
rect 7833 6704 7838 6760
rect 7894 6704 10414 6760
rect 10470 6704 10475 6760
rect 7833 6702 10475 6704
rect 7833 6699 7899 6702
rect 10409 6699 10475 6702
rect 3752 6560 4068 6561
rect 3752 6496 3758 6560
rect 3822 6496 3838 6560
rect 3902 6496 3918 6560
rect 3982 6496 3998 6560
rect 4062 6496 4068 6560
rect 3752 6495 4068 6496
rect 10468 6560 10784 6561
rect 10468 6496 10474 6560
rect 10538 6496 10554 6560
rect 10618 6496 10634 6560
rect 10698 6496 10714 6560
rect 10778 6496 10784 6560
rect 10468 6495 10784 6496
rect 17184 6560 17500 6561
rect 17184 6496 17190 6560
rect 17254 6496 17270 6560
rect 17334 6496 17350 6560
rect 17414 6496 17430 6560
rect 17494 6496 17500 6560
rect 17184 6495 17500 6496
rect 23900 6560 24216 6561
rect 23900 6496 23906 6560
rect 23970 6496 23986 6560
rect 24050 6496 24066 6560
rect 24130 6496 24146 6560
rect 24210 6496 24216 6560
rect 23900 6495 24216 6496
rect 7110 6016 7426 6017
rect 7110 5952 7116 6016
rect 7180 5952 7196 6016
rect 7260 5952 7276 6016
rect 7340 5952 7356 6016
rect 7420 5952 7426 6016
rect 7110 5951 7426 5952
rect 13826 6016 14142 6017
rect 13826 5952 13832 6016
rect 13896 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14142 6016
rect 13826 5951 14142 5952
rect 20542 6016 20858 6017
rect 20542 5952 20548 6016
rect 20612 5952 20628 6016
rect 20692 5952 20708 6016
rect 20772 5952 20788 6016
rect 20852 5952 20858 6016
rect 20542 5951 20858 5952
rect 27258 6016 27574 6017
rect 27258 5952 27264 6016
rect 27328 5952 27344 6016
rect 27408 5952 27424 6016
rect 27488 5952 27504 6016
rect 27568 5952 27574 6016
rect 27258 5951 27574 5952
rect 12249 5946 12315 5949
rect 12566 5946 12572 5948
rect 12249 5944 12572 5946
rect 12249 5888 12254 5944
rect 12310 5888 12572 5944
rect 12249 5886 12572 5888
rect 12249 5883 12315 5886
rect 12566 5884 12572 5886
rect 12636 5884 12642 5948
rect 7925 5538 7991 5541
rect 8334 5538 8340 5540
rect 7925 5536 8340 5538
rect 7925 5480 7930 5536
rect 7986 5480 8340 5536
rect 7925 5478 8340 5480
rect 7925 5475 7991 5478
rect 8334 5476 8340 5478
rect 8404 5476 8410 5540
rect 3752 5472 4068 5473
rect 3752 5408 3758 5472
rect 3822 5408 3838 5472
rect 3902 5408 3918 5472
rect 3982 5408 3998 5472
rect 4062 5408 4068 5472
rect 3752 5407 4068 5408
rect 10468 5472 10784 5473
rect 10468 5408 10474 5472
rect 10538 5408 10554 5472
rect 10618 5408 10634 5472
rect 10698 5408 10714 5472
rect 10778 5408 10784 5472
rect 10468 5407 10784 5408
rect 17184 5472 17500 5473
rect 17184 5408 17190 5472
rect 17254 5408 17270 5472
rect 17334 5408 17350 5472
rect 17414 5408 17430 5472
rect 17494 5408 17500 5472
rect 17184 5407 17500 5408
rect 23900 5472 24216 5473
rect 23900 5408 23906 5472
rect 23970 5408 23986 5472
rect 24050 5408 24066 5472
rect 24130 5408 24146 5472
rect 24210 5408 24216 5472
rect 23900 5407 24216 5408
rect 13445 5266 13511 5269
rect 17125 5266 17191 5269
rect 13445 5264 17191 5266
rect 13445 5208 13450 5264
rect 13506 5208 17130 5264
rect 17186 5208 17191 5264
rect 13445 5206 17191 5208
rect 13445 5203 13511 5206
rect 17125 5203 17191 5206
rect 7110 4928 7426 4929
rect 7110 4864 7116 4928
rect 7180 4864 7196 4928
rect 7260 4864 7276 4928
rect 7340 4864 7356 4928
rect 7420 4864 7426 4928
rect 7110 4863 7426 4864
rect 13826 4928 14142 4929
rect 13826 4864 13832 4928
rect 13896 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14142 4928
rect 13826 4863 14142 4864
rect 20542 4928 20858 4929
rect 20542 4864 20548 4928
rect 20612 4864 20628 4928
rect 20692 4864 20708 4928
rect 20772 4864 20788 4928
rect 20852 4864 20858 4928
rect 20542 4863 20858 4864
rect 27258 4928 27574 4929
rect 27258 4864 27264 4928
rect 27328 4864 27344 4928
rect 27408 4864 27424 4928
rect 27488 4864 27504 4928
rect 27568 4864 27574 4928
rect 27258 4863 27574 4864
rect 16389 4722 16455 4725
rect 17033 4722 17099 4725
rect 16389 4720 17099 4722
rect 16389 4664 16394 4720
rect 16450 4664 17038 4720
rect 17094 4664 17099 4720
rect 16389 4662 17099 4664
rect 16389 4659 16455 4662
rect 17033 4659 17099 4662
rect 3752 4384 4068 4385
rect 3752 4320 3758 4384
rect 3822 4320 3838 4384
rect 3902 4320 3918 4384
rect 3982 4320 3998 4384
rect 4062 4320 4068 4384
rect 3752 4319 4068 4320
rect 10468 4384 10784 4385
rect 10468 4320 10474 4384
rect 10538 4320 10554 4384
rect 10618 4320 10634 4384
rect 10698 4320 10714 4384
rect 10778 4320 10784 4384
rect 10468 4319 10784 4320
rect 17184 4384 17500 4385
rect 17184 4320 17190 4384
rect 17254 4320 17270 4384
rect 17334 4320 17350 4384
rect 17414 4320 17430 4384
rect 17494 4320 17500 4384
rect 17184 4319 17500 4320
rect 23900 4384 24216 4385
rect 23900 4320 23906 4384
rect 23970 4320 23986 4384
rect 24050 4320 24066 4384
rect 24130 4320 24146 4384
rect 24210 4320 24216 4384
rect 23900 4319 24216 4320
rect 9857 4042 9923 4045
rect 11053 4042 11119 4045
rect 11789 4042 11855 4045
rect 9857 4040 11855 4042
rect 9857 3984 9862 4040
rect 9918 3984 11058 4040
rect 11114 3984 11794 4040
rect 11850 3984 11855 4040
rect 9857 3982 11855 3984
rect 9857 3979 9923 3982
rect 11053 3979 11119 3982
rect 11789 3979 11855 3982
rect 7110 3840 7426 3841
rect 7110 3776 7116 3840
rect 7180 3776 7196 3840
rect 7260 3776 7276 3840
rect 7340 3776 7356 3840
rect 7420 3776 7426 3840
rect 7110 3775 7426 3776
rect 13826 3840 14142 3841
rect 13826 3776 13832 3840
rect 13896 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14142 3840
rect 13826 3775 14142 3776
rect 20542 3840 20858 3841
rect 20542 3776 20548 3840
rect 20612 3776 20628 3840
rect 20692 3776 20708 3840
rect 20772 3776 20788 3840
rect 20852 3776 20858 3840
rect 20542 3775 20858 3776
rect 27258 3840 27574 3841
rect 27258 3776 27264 3840
rect 27328 3776 27344 3840
rect 27408 3776 27424 3840
rect 27488 3776 27504 3840
rect 27568 3776 27574 3840
rect 27258 3775 27574 3776
rect 5073 3634 5139 3637
rect 8753 3634 8819 3637
rect 14273 3634 14339 3637
rect 5073 3632 14339 3634
rect 5073 3576 5078 3632
rect 5134 3576 8758 3632
rect 8814 3576 14278 3632
rect 14334 3576 14339 3632
rect 5073 3574 14339 3576
rect 5073 3571 5139 3574
rect 8753 3571 8819 3574
rect 14273 3571 14339 3574
rect 13905 3498 13971 3501
rect 16941 3498 17007 3501
rect 13905 3496 17007 3498
rect 13905 3440 13910 3496
rect 13966 3440 16946 3496
rect 17002 3440 17007 3496
rect 13905 3438 17007 3440
rect 13905 3435 13971 3438
rect 16941 3435 17007 3438
rect 3752 3296 4068 3297
rect 3752 3232 3758 3296
rect 3822 3232 3838 3296
rect 3902 3232 3918 3296
rect 3982 3232 3998 3296
rect 4062 3232 4068 3296
rect 3752 3231 4068 3232
rect 10468 3296 10784 3297
rect 10468 3232 10474 3296
rect 10538 3232 10554 3296
rect 10618 3232 10634 3296
rect 10698 3232 10714 3296
rect 10778 3232 10784 3296
rect 10468 3231 10784 3232
rect 17184 3296 17500 3297
rect 17184 3232 17190 3296
rect 17254 3232 17270 3296
rect 17334 3232 17350 3296
rect 17414 3232 17430 3296
rect 17494 3232 17500 3296
rect 17184 3231 17500 3232
rect 23900 3296 24216 3297
rect 23900 3232 23906 3296
rect 23970 3232 23986 3296
rect 24050 3232 24066 3296
rect 24130 3232 24146 3296
rect 24210 3232 24216 3296
rect 23900 3231 24216 3232
rect 8845 3090 8911 3093
rect 9305 3090 9371 3093
rect 8845 3088 9371 3090
rect 8845 3032 8850 3088
rect 8906 3032 9310 3088
rect 9366 3032 9371 3088
rect 8845 3030 9371 3032
rect 8845 3027 8911 3030
rect 9305 3027 9371 3030
rect 9673 3090 9739 3093
rect 17953 3090 18019 3093
rect 9673 3088 18019 3090
rect 9673 3032 9678 3088
rect 9734 3032 17958 3088
rect 18014 3032 18019 3088
rect 9673 3030 18019 3032
rect 9673 3027 9739 3030
rect 17953 3027 18019 3030
rect 7557 2954 7623 2957
rect 8109 2954 8175 2957
rect 7557 2952 8175 2954
rect 7557 2896 7562 2952
rect 7618 2896 8114 2952
rect 8170 2896 8175 2952
rect 7557 2894 8175 2896
rect 7557 2891 7623 2894
rect 8109 2891 8175 2894
rect 7110 2752 7426 2753
rect 7110 2688 7116 2752
rect 7180 2688 7196 2752
rect 7260 2688 7276 2752
rect 7340 2688 7356 2752
rect 7420 2688 7426 2752
rect 7110 2687 7426 2688
rect 13826 2752 14142 2753
rect 13826 2688 13832 2752
rect 13896 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14142 2752
rect 13826 2687 14142 2688
rect 20542 2752 20858 2753
rect 20542 2688 20548 2752
rect 20612 2688 20628 2752
rect 20692 2688 20708 2752
rect 20772 2688 20788 2752
rect 20852 2688 20858 2752
rect 20542 2687 20858 2688
rect 27258 2752 27574 2753
rect 27258 2688 27264 2752
rect 27328 2688 27344 2752
rect 27408 2688 27424 2752
rect 27488 2688 27504 2752
rect 27568 2688 27574 2752
rect 27258 2687 27574 2688
rect 8385 2546 8451 2549
rect 8518 2546 8524 2548
rect 8385 2544 8524 2546
rect 8385 2488 8390 2544
rect 8446 2488 8524 2544
rect 8385 2486 8524 2488
rect 8385 2483 8451 2486
rect 8518 2484 8524 2486
rect 8588 2484 8594 2548
rect 11145 2546 11211 2549
rect 20345 2546 20411 2549
rect 20621 2546 20687 2549
rect 11145 2544 20687 2546
rect 11145 2488 11150 2544
rect 11206 2488 20350 2544
rect 20406 2488 20626 2544
rect 20682 2488 20687 2544
rect 11145 2486 20687 2488
rect 11145 2483 11211 2486
rect 20345 2483 20411 2486
rect 20621 2483 20687 2486
rect 3752 2208 4068 2209
rect 3752 2144 3758 2208
rect 3822 2144 3838 2208
rect 3902 2144 3918 2208
rect 3982 2144 3998 2208
rect 4062 2144 4068 2208
rect 3752 2143 4068 2144
rect 10468 2208 10784 2209
rect 10468 2144 10474 2208
rect 10538 2144 10554 2208
rect 10618 2144 10634 2208
rect 10698 2144 10714 2208
rect 10778 2144 10784 2208
rect 10468 2143 10784 2144
rect 17184 2208 17500 2209
rect 17184 2144 17190 2208
rect 17254 2144 17270 2208
rect 17334 2144 17350 2208
rect 17414 2144 17430 2208
rect 17494 2144 17500 2208
rect 17184 2143 17500 2144
rect 23900 2208 24216 2209
rect 23900 2144 23906 2208
rect 23970 2144 23986 2208
rect 24050 2144 24066 2208
rect 24130 2144 24146 2208
rect 24210 2144 24216 2208
rect 23900 2143 24216 2144
rect 10918 2078 17050 2138
rect 7557 2002 7623 2005
rect 10918 2002 10978 2078
rect 15929 2002 15995 2005
rect 16798 2002 16804 2004
rect 7557 2000 10978 2002
rect 7557 1944 7562 2000
rect 7618 1944 10978 2000
rect 7557 1942 10978 1944
rect 12390 2000 16804 2002
rect 12390 1944 15934 2000
rect 15990 1944 16804 2000
rect 12390 1942 16804 1944
rect 7557 1939 7623 1942
rect 7649 1866 7715 1869
rect 12390 1866 12450 1942
rect 15929 1939 15995 1942
rect 16798 1940 16804 1942
rect 16868 1940 16874 2004
rect 16990 2002 17050 2078
rect 17953 2002 18019 2005
rect 16990 2000 18019 2002
rect 16990 1944 17958 2000
rect 18014 1944 18019 2000
rect 16990 1942 18019 1944
rect 17953 1939 18019 1942
rect 7649 1864 12450 1866
rect 7649 1808 7654 1864
rect 7710 1808 12450 1864
rect 7649 1806 12450 1808
rect 7649 1803 7715 1806
rect 7110 1664 7426 1665
rect 7110 1600 7116 1664
rect 7180 1600 7196 1664
rect 7260 1600 7276 1664
rect 7340 1600 7356 1664
rect 7420 1600 7426 1664
rect 7110 1599 7426 1600
rect 13826 1664 14142 1665
rect 13826 1600 13832 1664
rect 13896 1600 13912 1664
rect 13976 1600 13992 1664
rect 14056 1600 14072 1664
rect 14136 1600 14142 1664
rect 13826 1599 14142 1600
rect 20542 1664 20858 1665
rect 20542 1600 20548 1664
rect 20612 1600 20628 1664
rect 20692 1600 20708 1664
rect 20772 1600 20788 1664
rect 20852 1600 20858 1664
rect 20542 1599 20858 1600
rect 27258 1664 27574 1665
rect 27258 1600 27264 1664
rect 27328 1600 27344 1664
rect 27408 1600 27424 1664
rect 27488 1600 27504 1664
rect 27568 1600 27574 1664
rect 27258 1599 27574 1600
rect 8518 1396 8524 1460
rect 8588 1458 8594 1460
rect 19241 1458 19307 1461
rect 8588 1456 19307 1458
rect 8588 1400 19246 1456
rect 19302 1400 19307 1456
rect 8588 1398 19307 1400
rect 8588 1396 8594 1398
rect 19241 1395 19307 1398
rect 3752 1120 4068 1121
rect 3752 1056 3758 1120
rect 3822 1056 3838 1120
rect 3902 1056 3918 1120
rect 3982 1056 3998 1120
rect 4062 1056 4068 1120
rect 3752 1055 4068 1056
rect 10468 1120 10784 1121
rect 10468 1056 10474 1120
rect 10538 1056 10554 1120
rect 10618 1056 10634 1120
rect 10698 1056 10714 1120
rect 10778 1056 10784 1120
rect 10468 1055 10784 1056
rect 17184 1120 17500 1121
rect 17184 1056 17190 1120
rect 17254 1056 17270 1120
rect 17334 1056 17350 1120
rect 17414 1056 17430 1120
rect 17494 1056 17500 1120
rect 17184 1055 17500 1056
rect 23900 1120 24216 1121
rect 23900 1056 23906 1120
rect 23970 1056 23986 1120
rect 24050 1056 24066 1120
rect 24130 1056 24146 1120
rect 24210 1056 24216 1120
rect 23900 1055 24216 1056
rect 7110 576 7426 577
rect 7110 512 7116 576
rect 7180 512 7196 576
rect 7260 512 7276 576
rect 7340 512 7356 576
rect 7420 512 7426 576
rect 7110 511 7426 512
rect 13826 576 14142 577
rect 13826 512 13832 576
rect 13896 512 13912 576
rect 13976 512 13992 576
rect 14056 512 14072 576
rect 14136 512 14142 576
rect 13826 511 14142 512
rect 20542 576 20858 577
rect 20542 512 20548 576
rect 20612 512 20628 576
rect 20692 512 20708 576
rect 20772 512 20788 576
rect 20852 512 20858 576
rect 20542 511 20858 512
rect 27258 576 27574 577
rect 27258 512 27264 576
rect 27328 512 27344 576
rect 27408 512 27424 576
rect 27488 512 27504 576
rect 27568 512 27574 576
rect 27258 511 27574 512
<< via3 >>
rect 3758 17436 3822 17440
rect 3758 17380 3762 17436
rect 3762 17380 3818 17436
rect 3818 17380 3822 17436
rect 3758 17376 3822 17380
rect 3838 17436 3902 17440
rect 3838 17380 3842 17436
rect 3842 17380 3898 17436
rect 3898 17380 3902 17436
rect 3838 17376 3902 17380
rect 3918 17436 3982 17440
rect 3918 17380 3922 17436
rect 3922 17380 3978 17436
rect 3978 17380 3982 17436
rect 3918 17376 3982 17380
rect 3998 17436 4062 17440
rect 3998 17380 4002 17436
rect 4002 17380 4058 17436
rect 4058 17380 4062 17436
rect 3998 17376 4062 17380
rect 10474 17436 10538 17440
rect 10474 17380 10478 17436
rect 10478 17380 10534 17436
rect 10534 17380 10538 17436
rect 10474 17376 10538 17380
rect 10554 17436 10618 17440
rect 10554 17380 10558 17436
rect 10558 17380 10614 17436
rect 10614 17380 10618 17436
rect 10554 17376 10618 17380
rect 10634 17436 10698 17440
rect 10634 17380 10638 17436
rect 10638 17380 10694 17436
rect 10694 17380 10698 17436
rect 10634 17376 10698 17380
rect 10714 17436 10778 17440
rect 10714 17380 10718 17436
rect 10718 17380 10774 17436
rect 10774 17380 10778 17436
rect 10714 17376 10778 17380
rect 17190 17436 17254 17440
rect 17190 17380 17194 17436
rect 17194 17380 17250 17436
rect 17250 17380 17254 17436
rect 17190 17376 17254 17380
rect 17270 17436 17334 17440
rect 17270 17380 17274 17436
rect 17274 17380 17330 17436
rect 17330 17380 17334 17436
rect 17270 17376 17334 17380
rect 17350 17436 17414 17440
rect 17350 17380 17354 17436
rect 17354 17380 17410 17436
rect 17410 17380 17414 17436
rect 17350 17376 17414 17380
rect 17430 17436 17494 17440
rect 17430 17380 17434 17436
rect 17434 17380 17490 17436
rect 17490 17380 17494 17436
rect 17430 17376 17494 17380
rect 23906 17436 23970 17440
rect 23906 17380 23910 17436
rect 23910 17380 23966 17436
rect 23966 17380 23970 17436
rect 23906 17376 23970 17380
rect 23986 17436 24050 17440
rect 23986 17380 23990 17436
rect 23990 17380 24046 17436
rect 24046 17380 24050 17436
rect 23986 17376 24050 17380
rect 24066 17436 24130 17440
rect 24066 17380 24070 17436
rect 24070 17380 24126 17436
rect 24126 17380 24130 17436
rect 24066 17376 24130 17380
rect 24146 17436 24210 17440
rect 24146 17380 24150 17436
rect 24150 17380 24206 17436
rect 24206 17380 24210 17436
rect 24146 17376 24210 17380
rect 7116 16892 7180 16896
rect 7116 16836 7120 16892
rect 7120 16836 7176 16892
rect 7176 16836 7180 16892
rect 7116 16832 7180 16836
rect 7196 16892 7260 16896
rect 7196 16836 7200 16892
rect 7200 16836 7256 16892
rect 7256 16836 7260 16892
rect 7196 16832 7260 16836
rect 7276 16892 7340 16896
rect 7276 16836 7280 16892
rect 7280 16836 7336 16892
rect 7336 16836 7340 16892
rect 7276 16832 7340 16836
rect 7356 16892 7420 16896
rect 7356 16836 7360 16892
rect 7360 16836 7416 16892
rect 7416 16836 7420 16892
rect 7356 16832 7420 16836
rect 13832 16892 13896 16896
rect 13832 16836 13836 16892
rect 13836 16836 13892 16892
rect 13892 16836 13896 16892
rect 13832 16832 13896 16836
rect 13912 16892 13976 16896
rect 13912 16836 13916 16892
rect 13916 16836 13972 16892
rect 13972 16836 13976 16892
rect 13912 16832 13976 16836
rect 13992 16892 14056 16896
rect 13992 16836 13996 16892
rect 13996 16836 14052 16892
rect 14052 16836 14056 16892
rect 13992 16832 14056 16836
rect 14072 16892 14136 16896
rect 14072 16836 14076 16892
rect 14076 16836 14132 16892
rect 14132 16836 14136 16892
rect 14072 16832 14136 16836
rect 20548 16892 20612 16896
rect 20548 16836 20552 16892
rect 20552 16836 20608 16892
rect 20608 16836 20612 16892
rect 20548 16832 20612 16836
rect 20628 16892 20692 16896
rect 20628 16836 20632 16892
rect 20632 16836 20688 16892
rect 20688 16836 20692 16892
rect 20628 16832 20692 16836
rect 20708 16892 20772 16896
rect 20708 16836 20712 16892
rect 20712 16836 20768 16892
rect 20768 16836 20772 16892
rect 20708 16832 20772 16836
rect 20788 16892 20852 16896
rect 20788 16836 20792 16892
rect 20792 16836 20848 16892
rect 20848 16836 20852 16892
rect 20788 16832 20852 16836
rect 27264 16892 27328 16896
rect 27264 16836 27268 16892
rect 27268 16836 27324 16892
rect 27324 16836 27328 16892
rect 27264 16832 27328 16836
rect 27344 16892 27408 16896
rect 27344 16836 27348 16892
rect 27348 16836 27404 16892
rect 27404 16836 27408 16892
rect 27344 16832 27408 16836
rect 27424 16892 27488 16896
rect 27424 16836 27428 16892
rect 27428 16836 27484 16892
rect 27484 16836 27488 16892
rect 27424 16832 27488 16836
rect 27504 16892 27568 16896
rect 27504 16836 27508 16892
rect 27508 16836 27564 16892
rect 27564 16836 27568 16892
rect 27504 16832 27568 16836
rect 12572 16628 12636 16692
rect 16804 16628 16868 16692
rect 3758 16348 3822 16352
rect 3758 16292 3762 16348
rect 3762 16292 3818 16348
rect 3818 16292 3822 16348
rect 3758 16288 3822 16292
rect 3838 16348 3902 16352
rect 3838 16292 3842 16348
rect 3842 16292 3898 16348
rect 3898 16292 3902 16348
rect 3838 16288 3902 16292
rect 3918 16348 3982 16352
rect 3918 16292 3922 16348
rect 3922 16292 3978 16348
rect 3978 16292 3982 16348
rect 3918 16288 3982 16292
rect 3998 16348 4062 16352
rect 3998 16292 4002 16348
rect 4002 16292 4058 16348
rect 4058 16292 4062 16348
rect 3998 16288 4062 16292
rect 10474 16348 10538 16352
rect 10474 16292 10478 16348
rect 10478 16292 10534 16348
rect 10534 16292 10538 16348
rect 10474 16288 10538 16292
rect 10554 16348 10618 16352
rect 10554 16292 10558 16348
rect 10558 16292 10614 16348
rect 10614 16292 10618 16348
rect 10554 16288 10618 16292
rect 10634 16348 10698 16352
rect 10634 16292 10638 16348
rect 10638 16292 10694 16348
rect 10694 16292 10698 16348
rect 10634 16288 10698 16292
rect 10714 16348 10778 16352
rect 10714 16292 10718 16348
rect 10718 16292 10774 16348
rect 10774 16292 10778 16348
rect 10714 16288 10778 16292
rect 17190 16348 17254 16352
rect 17190 16292 17194 16348
rect 17194 16292 17250 16348
rect 17250 16292 17254 16348
rect 17190 16288 17254 16292
rect 17270 16348 17334 16352
rect 17270 16292 17274 16348
rect 17274 16292 17330 16348
rect 17330 16292 17334 16348
rect 17270 16288 17334 16292
rect 17350 16348 17414 16352
rect 17350 16292 17354 16348
rect 17354 16292 17410 16348
rect 17410 16292 17414 16348
rect 17350 16288 17414 16292
rect 17430 16348 17494 16352
rect 17430 16292 17434 16348
rect 17434 16292 17490 16348
rect 17490 16292 17494 16348
rect 17430 16288 17494 16292
rect 23906 16348 23970 16352
rect 23906 16292 23910 16348
rect 23910 16292 23966 16348
rect 23966 16292 23970 16348
rect 23906 16288 23970 16292
rect 23986 16348 24050 16352
rect 23986 16292 23990 16348
rect 23990 16292 24046 16348
rect 24046 16292 24050 16348
rect 23986 16288 24050 16292
rect 24066 16348 24130 16352
rect 24066 16292 24070 16348
rect 24070 16292 24126 16348
rect 24126 16292 24130 16348
rect 24066 16288 24130 16292
rect 24146 16348 24210 16352
rect 24146 16292 24150 16348
rect 24150 16292 24206 16348
rect 24206 16292 24210 16348
rect 24146 16288 24210 16292
rect 7116 15804 7180 15808
rect 7116 15748 7120 15804
rect 7120 15748 7176 15804
rect 7176 15748 7180 15804
rect 7116 15744 7180 15748
rect 7196 15804 7260 15808
rect 7196 15748 7200 15804
rect 7200 15748 7256 15804
rect 7256 15748 7260 15804
rect 7196 15744 7260 15748
rect 7276 15804 7340 15808
rect 7276 15748 7280 15804
rect 7280 15748 7336 15804
rect 7336 15748 7340 15804
rect 7276 15744 7340 15748
rect 7356 15804 7420 15808
rect 7356 15748 7360 15804
rect 7360 15748 7416 15804
rect 7416 15748 7420 15804
rect 7356 15744 7420 15748
rect 13832 15804 13896 15808
rect 13832 15748 13836 15804
rect 13836 15748 13892 15804
rect 13892 15748 13896 15804
rect 13832 15744 13896 15748
rect 13912 15804 13976 15808
rect 13912 15748 13916 15804
rect 13916 15748 13972 15804
rect 13972 15748 13976 15804
rect 13912 15744 13976 15748
rect 13992 15804 14056 15808
rect 13992 15748 13996 15804
rect 13996 15748 14052 15804
rect 14052 15748 14056 15804
rect 13992 15744 14056 15748
rect 14072 15804 14136 15808
rect 14072 15748 14076 15804
rect 14076 15748 14132 15804
rect 14132 15748 14136 15804
rect 14072 15744 14136 15748
rect 20548 15804 20612 15808
rect 20548 15748 20552 15804
rect 20552 15748 20608 15804
rect 20608 15748 20612 15804
rect 20548 15744 20612 15748
rect 20628 15804 20692 15808
rect 20628 15748 20632 15804
rect 20632 15748 20688 15804
rect 20688 15748 20692 15804
rect 20628 15744 20692 15748
rect 20708 15804 20772 15808
rect 20708 15748 20712 15804
rect 20712 15748 20768 15804
rect 20768 15748 20772 15804
rect 20708 15744 20772 15748
rect 20788 15804 20852 15808
rect 20788 15748 20792 15804
rect 20792 15748 20848 15804
rect 20848 15748 20852 15804
rect 20788 15744 20852 15748
rect 27264 15804 27328 15808
rect 27264 15748 27268 15804
rect 27268 15748 27324 15804
rect 27324 15748 27328 15804
rect 27264 15744 27328 15748
rect 27344 15804 27408 15808
rect 27344 15748 27348 15804
rect 27348 15748 27404 15804
rect 27404 15748 27408 15804
rect 27344 15744 27408 15748
rect 27424 15804 27488 15808
rect 27424 15748 27428 15804
rect 27428 15748 27484 15804
rect 27484 15748 27488 15804
rect 27424 15744 27488 15748
rect 27504 15804 27568 15808
rect 27504 15748 27508 15804
rect 27508 15748 27564 15804
rect 27564 15748 27568 15804
rect 27504 15744 27568 15748
rect 3758 15260 3822 15264
rect 3758 15204 3762 15260
rect 3762 15204 3818 15260
rect 3818 15204 3822 15260
rect 3758 15200 3822 15204
rect 3838 15260 3902 15264
rect 3838 15204 3842 15260
rect 3842 15204 3898 15260
rect 3898 15204 3902 15260
rect 3838 15200 3902 15204
rect 3918 15260 3982 15264
rect 3918 15204 3922 15260
rect 3922 15204 3978 15260
rect 3978 15204 3982 15260
rect 3918 15200 3982 15204
rect 3998 15260 4062 15264
rect 3998 15204 4002 15260
rect 4002 15204 4058 15260
rect 4058 15204 4062 15260
rect 3998 15200 4062 15204
rect 10474 15260 10538 15264
rect 10474 15204 10478 15260
rect 10478 15204 10534 15260
rect 10534 15204 10538 15260
rect 10474 15200 10538 15204
rect 10554 15260 10618 15264
rect 10554 15204 10558 15260
rect 10558 15204 10614 15260
rect 10614 15204 10618 15260
rect 10554 15200 10618 15204
rect 10634 15260 10698 15264
rect 10634 15204 10638 15260
rect 10638 15204 10694 15260
rect 10694 15204 10698 15260
rect 10634 15200 10698 15204
rect 10714 15260 10778 15264
rect 10714 15204 10718 15260
rect 10718 15204 10774 15260
rect 10774 15204 10778 15260
rect 10714 15200 10778 15204
rect 17190 15260 17254 15264
rect 17190 15204 17194 15260
rect 17194 15204 17250 15260
rect 17250 15204 17254 15260
rect 17190 15200 17254 15204
rect 17270 15260 17334 15264
rect 17270 15204 17274 15260
rect 17274 15204 17330 15260
rect 17330 15204 17334 15260
rect 17270 15200 17334 15204
rect 17350 15260 17414 15264
rect 17350 15204 17354 15260
rect 17354 15204 17410 15260
rect 17410 15204 17414 15260
rect 17350 15200 17414 15204
rect 17430 15260 17494 15264
rect 17430 15204 17434 15260
rect 17434 15204 17490 15260
rect 17490 15204 17494 15260
rect 17430 15200 17494 15204
rect 23906 15260 23970 15264
rect 23906 15204 23910 15260
rect 23910 15204 23966 15260
rect 23966 15204 23970 15260
rect 23906 15200 23970 15204
rect 23986 15260 24050 15264
rect 23986 15204 23990 15260
rect 23990 15204 24046 15260
rect 24046 15204 24050 15260
rect 23986 15200 24050 15204
rect 24066 15260 24130 15264
rect 24066 15204 24070 15260
rect 24070 15204 24126 15260
rect 24126 15204 24130 15260
rect 24066 15200 24130 15204
rect 24146 15260 24210 15264
rect 24146 15204 24150 15260
rect 24150 15204 24206 15260
rect 24206 15204 24210 15260
rect 24146 15200 24210 15204
rect 7116 14716 7180 14720
rect 7116 14660 7120 14716
rect 7120 14660 7176 14716
rect 7176 14660 7180 14716
rect 7116 14656 7180 14660
rect 7196 14716 7260 14720
rect 7196 14660 7200 14716
rect 7200 14660 7256 14716
rect 7256 14660 7260 14716
rect 7196 14656 7260 14660
rect 7276 14716 7340 14720
rect 7276 14660 7280 14716
rect 7280 14660 7336 14716
rect 7336 14660 7340 14716
rect 7276 14656 7340 14660
rect 7356 14716 7420 14720
rect 7356 14660 7360 14716
rect 7360 14660 7416 14716
rect 7416 14660 7420 14716
rect 7356 14656 7420 14660
rect 13832 14716 13896 14720
rect 13832 14660 13836 14716
rect 13836 14660 13892 14716
rect 13892 14660 13896 14716
rect 13832 14656 13896 14660
rect 13912 14716 13976 14720
rect 13912 14660 13916 14716
rect 13916 14660 13972 14716
rect 13972 14660 13976 14716
rect 13912 14656 13976 14660
rect 13992 14716 14056 14720
rect 13992 14660 13996 14716
rect 13996 14660 14052 14716
rect 14052 14660 14056 14716
rect 13992 14656 14056 14660
rect 14072 14716 14136 14720
rect 14072 14660 14076 14716
rect 14076 14660 14132 14716
rect 14132 14660 14136 14716
rect 14072 14656 14136 14660
rect 20548 14716 20612 14720
rect 20548 14660 20552 14716
rect 20552 14660 20608 14716
rect 20608 14660 20612 14716
rect 20548 14656 20612 14660
rect 20628 14716 20692 14720
rect 20628 14660 20632 14716
rect 20632 14660 20688 14716
rect 20688 14660 20692 14716
rect 20628 14656 20692 14660
rect 20708 14716 20772 14720
rect 20708 14660 20712 14716
rect 20712 14660 20768 14716
rect 20768 14660 20772 14716
rect 20708 14656 20772 14660
rect 20788 14716 20852 14720
rect 20788 14660 20792 14716
rect 20792 14660 20848 14716
rect 20848 14660 20852 14716
rect 20788 14656 20852 14660
rect 27264 14716 27328 14720
rect 27264 14660 27268 14716
rect 27268 14660 27324 14716
rect 27324 14660 27328 14716
rect 27264 14656 27328 14660
rect 27344 14716 27408 14720
rect 27344 14660 27348 14716
rect 27348 14660 27404 14716
rect 27404 14660 27408 14716
rect 27344 14656 27408 14660
rect 27424 14716 27488 14720
rect 27424 14660 27428 14716
rect 27428 14660 27484 14716
rect 27484 14660 27488 14716
rect 27424 14656 27488 14660
rect 27504 14716 27568 14720
rect 27504 14660 27508 14716
rect 27508 14660 27564 14716
rect 27564 14660 27568 14716
rect 27504 14656 27568 14660
rect 3758 14172 3822 14176
rect 3758 14116 3762 14172
rect 3762 14116 3818 14172
rect 3818 14116 3822 14172
rect 3758 14112 3822 14116
rect 3838 14172 3902 14176
rect 3838 14116 3842 14172
rect 3842 14116 3898 14172
rect 3898 14116 3902 14172
rect 3838 14112 3902 14116
rect 3918 14172 3982 14176
rect 3918 14116 3922 14172
rect 3922 14116 3978 14172
rect 3978 14116 3982 14172
rect 3918 14112 3982 14116
rect 3998 14172 4062 14176
rect 3998 14116 4002 14172
rect 4002 14116 4058 14172
rect 4058 14116 4062 14172
rect 3998 14112 4062 14116
rect 10474 14172 10538 14176
rect 10474 14116 10478 14172
rect 10478 14116 10534 14172
rect 10534 14116 10538 14172
rect 10474 14112 10538 14116
rect 10554 14172 10618 14176
rect 10554 14116 10558 14172
rect 10558 14116 10614 14172
rect 10614 14116 10618 14172
rect 10554 14112 10618 14116
rect 10634 14172 10698 14176
rect 10634 14116 10638 14172
rect 10638 14116 10694 14172
rect 10694 14116 10698 14172
rect 10634 14112 10698 14116
rect 10714 14172 10778 14176
rect 10714 14116 10718 14172
rect 10718 14116 10774 14172
rect 10774 14116 10778 14172
rect 10714 14112 10778 14116
rect 17190 14172 17254 14176
rect 17190 14116 17194 14172
rect 17194 14116 17250 14172
rect 17250 14116 17254 14172
rect 17190 14112 17254 14116
rect 17270 14172 17334 14176
rect 17270 14116 17274 14172
rect 17274 14116 17330 14172
rect 17330 14116 17334 14172
rect 17270 14112 17334 14116
rect 17350 14172 17414 14176
rect 17350 14116 17354 14172
rect 17354 14116 17410 14172
rect 17410 14116 17414 14172
rect 17350 14112 17414 14116
rect 17430 14172 17494 14176
rect 17430 14116 17434 14172
rect 17434 14116 17490 14172
rect 17490 14116 17494 14172
rect 17430 14112 17494 14116
rect 23906 14172 23970 14176
rect 23906 14116 23910 14172
rect 23910 14116 23966 14172
rect 23966 14116 23970 14172
rect 23906 14112 23970 14116
rect 23986 14172 24050 14176
rect 23986 14116 23990 14172
rect 23990 14116 24046 14172
rect 24046 14116 24050 14172
rect 23986 14112 24050 14116
rect 24066 14172 24130 14176
rect 24066 14116 24070 14172
rect 24070 14116 24126 14172
rect 24126 14116 24130 14172
rect 24066 14112 24130 14116
rect 24146 14172 24210 14176
rect 24146 14116 24150 14172
rect 24150 14116 24206 14172
rect 24206 14116 24210 14172
rect 24146 14112 24210 14116
rect 7116 13628 7180 13632
rect 7116 13572 7120 13628
rect 7120 13572 7176 13628
rect 7176 13572 7180 13628
rect 7116 13568 7180 13572
rect 7196 13628 7260 13632
rect 7196 13572 7200 13628
rect 7200 13572 7256 13628
rect 7256 13572 7260 13628
rect 7196 13568 7260 13572
rect 7276 13628 7340 13632
rect 7276 13572 7280 13628
rect 7280 13572 7336 13628
rect 7336 13572 7340 13628
rect 7276 13568 7340 13572
rect 7356 13628 7420 13632
rect 7356 13572 7360 13628
rect 7360 13572 7416 13628
rect 7416 13572 7420 13628
rect 7356 13568 7420 13572
rect 13832 13628 13896 13632
rect 13832 13572 13836 13628
rect 13836 13572 13892 13628
rect 13892 13572 13896 13628
rect 13832 13568 13896 13572
rect 13912 13628 13976 13632
rect 13912 13572 13916 13628
rect 13916 13572 13972 13628
rect 13972 13572 13976 13628
rect 13912 13568 13976 13572
rect 13992 13628 14056 13632
rect 13992 13572 13996 13628
rect 13996 13572 14052 13628
rect 14052 13572 14056 13628
rect 13992 13568 14056 13572
rect 14072 13628 14136 13632
rect 14072 13572 14076 13628
rect 14076 13572 14132 13628
rect 14132 13572 14136 13628
rect 14072 13568 14136 13572
rect 20548 13628 20612 13632
rect 20548 13572 20552 13628
rect 20552 13572 20608 13628
rect 20608 13572 20612 13628
rect 20548 13568 20612 13572
rect 20628 13628 20692 13632
rect 20628 13572 20632 13628
rect 20632 13572 20688 13628
rect 20688 13572 20692 13628
rect 20628 13568 20692 13572
rect 20708 13628 20772 13632
rect 20708 13572 20712 13628
rect 20712 13572 20768 13628
rect 20768 13572 20772 13628
rect 20708 13568 20772 13572
rect 20788 13628 20852 13632
rect 20788 13572 20792 13628
rect 20792 13572 20848 13628
rect 20848 13572 20852 13628
rect 20788 13568 20852 13572
rect 27264 13628 27328 13632
rect 27264 13572 27268 13628
rect 27268 13572 27324 13628
rect 27324 13572 27328 13628
rect 27264 13568 27328 13572
rect 27344 13628 27408 13632
rect 27344 13572 27348 13628
rect 27348 13572 27404 13628
rect 27404 13572 27408 13628
rect 27344 13568 27408 13572
rect 27424 13628 27488 13632
rect 27424 13572 27428 13628
rect 27428 13572 27484 13628
rect 27484 13572 27488 13628
rect 27424 13568 27488 13572
rect 27504 13628 27568 13632
rect 27504 13572 27508 13628
rect 27508 13572 27564 13628
rect 27564 13572 27568 13628
rect 27504 13568 27568 13572
rect 3758 13084 3822 13088
rect 3758 13028 3762 13084
rect 3762 13028 3818 13084
rect 3818 13028 3822 13084
rect 3758 13024 3822 13028
rect 3838 13084 3902 13088
rect 3838 13028 3842 13084
rect 3842 13028 3898 13084
rect 3898 13028 3902 13084
rect 3838 13024 3902 13028
rect 3918 13084 3982 13088
rect 3918 13028 3922 13084
rect 3922 13028 3978 13084
rect 3978 13028 3982 13084
rect 3918 13024 3982 13028
rect 3998 13084 4062 13088
rect 3998 13028 4002 13084
rect 4002 13028 4058 13084
rect 4058 13028 4062 13084
rect 3998 13024 4062 13028
rect 10474 13084 10538 13088
rect 10474 13028 10478 13084
rect 10478 13028 10534 13084
rect 10534 13028 10538 13084
rect 10474 13024 10538 13028
rect 10554 13084 10618 13088
rect 10554 13028 10558 13084
rect 10558 13028 10614 13084
rect 10614 13028 10618 13084
rect 10554 13024 10618 13028
rect 10634 13084 10698 13088
rect 10634 13028 10638 13084
rect 10638 13028 10694 13084
rect 10694 13028 10698 13084
rect 10634 13024 10698 13028
rect 10714 13084 10778 13088
rect 10714 13028 10718 13084
rect 10718 13028 10774 13084
rect 10774 13028 10778 13084
rect 10714 13024 10778 13028
rect 17190 13084 17254 13088
rect 17190 13028 17194 13084
rect 17194 13028 17250 13084
rect 17250 13028 17254 13084
rect 17190 13024 17254 13028
rect 17270 13084 17334 13088
rect 17270 13028 17274 13084
rect 17274 13028 17330 13084
rect 17330 13028 17334 13084
rect 17270 13024 17334 13028
rect 17350 13084 17414 13088
rect 17350 13028 17354 13084
rect 17354 13028 17410 13084
rect 17410 13028 17414 13084
rect 17350 13024 17414 13028
rect 17430 13084 17494 13088
rect 17430 13028 17434 13084
rect 17434 13028 17490 13084
rect 17490 13028 17494 13084
rect 17430 13024 17494 13028
rect 23906 13084 23970 13088
rect 23906 13028 23910 13084
rect 23910 13028 23966 13084
rect 23966 13028 23970 13084
rect 23906 13024 23970 13028
rect 23986 13084 24050 13088
rect 23986 13028 23990 13084
rect 23990 13028 24046 13084
rect 24046 13028 24050 13084
rect 23986 13024 24050 13028
rect 24066 13084 24130 13088
rect 24066 13028 24070 13084
rect 24070 13028 24126 13084
rect 24126 13028 24130 13084
rect 24066 13024 24130 13028
rect 24146 13084 24210 13088
rect 24146 13028 24150 13084
rect 24150 13028 24206 13084
rect 24206 13028 24210 13084
rect 24146 13024 24210 13028
rect 7116 12540 7180 12544
rect 7116 12484 7120 12540
rect 7120 12484 7176 12540
rect 7176 12484 7180 12540
rect 7116 12480 7180 12484
rect 7196 12540 7260 12544
rect 7196 12484 7200 12540
rect 7200 12484 7256 12540
rect 7256 12484 7260 12540
rect 7196 12480 7260 12484
rect 7276 12540 7340 12544
rect 7276 12484 7280 12540
rect 7280 12484 7336 12540
rect 7336 12484 7340 12540
rect 7276 12480 7340 12484
rect 7356 12540 7420 12544
rect 7356 12484 7360 12540
rect 7360 12484 7416 12540
rect 7416 12484 7420 12540
rect 7356 12480 7420 12484
rect 13832 12540 13896 12544
rect 13832 12484 13836 12540
rect 13836 12484 13892 12540
rect 13892 12484 13896 12540
rect 13832 12480 13896 12484
rect 13912 12540 13976 12544
rect 13912 12484 13916 12540
rect 13916 12484 13972 12540
rect 13972 12484 13976 12540
rect 13912 12480 13976 12484
rect 13992 12540 14056 12544
rect 13992 12484 13996 12540
rect 13996 12484 14052 12540
rect 14052 12484 14056 12540
rect 13992 12480 14056 12484
rect 14072 12540 14136 12544
rect 14072 12484 14076 12540
rect 14076 12484 14132 12540
rect 14132 12484 14136 12540
rect 14072 12480 14136 12484
rect 20548 12540 20612 12544
rect 20548 12484 20552 12540
rect 20552 12484 20608 12540
rect 20608 12484 20612 12540
rect 20548 12480 20612 12484
rect 20628 12540 20692 12544
rect 20628 12484 20632 12540
rect 20632 12484 20688 12540
rect 20688 12484 20692 12540
rect 20628 12480 20692 12484
rect 20708 12540 20772 12544
rect 20708 12484 20712 12540
rect 20712 12484 20768 12540
rect 20768 12484 20772 12540
rect 20708 12480 20772 12484
rect 20788 12540 20852 12544
rect 20788 12484 20792 12540
rect 20792 12484 20848 12540
rect 20848 12484 20852 12540
rect 20788 12480 20852 12484
rect 27264 12540 27328 12544
rect 27264 12484 27268 12540
rect 27268 12484 27324 12540
rect 27324 12484 27328 12540
rect 27264 12480 27328 12484
rect 27344 12540 27408 12544
rect 27344 12484 27348 12540
rect 27348 12484 27404 12540
rect 27404 12484 27408 12540
rect 27344 12480 27408 12484
rect 27424 12540 27488 12544
rect 27424 12484 27428 12540
rect 27428 12484 27484 12540
rect 27484 12484 27488 12540
rect 27424 12480 27488 12484
rect 27504 12540 27568 12544
rect 27504 12484 27508 12540
rect 27508 12484 27564 12540
rect 27564 12484 27568 12540
rect 27504 12480 27568 12484
rect 10916 12336 10980 12340
rect 10916 12280 10966 12336
rect 10966 12280 10980 12336
rect 10916 12276 10980 12280
rect 26188 12336 26252 12340
rect 26188 12280 26202 12336
rect 26202 12280 26252 12336
rect 26188 12276 26252 12280
rect 3758 11996 3822 12000
rect 3758 11940 3762 11996
rect 3762 11940 3818 11996
rect 3818 11940 3822 11996
rect 3758 11936 3822 11940
rect 3838 11996 3902 12000
rect 3838 11940 3842 11996
rect 3842 11940 3898 11996
rect 3898 11940 3902 11996
rect 3838 11936 3902 11940
rect 3918 11996 3982 12000
rect 3918 11940 3922 11996
rect 3922 11940 3978 11996
rect 3978 11940 3982 11996
rect 3918 11936 3982 11940
rect 3998 11996 4062 12000
rect 3998 11940 4002 11996
rect 4002 11940 4058 11996
rect 4058 11940 4062 11996
rect 3998 11936 4062 11940
rect 10474 11996 10538 12000
rect 10474 11940 10478 11996
rect 10478 11940 10534 11996
rect 10534 11940 10538 11996
rect 10474 11936 10538 11940
rect 10554 11996 10618 12000
rect 10554 11940 10558 11996
rect 10558 11940 10614 11996
rect 10614 11940 10618 11996
rect 10554 11936 10618 11940
rect 10634 11996 10698 12000
rect 10634 11940 10638 11996
rect 10638 11940 10694 11996
rect 10694 11940 10698 11996
rect 10634 11936 10698 11940
rect 10714 11996 10778 12000
rect 10714 11940 10718 11996
rect 10718 11940 10774 11996
rect 10774 11940 10778 11996
rect 10714 11936 10778 11940
rect 17190 11996 17254 12000
rect 17190 11940 17194 11996
rect 17194 11940 17250 11996
rect 17250 11940 17254 11996
rect 17190 11936 17254 11940
rect 17270 11996 17334 12000
rect 17270 11940 17274 11996
rect 17274 11940 17330 11996
rect 17330 11940 17334 11996
rect 17270 11936 17334 11940
rect 17350 11996 17414 12000
rect 17350 11940 17354 11996
rect 17354 11940 17410 11996
rect 17410 11940 17414 11996
rect 17350 11936 17414 11940
rect 17430 11996 17494 12000
rect 17430 11940 17434 11996
rect 17434 11940 17490 11996
rect 17490 11940 17494 11996
rect 17430 11936 17494 11940
rect 23906 11996 23970 12000
rect 23906 11940 23910 11996
rect 23910 11940 23966 11996
rect 23966 11940 23970 11996
rect 23906 11936 23970 11940
rect 23986 11996 24050 12000
rect 23986 11940 23990 11996
rect 23990 11940 24046 11996
rect 24046 11940 24050 11996
rect 23986 11936 24050 11940
rect 24066 11996 24130 12000
rect 24066 11940 24070 11996
rect 24070 11940 24126 11996
rect 24126 11940 24130 11996
rect 24066 11936 24130 11940
rect 24146 11996 24210 12000
rect 24146 11940 24150 11996
rect 24150 11940 24206 11996
rect 24206 11940 24210 11996
rect 24146 11936 24210 11940
rect 7116 11452 7180 11456
rect 7116 11396 7120 11452
rect 7120 11396 7176 11452
rect 7176 11396 7180 11452
rect 7116 11392 7180 11396
rect 7196 11452 7260 11456
rect 7196 11396 7200 11452
rect 7200 11396 7256 11452
rect 7256 11396 7260 11452
rect 7196 11392 7260 11396
rect 7276 11452 7340 11456
rect 7276 11396 7280 11452
rect 7280 11396 7336 11452
rect 7336 11396 7340 11452
rect 7276 11392 7340 11396
rect 7356 11452 7420 11456
rect 7356 11396 7360 11452
rect 7360 11396 7416 11452
rect 7416 11396 7420 11452
rect 7356 11392 7420 11396
rect 13832 11452 13896 11456
rect 13832 11396 13836 11452
rect 13836 11396 13892 11452
rect 13892 11396 13896 11452
rect 13832 11392 13896 11396
rect 13912 11452 13976 11456
rect 13912 11396 13916 11452
rect 13916 11396 13972 11452
rect 13972 11396 13976 11452
rect 13912 11392 13976 11396
rect 13992 11452 14056 11456
rect 13992 11396 13996 11452
rect 13996 11396 14052 11452
rect 14052 11396 14056 11452
rect 13992 11392 14056 11396
rect 14072 11452 14136 11456
rect 14072 11396 14076 11452
rect 14076 11396 14132 11452
rect 14132 11396 14136 11452
rect 14072 11392 14136 11396
rect 20548 11452 20612 11456
rect 20548 11396 20552 11452
rect 20552 11396 20608 11452
rect 20608 11396 20612 11452
rect 20548 11392 20612 11396
rect 20628 11452 20692 11456
rect 20628 11396 20632 11452
rect 20632 11396 20688 11452
rect 20688 11396 20692 11452
rect 20628 11392 20692 11396
rect 20708 11452 20772 11456
rect 20708 11396 20712 11452
rect 20712 11396 20768 11452
rect 20768 11396 20772 11452
rect 20708 11392 20772 11396
rect 20788 11452 20852 11456
rect 20788 11396 20792 11452
rect 20792 11396 20848 11452
rect 20848 11396 20852 11452
rect 20788 11392 20852 11396
rect 27264 11452 27328 11456
rect 27264 11396 27268 11452
rect 27268 11396 27324 11452
rect 27324 11396 27328 11452
rect 27264 11392 27328 11396
rect 27344 11452 27408 11456
rect 27344 11396 27348 11452
rect 27348 11396 27404 11452
rect 27404 11396 27408 11452
rect 27344 11392 27408 11396
rect 27424 11452 27488 11456
rect 27424 11396 27428 11452
rect 27428 11396 27484 11452
rect 27484 11396 27488 11452
rect 27424 11392 27488 11396
rect 27504 11452 27568 11456
rect 27504 11396 27508 11452
rect 27508 11396 27564 11452
rect 27564 11396 27568 11452
rect 27504 11392 27568 11396
rect 3758 10908 3822 10912
rect 3758 10852 3762 10908
rect 3762 10852 3818 10908
rect 3818 10852 3822 10908
rect 3758 10848 3822 10852
rect 3838 10908 3902 10912
rect 3838 10852 3842 10908
rect 3842 10852 3898 10908
rect 3898 10852 3902 10908
rect 3838 10848 3902 10852
rect 3918 10908 3982 10912
rect 3918 10852 3922 10908
rect 3922 10852 3978 10908
rect 3978 10852 3982 10908
rect 3918 10848 3982 10852
rect 3998 10908 4062 10912
rect 3998 10852 4002 10908
rect 4002 10852 4058 10908
rect 4058 10852 4062 10908
rect 3998 10848 4062 10852
rect 10474 10908 10538 10912
rect 10474 10852 10478 10908
rect 10478 10852 10534 10908
rect 10534 10852 10538 10908
rect 10474 10848 10538 10852
rect 10554 10908 10618 10912
rect 10554 10852 10558 10908
rect 10558 10852 10614 10908
rect 10614 10852 10618 10908
rect 10554 10848 10618 10852
rect 10634 10908 10698 10912
rect 10634 10852 10638 10908
rect 10638 10852 10694 10908
rect 10694 10852 10698 10908
rect 10634 10848 10698 10852
rect 10714 10908 10778 10912
rect 10714 10852 10718 10908
rect 10718 10852 10774 10908
rect 10774 10852 10778 10908
rect 10714 10848 10778 10852
rect 17190 10908 17254 10912
rect 17190 10852 17194 10908
rect 17194 10852 17250 10908
rect 17250 10852 17254 10908
rect 17190 10848 17254 10852
rect 17270 10908 17334 10912
rect 17270 10852 17274 10908
rect 17274 10852 17330 10908
rect 17330 10852 17334 10908
rect 17270 10848 17334 10852
rect 17350 10908 17414 10912
rect 17350 10852 17354 10908
rect 17354 10852 17410 10908
rect 17410 10852 17414 10908
rect 17350 10848 17414 10852
rect 17430 10908 17494 10912
rect 17430 10852 17434 10908
rect 17434 10852 17490 10908
rect 17490 10852 17494 10908
rect 17430 10848 17494 10852
rect 23906 10908 23970 10912
rect 23906 10852 23910 10908
rect 23910 10852 23966 10908
rect 23966 10852 23970 10908
rect 23906 10848 23970 10852
rect 23986 10908 24050 10912
rect 23986 10852 23990 10908
rect 23990 10852 24046 10908
rect 24046 10852 24050 10908
rect 23986 10848 24050 10852
rect 24066 10908 24130 10912
rect 24066 10852 24070 10908
rect 24070 10852 24126 10908
rect 24126 10852 24130 10908
rect 24066 10848 24130 10852
rect 24146 10908 24210 10912
rect 24146 10852 24150 10908
rect 24150 10852 24206 10908
rect 24206 10852 24210 10908
rect 24146 10848 24210 10852
rect 7116 10364 7180 10368
rect 7116 10308 7120 10364
rect 7120 10308 7176 10364
rect 7176 10308 7180 10364
rect 7116 10304 7180 10308
rect 7196 10364 7260 10368
rect 7196 10308 7200 10364
rect 7200 10308 7256 10364
rect 7256 10308 7260 10364
rect 7196 10304 7260 10308
rect 7276 10364 7340 10368
rect 7276 10308 7280 10364
rect 7280 10308 7336 10364
rect 7336 10308 7340 10364
rect 7276 10304 7340 10308
rect 7356 10364 7420 10368
rect 7356 10308 7360 10364
rect 7360 10308 7416 10364
rect 7416 10308 7420 10364
rect 7356 10304 7420 10308
rect 13832 10364 13896 10368
rect 13832 10308 13836 10364
rect 13836 10308 13892 10364
rect 13892 10308 13896 10364
rect 13832 10304 13896 10308
rect 13912 10364 13976 10368
rect 13912 10308 13916 10364
rect 13916 10308 13972 10364
rect 13972 10308 13976 10364
rect 13912 10304 13976 10308
rect 13992 10364 14056 10368
rect 13992 10308 13996 10364
rect 13996 10308 14052 10364
rect 14052 10308 14056 10364
rect 13992 10304 14056 10308
rect 14072 10364 14136 10368
rect 14072 10308 14076 10364
rect 14076 10308 14132 10364
rect 14132 10308 14136 10364
rect 14072 10304 14136 10308
rect 20548 10364 20612 10368
rect 20548 10308 20552 10364
rect 20552 10308 20608 10364
rect 20608 10308 20612 10364
rect 20548 10304 20612 10308
rect 20628 10364 20692 10368
rect 20628 10308 20632 10364
rect 20632 10308 20688 10364
rect 20688 10308 20692 10364
rect 20628 10304 20692 10308
rect 20708 10364 20772 10368
rect 20708 10308 20712 10364
rect 20712 10308 20768 10364
rect 20768 10308 20772 10364
rect 20708 10304 20772 10308
rect 20788 10364 20852 10368
rect 20788 10308 20792 10364
rect 20792 10308 20848 10364
rect 20848 10308 20852 10364
rect 20788 10304 20852 10308
rect 27264 10364 27328 10368
rect 27264 10308 27268 10364
rect 27268 10308 27324 10364
rect 27324 10308 27328 10364
rect 27264 10304 27328 10308
rect 27344 10364 27408 10368
rect 27344 10308 27348 10364
rect 27348 10308 27404 10364
rect 27404 10308 27408 10364
rect 27344 10304 27408 10308
rect 27424 10364 27488 10368
rect 27424 10308 27428 10364
rect 27428 10308 27484 10364
rect 27484 10308 27488 10364
rect 27424 10304 27488 10308
rect 27504 10364 27568 10368
rect 27504 10308 27508 10364
rect 27508 10308 27564 10364
rect 27564 10308 27568 10364
rect 27504 10304 27568 10308
rect 3758 9820 3822 9824
rect 3758 9764 3762 9820
rect 3762 9764 3818 9820
rect 3818 9764 3822 9820
rect 3758 9760 3822 9764
rect 3838 9820 3902 9824
rect 3838 9764 3842 9820
rect 3842 9764 3898 9820
rect 3898 9764 3902 9820
rect 3838 9760 3902 9764
rect 3918 9820 3982 9824
rect 3918 9764 3922 9820
rect 3922 9764 3978 9820
rect 3978 9764 3982 9820
rect 3918 9760 3982 9764
rect 3998 9820 4062 9824
rect 3998 9764 4002 9820
rect 4002 9764 4058 9820
rect 4058 9764 4062 9820
rect 3998 9760 4062 9764
rect 10474 9820 10538 9824
rect 10474 9764 10478 9820
rect 10478 9764 10534 9820
rect 10534 9764 10538 9820
rect 10474 9760 10538 9764
rect 10554 9820 10618 9824
rect 10554 9764 10558 9820
rect 10558 9764 10614 9820
rect 10614 9764 10618 9820
rect 10554 9760 10618 9764
rect 10634 9820 10698 9824
rect 10634 9764 10638 9820
rect 10638 9764 10694 9820
rect 10694 9764 10698 9820
rect 10634 9760 10698 9764
rect 10714 9820 10778 9824
rect 10714 9764 10718 9820
rect 10718 9764 10774 9820
rect 10774 9764 10778 9820
rect 10714 9760 10778 9764
rect 17190 9820 17254 9824
rect 17190 9764 17194 9820
rect 17194 9764 17250 9820
rect 17250 9764 17254 9820
rect 17190 9760 17254 9764
rect 17270 9820 17334 9824
rect 17270 9764 17274 9820
rect 17274 9764 17330 9820
rect 17330 9764 17334 9820
rect 17270 9760 17334 9764
rect 17350 9820 17414 9824
rect 17350 9764 17354 9820
rect 17354 9764 17410 9820
rect 17410 9764 17414 9820
rect 17350 9760 17414 9764
rect 17430 9820 17494 9824
rect 17430 9764 17434 9820
rect 17434 9764 17490 9820
rect 17490 9764 17494 9820
rect 17430 9760 17494 9764
rect 23906 9820 23970 9824
rect 23906 9764 23910 9820
rect 23910 9764 23966 9820
rect 23966 9764 23970 9820
rect 23906 9760 23970 9764
rect 23986 9820 24050 9824
rect 23986 9764 23990 9820
rect 23990 9764 24046 9820
rect 24046 9764 24050 9820
rect 23986 9760 24050 9764
rect 24066 9820 24130 9824
rect 24066 9764 24070 9820
rect 24070 9764 24126 9820
rect 24126 9764 24130 9820
rect 24066 9760 24130 9764
rect 24146 9820 24210 9824
rect 24146 9764 24150 9820
rect 24150 9764 24206 9820
rect 24206 9764 24210 9820
rect 24146 9760 24210 9764
rect 10916 9556 10980 9620
rect 26188 9420 26252 9484
rect 7116 9276 7180 9280
rect 7116 9220 7120 9276
rect 7120 9220 7176 9276
rect 7176 9220 7180 9276
rect 7116 9216 7180 9220
rect 7196 9276 7260 9280
rect 7196 9220 7200 9276
rect 7200 9220 7256 9276
rect 7256 9220 7260 9276
rect 7196 9216 7260 9220
rect 7276 9276 7340 9280
rect 7276 9220 7280 9276
rect 7280 9220 7336 9276
rect 7336 9220 7340 9276
rect 7276 9216 7340 9220
rect 7356 9276 7420 9280
rect 7356 9220 7360 9276
rect 7360 9220 7416 9276
rect 7416 9220 7420 9276
rect 7356 9216 7420 9220
rect 13832 9276 13896 9280
rect 13832 9220 13836 9276
rect 13836 9220 13892 9276
rect 13892 9220 13896 9276
rect 13832 9216 13896 9220
rect 13912 9276 13976 9280
rect 13912 9220 13916 9276
rect 13916 9220 13972 9276
rect 13972 9220 13976 9276
rect 13912 9216 13976 9220
rect 13992 9276 14056 9280
rect 13992 9220 13996 9276
rect 13996 9220 14052 9276
rect 14052 9220 14056 9276
rect 13992 9216 14056 9220
rect 14072 9276 14136 9280
rect 14072 9220 14076 9276
rect 14076 9220 14132 9276
rect 14132 9220 14136 9276
rect 14072 9216 14136 9220
rect 20548 9276 20612 9280
rect 20548 9220 20552 9276
rect 20552 9220 20608 9276
rect 20608 9220 20612 9276
rect 20548 9216 20612 9220
rect 20628 9276 20692 9280
rect 20628 9220 20632 9276
rect 20632 9220 20688 9276
rect 20688 9220 20692 9276
rect 20628 9216 20692 9220
rect 20708 9276 20772 9280
rect 20708 9220 20712 9276
rect 20712 9220 20768 9276
rect 20768 9220 20772 9276
rect 20708 9216 20772 9220
rect 20788 9276 20852 9280
rect 20788 9220 20792 9276
rect 20792 9220 20848 9276
rect 20848 9220 20852 9276
rect 20788 9216 20852 9220
rect 27264 9276 27328 9280
rect 27264 9220 27268 9276
rect 27268 9220 27324 9276
rect 27324 9220 27328 9276
rect 27264 9216 27328 9220
rect 27344 9276 27408 9280
rect 27344 9220 27348 9276
rect 27348 9220 27404 9276
rect 27404 9220 27408 9276
rect 27344 9216 27408 9220
rect 27424 9276 27488 9280
rect 27424 9220 27428 9276
rect 27428 9220 27484 9276
rect 27484 9220 27488 9276
rect 27424 9216 27488 9220
rect 27504 9276 27568 9280
rect 27504 9220 27508 9276
rect 27508 9220 27564 9276
rect 27564 9220 27568 9276
rect 27504 9216 27568 9220
rect 8340 8936 8404 8940
rect 8340 8880 8354 8936
rect 8354 8880 8404 8936
rect 8340 8876 8404 8880
rect 3758 8732 3822 8736
rect 3758 8676 3762 8732
rect 3762 8676 3818 8732
rect 3818 8676 3822 8732
rect 3758 8672 3822 8676
rect 3838 8732 3902 8736
rect 3838 8676 3842 8732
rect 3842 8676 3898 8732
rect 3898 8676 3902 8732
rect 3838 8672 3902 8676
rect 3918 8732 3982 8736
rect 3918 8676 3922 8732
rect 3922 8676 3978 8732
rect 3978 8676 3982 8732
rect 3918 8672 3982 8676
rect 3998 8732 4062 8736
rect 3998 8676 4002 8732
rect 4002 8676 4058 8732
rect 4058 8676 4062 8732
rect 3998 8672 4062 8676
rect 10474 8732 10538 8736
rect 10474 8676 10478 8732
rect 10478 8676 10534 8732
rect 10534 8676 10538 8732
rect 10474 8672 10538 8676
rect 10554 8732 10618 8736
rect 10554 8676 10558 8732
rect 10558 8676 10614 8732
rect 10614 8676 10618 8732
rect 10554 8672 10618 8676
rect 10634 8732 10698 8736
rect 10634 8676 10638 8732
rect 10638 8676 10694 8732
rect 10694 8676 10698 8732
rect 10634 8672 10698 8676
rect 10714 8732 10778 8736
rect 10714 8676 10718 8732
rect 10718 8676 10774 8732
rect 10774 8676 10778 8732
rect 10714 8672 10778 8676
rect 17190 8732 17254 8736
rect 17190 8676 17194 8732
rect 17194 8676 17250 8732
rect 17250 8676 17254 8732
rect 17190 8672 17254 8676
rect 17270 8732 17334 8736
rect 17270 8676 17274 8732
rect 17274 8676 17330 8732
rect 17330 8676 17334 8732
rect 17270 8672 17334 8676
rect 17350 8732 17414 8736
rect 17350 8676 17354 8732
rect 17354 8676 17410 8732
rect 17410 8676 17414 8732
rect 17350 8672 17414 8676
rect 17430 8732 17494 8736
rect 17430 8676 17434 8732
rect 17434 8676 17490 8732
rect 17490 8676 17494 8732
rect 17430 8672 17494 8676
rect 23906 8732 23970 8736
rect 23906 8676 23910 8732
rect 23910 8676 23966 8732
rect 23966 8676 23970 8732
rect 23906 8672 23970 8676
rect 23986 8732 24050 8736
rect 23986 8676 23990 8732
rect 23990 8676 24046 8732
rect 24046 8676 24050 8732
rect 23986 8672 24050 8676
rect 24066 8732 24130 8736
rect 24066 8676 24070 8732
rect 24070 8676 24126 8732
rect 24126 8676 24130 8732
rect 24066 8672 24130 8676
rect 24146 8732 24210 8736
rect 24146 8676 24150 8732
rect 24150 8676 24206 8732
rect 24206 8676 24210 8732
rect 24146 8672 24210 8676
rect 8524 8332 8588 8396
rect 7116 8188 7180 8192
rect 7116 8132 7120 8188
rect 7120 8132 7176 8188
rect 7176 8132 7180 8188
rect 7116 8128 7180 8132
rect 7196 8188 7260 8192
rect 7196 8132 7200 8188
rect 7200 8132 7256 8188
rect 7256 8132 7260 8188
rect 7196 8128 7260 8132
rect 7276 8188 7340 8192
rect 7276 8132 7280 8188
rect 7280 8132 7336 8188
rect 7336 8132 7340 8188
rect 7276 8128 7340 8132
rect 7356 8188 7420 8192
rect 7356 8132 7360 8188
rect 7360 8132 7416 8188
rect 7416 8132 7420 8188
rect 7356 8128 7420 8132
rect 13832 8188 13896 8192
rect 13832 8132 13836 8188
rect 13836 8132 13892 8188
rect 13892 8132 13896 8188
rect 13832 8128 13896 8132
rect 13912 8188 13976 8192
rect 13912 8132 13916 8188
rect 13916 8132 13972 8188
rect 13972 8132 13976 8188
rect 13912 8128 13976 8132
rect 13992 8188 14056 8192
rect 13992 8132 13996 8188
rect 13996 8132 14052 8188
rect 14052 8132 14056 8188
rect 13992 8128 14056 8132
rect 14072 8188 14136 8192
rect 14072 8132 14076 8188
rect 14076 8132 14132 8188
rect 14132 8132 14136 8188
rect 14072 8128 14136 8132
rect 20548 8188 20612 8192
rect 20548 8132 20552 8188
rect 20552 8132 20608 8188
rect 20608 8132 20612 8188
rect 20548 8128 20612 8132
rect 20628 8188 20692 8192
rect 20628 8132 20632 8188
rect 20632 8132 20688 8188
rect 20688 8132 20692 8188
rect 20628 8128 20692 8132
rect 20708 8188 20772 8192
rect 20708 8132 20712 8188
rect 20712 8132 20768 8188
rect 20768 8132 20772 8188
rect 20708 8128 20772 8132
rect 20788 8188 20852 8192
rect 20788 8132 20792 8188
rect 20792 8132 20848 8188
rect 20848 8132 20852 8188
rect 20788 8128 20852 8132
rect 27264 8188 27328 8192
rect 27264 8132 27268 8188
rect 27268 8132 27324 8188
rect 27324 8132 27328 8188
rect 27264 8128 27328 8132
rect 27344 8188 27408 8192
rect 27344 8132 27348 8188
rect 27348 8132 27404 8188
rect 27404 8132 27408 8188
rect 27344 8128 27408 8132
rect 27424 8188 27488 8192
rect 27424 8132 27428 8188
rect 27428 8132 27484 8188
rect 27484 8132 27488 8188
rect 27424 8128 27488 8132
rect 27504 8188 27568 8192
rect 27504 8132 27508 8188
rect 27508 8132 27564 8188
rect 27564 8132 27568 8188
rect 27504 8128 27568 8132
rect 3758 7644 3822 7648
rect 3758 7588 3762 7644
rect 3762 7588 3818 7644
rect 3818 7588 3822 7644
rect 3758 7584 3822 7588
rect 3838 7644 3902 7648
rect 3838 7588 3842 7644
rect 3842 7588 3898 7644
rect 3898 7588 3902 7644
rect 3838 7584 3902 7588
rect 3918 7644 3982 7648
rect 3918 7588 3922 7644
rect 3922 7588 3978 7644
rect 3978 7588 3982 7644
rect 3918 7584 3982 7588
rect 3998 7644 4062 7648
rect 3998 7588 4002 7644
rect 4002 7588 4058 7644
rect 4058 7588 4062 7644
rect 3998 7584 4062 7588
rect 10474 7644 10538 7648
rect 10474 7588 10478 7644
rect 10478 7588 10534 7644
rect 10534 7588 10538 7644
rect 10474 7584 10538 7588
rect 10554 7644 10618 7648
rect 10554 7588 10558 7644
rect 10558 7588 10614 7644
rect 10614 7588 10618 7644
rect 10554 7584 10618 7588
rect 10634 7644 10698 7648
rect 10634 7588 10638 7644
rect 10638 7588 10694 7644
rect 10694 7588 10698 7644
rect 10634 7584 10698 7588
rect 10714 7644 10778 7648
rect 10714 7588 10718 7644
rect 10718 7588 10774 7644
rect 10774 7588 10778 7644
rect 10714 7584 10778 7588
rect 17190 7644 17254 7648
rect 17190 7588 17194 7644
rect 17194 7588 17250 7644
rect 17250 7588 17254 7644
rect 17190 7584 17254 7588
rect 17270 7644 17334 7648
rect 17270 7588 17274 7644
rect 17274 7588 17330 7644
rect 17330 7588 17334 7644
rect 17270 7584 17334 7588
rect 17350 7644 17414 7648
rect 17350 7588 17354 7644
rect 17354 7588 17410 7644
rect 17410 7588 17414 7644
rect 17350 7584 17414 7588
rect 17430 7644 17494 7648
rect 17430 7588 17434 7644
rect 17434 7588 17490 7644
rect 17490 7588 17494 7644
rect 17430 7584 17494 7588
rect 23906 7644 23970 7648
rect 23906 7588 23910 7644
rect 23910 7588 23966 7644
rect 23966 7588 23970 7644
rect 23906 7584 23970 7588
rect 23986 7644 24050 7648
rect 23986 7588 23990 7644
rect 23990 7588 24046 7644
rect 24046 7588 24050 7644
rect 23986 7584 24050 7588
rect 24066 7644 24130 7648
rect 24066 7588 24070 7644
rect 24070 7588 24126 7644
rect 24126 7588 24130 7644
rect 24066 7584 24130 7588
rect 24146 7644 24210 7648
rect 24146 7588 24150 7644
rect 24150 7588 24206 7644
rect 24206 7588 24210 7644
rect 24146 7584 24210 7588
rect 7116 7100 7180 7104
rect 7116 7044 7120 7100
rect 7120 7044 7176 7100
rect 7176 7044 7180 7100
rect 7116 7040 7180 7044
rect 7196 7100 7260 7104
rect 7196 7044 7200 7100
rect 7200 7044 7256 7100
rect 7256 7044 7260 7100
rect 7196 7040 7260 7044
rect 7276 7100 7340 7104
rect 7276 7044 7280 7100
rect 7280 7044 7336 7100
rect 7336 7044 7340 7100
rect 7276 7040 7340 7044
rect 7356 7100 7420 7104
rect 7356 7044 7360 7100
rect 7360 7044 7416 7100
rect 7416 7044 7420 7100
rect 7356 7040 7420 7044
rect 13832 7100 13896 7104
rect 13832 7044 13836 7100
rect 13836 7044 13892 7100
rect 13892 7044 13896 7100
rect 13832 7040 13896 7044
rect 13912 7100 13976 7104
rect 13912 7044 13916 7100
rect 13916 7044 13972 7100
rect 13972 7044 13976 7100
rect 13912 7040 13976 7044
rect 13992 7100 14056 7104
rect 13992 7044 13996 7100
rect 13996 7044 14052 7100
rect 14052 7044 14056 7100
rect 13992 7040 14056 7044
rect 14072 7100 14136 7104
rect 14072 7044 14076 7100
rect 14076 7044 14132 7100
rect 14132 7044 14136 7100
rect 14072 7040 14136 7044
rect 20548 7100 20612 7104
rect 20548 7044 20552 7100
rect 20552 7044 20608 7100
rect 20608 7044 20612 7100
rect 20548 7040 20612 7044
rect 20628 7100 20692 7104
rect 20628 7044 20632 7100
rect 20632 7044 20688 7100
rect 20688 7044 20692 7100
rect 20628 7040 20692 7044
rect 20708 7100 20772 7104
rect 20708 7044 20712 7100
rect 20712 7044 20768 7100
rect 20768 7044 20772 7100
rect 20708 7040 20772 7044
rect 20788 7100 20852 7104
rect 20788 7044 20792 7100
rect 20792 7044 20848 7100
rect 20848 7044 20852 7100
rect 20788 7040 20852 7044
rect 27264 7100 27328 7104
rect 27264 7044 27268 7100
rect 27268 7044 27324 7100
rect 27324 7044 27328 7100
rect 27264 7040 27328 7044
rect 27344 7100 27408 7104
rect 27344 7044 27348 7100
rect 27348 7044 27404 7100
rect 27404 7044 27408 7100
rect 27344 7040 27408 7044
rect 27424 7100 27488 7104
rect 27424 7044 27428 7100
rect 27428 7044 27484 7100
rect 27484 7044 27488 7100
rect 27424 7040 27488 7044
rect 27504 7100 27568 7104
rect 27504 7044 27508 7100
rect 27508 7044 27564 7100
rect 27564 7044 27568 7100
rect 27504 7040 27568 7044
rect 10916 6896 10980 6900
rect 10916 6840 10930 6896
rect 10930 6840 10980 6896
rect 10916 6836 10980 6840
rect 3758 6556 3822 6560
rect 3758 6500 3762 6556
rect 3762 6500 3818 6556
rect 3818 6500 3822 6556
rect 3758 6496 3822 6500
rect 3838 6556 3902 6560
rect 3838 6500 3842 6556
rect 3842 6500 3898 6556
rect 3898 6500 3902 6556
rect 3838 6496 3902 6500
rect 3918 6556 3982 6560
rect 3918 6500 3922 6556
rect 3922 6500 3978 6556
rect 3978 6500 3982 6556
rect 3918 6496 3982 6500
rect 3998 6556 4062 6560
rect 3998 6500 4002 6556
rect 4002 6500 4058 6556
rect 4058 6500 4062 6556
rect 3998 6496 4062 6500
rect 10474 6556 10538 6560
rect 10474 6500 10478 6556
rect 10478 6500 10534 6556
rect 10534 6500 10538 6556
rect 10474 6496 10538 6500
rect 10554 6556 10618 6560
rect 10554 6500 10558 6556
rect 10558 6500 10614 6556
rect 10614 6500 10618 6556
rect 10554 6496 10618 6500
rect 10634 6556 10698 6560
rect 10634 6500 10638 6556
rect 10638 6500 10694 6556
rect 10694 6500 10698 6556
rect 10634 6496 10698 6500
rect 10714 6556 10778 6560
rect 10714 6500 10718 6556
rect 10718 6500 10774 6556
rect 10774 6500 10778 6556
rect 10714 6496 10778 6500
rect 17190 6556 17254 6560
rect 17190 6500 17194 6556
rect 17194 6500 17250 6556
rect 17250 6500 17254 6556
rect 17190 6496 17254 6500
rect 17270 6556 17334 6560
rect 17270 6500 17274 6556
rect 17274 6500 17330 6556
rect 17330 6500 17334 6556
rect 17270 6496 17334 6500
rect 17350 6556 17414 6560
rect 17350 6500 17354 6556
rect 17354 6500 17410 6556
rect 17410 6500 17414 6556
rect 17350 6496 17414 6500
rect 17430 6556 17494 6560
rect 17430 6500 17434 6556
rect 17434 6500 17490 6556
rect 17490 6500 17494 6556
rect 17430 6496 17494 6500
rect 23906 6556 23970 6560
rect 23906 6500 23910 6556
rect 23910 6500 23966 6556
rect 23966 6500 23970 6556
rect 23906 6496 23970 6500
rect 23986 6556 24050 6560
rect 23986 6500 23990 6556
rect 23990 6500 24046 6556
rect 24046 6500 24050 6556
rect 23986 6496 24050 6500
rect 24066 6556 24130 6560
rect 24066 6500 24070 6556
rect 24070 6500 24126 6556
rect 24126 6500 24130 6556
rect 24066 6496 24130 6500
rect 24146 6556 24210 6560
rect 24146 6500 24150 6556
rect 24150 6500 24206 6556
rect 24206 6500 24210 6556
rect 24146 6496 24210 6500
rect 7116 6012 7180 6016
rect 7116 5956 7120 6012
rect 7120 5956 7176 6012
rect 7176 5956 7180 6012
rect 7116 5952 7180 5956
rect 7196 6012 7260 6016
rect 7196 5956 7200 6012
rect 7200 5956 7256 6012
rect 7256 5956 7260 6012
rect 7196 5952 7260 5956
rect 7276 6012 7340 6016
rect 7276 5956 7280 6012
rect 7280 5956 7336 6012
rect 7336 5956 7340 6012
rect 7276 5952 7340 5956
rect 7356 6012 7420 6016
rect 7356 5956 7360 6012
rect 7360 5956 7416 6012
rect 7416 5956 7420 6012
rect 7356 5952 7420 5956
rect 13832 6012 13896 6016
rect 13832 5956 13836 6012
rect 13836 5956 13892 6012
rect 13892 5956 13896 6012
rect 13832 5952 13896 5956
rect 13912 6012 13976 6016
rect 13912 5956 13916 6012
rect 13916 5956 13972 6012
rect 13972 5956 13976 6012
rect 13912 5952 13976 5956
rect 13992 6012 14056 6016
rect 13992 5956 13996 6012
rect 13996 5956 14052 6012
rect 14052 5956 14056 6012
rect 13992 5952 14056 5956
rect 14072 6012 14136 6016
rect 14072 5956 14076 6012
rect 14076 5956 14132 6012
rect 14132 5956 14136 6012
rect 14072 5952 14136 5956
rect 20548 6012 20612 6016
rect 20548 5956 20552 6012
rect 20552 5956 20608 6012
rect 20608 5956 20612 6012
rect 20548 5952 20612 5956
rect 20628 6012 20692 6016
rect 20628 5956 20632 6012
rect 20632 5956 20688 6012
rect 20688 5956 20692 6012
rect 20628 5952 20692 5956
rect 20708 6012 20772 6016
rect 20708 5956 20712 6012
rect 20712 5956 20768 6012
rect 20768 5956 20772 6012
rect 20708 5952 20772 5956
rect 20788 6012 20852 6016
rect 20788 5956 20792 6012
rect 20792 5956 20848 6012
rect 20848 5956 20852 6012
rect 20788 5952 20852 5956
rect 27264 6012 27328 6016
rect 27264 5956 27268 6012
rect 27268 5956 27324 6012
rect 27324 5956 27328 6012
rect 27264 5952 27328 5956
rect 27344 6012 27408 6016
rect 27344 5956 27348 6012
rect 27348 5956 27404 6012
rect 27404 5956 27408 6012
rect 27344 5952 27408 5956
rect 27424 6012 27488 6016
rect 27424 5956 27428 6012
rect 27428 5956 27484 6012
rect 27484 5956 27488 6012
rect 27424 5952 27488 5956
rect 27504 6012 27568 6016
rect 27504 5956 27508 6012
rect 27508 5956 27564 6012
rect 27564 5956 27568 6012
rect 27504 5952 27568 5956
rect 12572 5884 12636 5948
rect 8340 5476 8404 5540
rect 3758 5468 3822 5472
rect 3758 5412 3762 5468
rect 3762 5412 3818 5468
rect 3818 5412 3822 5468
rect 3758 5408 3822 5412
rect 3838 5468 3902 5472
rect 3838 5412 3842 5468
rect 3842 5412 3898 5468
rect 3898 5412 3902 5468
rect 3838 5408 3902 5412
rect 3918 5468 3982 5472
rect 3918 5412 3922 5468
rect 3922 5412 3978 5468
rect 3978 5412 3982 5468
rect 3918 5408 3982 5412
rect 3998 5468 4062 5472
rect 3998 5412 4002 5468
rect 4002 5412 4058 5468
rect 4058 5412 4062 5468
rect 3998 5408 4062 5412
rect 10474 5468 10538 5472
rect 10474 5412 10478 5468
rect 10478 5412 10534 5468
rect 10534 5412 10538 5468
rect 10474 5408 10538 5412
rect 10554 5468 10618 5472
rect 10554 5412 10558 5468
rect 10558 5412 10614 5468
rect 10614 5412 10618 5468
rect 10554 5408 10618 5412
rect 10634 5468 10698 5472
rect 10634 5412 10638 5468
rect 10638 5412 10694 5468
rect 10694 5412 10698 5468
rect 10634 5408 10698 5412
rect 10714 5468 10778 5472
rect 10714 5412 10718 5468
rect 10718 5412 10774 5468
rect 10774 5412 10778 5468
rect 10714 5408 10778 5412
rect 17190 5468 17254 5472
rect 17190 5412 17194 5468
rect 17194 5412 17250 5468
rect 17250 5412 17254 5468
rect 17190 5408 17254 5412
rect 17270 5468 17334 5472
rect 17270 5412 17274 5468
rect 17274 5412 17330 5468
rect 17330 5412 17334 5468
rect 17270 5408 17334 5412
rect 17350 5468 17414 5472
rect 17350 5412 17354 5468
rect 17354 5412 17410 5468
rect 17410 5412 17414 5468
rect 17350 5408 17414 5412
rect 17430 5468 17494 5472
rect 17430 5412 17434 5468
rect 17434 5412 17490 5468
rect 17490 5412 17494 5468
rect 17430 5408 17494 5412
rect 23906 5468 23970 5472
rect 23906 5412 23910 5468
rect 23910 5412 23966 5468
rect 23966 5412 23970 5468
rect 23906 5408 23970 5412
rect 23986 5468 24050 5472
rect 23986 5412 23990 5468
rect 23990 5412 24046 5468
rect 24046 5412 24050 5468
rect 23986 5408 24050 5412
rect 24066 5468 24130 5472
rect 24066 5412 24070 5468
rect 24070 5412 24126 5468
rect 24126 5412 24130 5468
rect 24066 5408 24130 5412
rect 24146 5468 24210 5472
rect 24146 5412 24150 5468
rect 24150 5412 24206 5468
rect 24206 5412 24210 5468
rect 24146 5408 24210 5412
rect 7116 4924 7180 4928
rect 7116 4868 7120 4924
rect 7120 4868 7176 4924
rect 7176 4868 7180 4924
rect 7116 4864 7180 4868
rect 7196 4924 7260 4928
rect 7196 4868 7200 4924
rect 7200 4868 7256 4924
rect 7256 4868 7260 4924
rect 7196 4864 7260 4868
rect 7276 4924 7340 4928
rect 7276 4868 7280 4924
rect 7280 4868 7336 4924
rect 7336 4868 7340 4924
rect 7276 4864 7340 4868
rect 7356 4924 7420 4928
rect 7356 4868 7360 4924
rect 7360 4868 7416 4924
rect 7416 4868 7420 4924
rect 7356 4864 7420 4868
rect 13832 4924 13896 4928
rect 13832 4868 13836 4924
rect 13836 4868 13892 4924
rect 13892 4868 13896 4924
rect 13832 4864 13896 4868
rect 13912 4924 13976 4928
rect 13912 4868 13916 4924
rect 13916 4868 13972 4924
rect 13972 4868 13976 4924
rect 13912 4864 13976 4868
rect 13992 4924 14056 4928
rect 13992 4868 13996 4924
rect 13996 4868 14052 4924
rect 14052 4868 14056 4924
rect 13992 4864 14056 4868
rect 14072 4924 14136 4928
rect 14072 4868 14076 4924
rect 14076 4868 14132 4924
rect 14132 4868 14136 4924
rect 14072 4864 14136 4868
rect 20548 4924 20612 4928
rect 20548 4868 20552 4924
rect 20552 4868 20608 4924
rect 20608 4868 20612 4924
rect 20548 4864 20612 4868
rect 20628 4924 20692 4928
rect 20628 4868 20632 4924
rect 20632 4868 20688 4924
rect 20688 4868 20692 4924
rect 20628 4864 20692 4868
rect 20708 4924 20772 4928
rect 20708 4868 20712 4924
rect 20712 4868 20768 4924
rect 20768 4868 20772 4924
rect 20708 4864 20772 4868
rect 20788 4924 20852 4928
rect 20788 4868 20792 4924
rect 20792 4868 20848 4924
rect 20848 4868 20852 4924
rect 20788 4864 20852 4868
rect 27264 4924 27328 4928
rect 27264 4868 27268 4924
rect 27268 4868 27324 4924
rect 27324 4868 27328 4924
rect 27264 4864 27328 4868
rect 27344 4924 27408 4928
rect 27344 4868 27348 4924
rect 27348 4868 27404 4924
rect 27404 4868 27408 4924
rect 27344 4864 27408 4868
rect 27424 4924 27488 4928
rect 27424 4868 27428 4924
rect 27428 4868 27484 4924
rect 27484 4868 27488 4924
rect 27424 4864 27488 4868
rect 27504 4924 27568 4928
rect 27504 4868 27508 4924
rect 27508 4868 27564 4924
rect 27564 4868 27568 4924
rect 27504 4864 27568 4868
rect 3758 4380 3822 4384
rect 3758 4324 3762 4380
rect 3762 4324 3818 4380
rect 3818 4324 3822 4380
rect 3758 4320 3822 4324
rect 3838 4380 3902 4384
rect 3838 4324 3842 4380
rect 3842 4324 3898 4380
rect 3898 4324 3902 4380
rect 3838 4320 3902 4324
rect 3918 4380 3982 4384
rect 3918 4324 3922 4380
rect 3922 4324 3978 4380
rect 3978 4324 3982 4380
rect 3918 4320 3982 4324
rect 3998 4380 4062 4384
rect 3998 4324 4002 4380
rect 4002 4324 4058 4380
rect 4058 4324 4062 4380
rect 3998 4320 4062 4324
rect 10474 4380 10538 4384
rect 10474 4324 10478 4380
rect 10478 4324 10534 4380
rect 10534 4324 10538 4380
rect 10474 4320 10538 4324
rect 10554 4380 10618 4384
rect 10554 4324 10558 4380
rect 10558 4324 10614 4380
rect 10614 4324 10618 4380
rect 10554 4320 10618 4324
rect 10634 4380 10698 4384
rect 10634 4324 10638 4380
rect 10638 4324 10694 4380
rect 10694 4324 10698 4380
rect 10634 4320 10698 4324
rect 10714 4380 10778 4384
rect 10714 4324 10718 4380
rect 10718 4324 10774 4380
rect 10774 4324 10778 4380
rect 10714 4320 10778 4324
rect 17190 4380 17254 4384
rect 17190 4324 17194 4380
rect 17194 4324 17250 4380
rect 17250 4324 17254 4380
rect 17190 4320 17254 4324
rect 17270 4380 17334 4384
rect 17270 4324 17274 4380
rect 17274 4324 17330 4380
rect 17330 4324 17334 4380
rect 17270 4320 17334 4324
rect 17350 4380 17414 4384
rect 17350 4324 17354 4380
rect 17354 4324 17410 4380
rect 17410 4324 17414 4380
rect 17350 4320 17414 4324
rect 17430 4380 17494 4384
rect 17430 4324 17434 4380
rect 17434 4324 17490 4380
rect 17490 4324 17494 4380
rect 17430 4320 17494 4324
rect 23906 4380 23970 4384
rect 23906 4324 23910 4380
rect 23910 4324 23966 4380
rect 23966 4324 23970 4380
rect 23906 4320 23970 4324
rect 23986 4380 24050 4384
rect 23986 4324 23990 4380
rect 23990 4324 24046 4380
rect 24046 4324 24050 4380
rect 23986 4320 24050 4324
rect 24066 4380 24130 4384
rect 24066 4324 24070 4380
rect 24070 4324 24126 4380
rect 24126 4324 24130 4380
rect 24066 4320 24130 4324
rect 24146 4380 24210 4384
rect 24146 4324 24150 4380
rect 24150 4324 24206 4380
rect 24206 4324 24210 4380
rect 24146 4320 24210 4324
rect 7116 3836 7180 3840
rect 7116 3780 7120 3836
rect 7120 3780 7176 3836
rect 7176 3780 7180 3836
rect 7116 3776 7180 3780
rect 7196 3836 7260 3840
rect 7196 3780 7200 3836
rect 7200 3780 7256 3836
rect 7256 3780 7260 3836
rect 7196 3776 7260 3780
rect 7276 3836 7340 3840
rect 7276 3780 7280 3836
rect 7280 3780 7336 3836
rect 7336 3780 7340 3836
rect 7276 3776 7340 3780
rect 7356 3836 7420 3840
rect 7356 3780 7360 3836
rect 7360 3780 7416 3836
rect 7416 3780 7420 3836
rect 7356 3776 7420 3780
rect 13832 3836 13896 3840
rect 13832 3780 13836 3836
rect 13836 3780 13892 3836
rect 13892 3780 13896 3836
rect 13832 3776 13896 3780
rect 13912 3836 13976 3840
rect 13912 3780 13916 3836
rect 13916 3780 13972 3836
rect 13972 3780 13976 3836
rect 13912 3776 13976 3780
rect 13992 3836 14056 3840
rect 13992 3780 13996 3836
rect 13996 3780 14052 3836
rect 14052 3780 14056 3836
rect 13992 3776 14056 3780
rect 14072 3836 14136 3840
rect 14072 3780 14076 3836
rect 14076 3780 14132 3836
rect 14132 3780 14136 3836
rect 14072 3776 14136 3780
rect 20548 3836 20612 3840
rect 20548 3780 20552 3836
rect 20552 3780 20608 3836
rect 20608 3780 20612 3836
rect 20548 3776 20612 3780
rect 20628 3836 20692 3840
rect 20628 3780 20632 3836
rect 20632 3780 20688 3836
rect 20688 3780 20692 3836
rect 20628 3776 20692 3780
rect 20708 3836 20772 3840
rect 20708 3780 20712 3836
rect 20712 3780 20768 3836
rect 20768 3780 20772 3836
rect 20708 3776 20772 3780
rect 20788 3836 20852 3840
rect 20788 3780 20792 3836
rect 20792 3780 20848 3836
rect 20848 3780 20852 3836
rect 20788 3776 20852 3780
rect 27264 3836 27328 3840
rect 27264 3780 27268 3836
rect 27268 3780 27324 3836
rect 27324 3780 27328 3836
rect 27264 3776 27328 3780
rect 27344 3836 27408 3840
rect 27344 3780 27348 3836
rect 27348 3780 27404 3836
rect 27404 3780 27408 3836
rect 27344 3776 27408 3780
rect 27424 3836 27488 3840
rect 27424 3780 27428 3836
rect 27428 3780 27484 3836
rect 27484 3780 27488 3836
rect 27424 3776 27488 3780
rect 27504 3836 27568 3840
rect 27504 3780 27508 3836
rect 27508 3780 27564 3836
rect 27564 3780 27568 3836
rect 27504 3776 27568 3780
rect 3758 3292 3822 3296
rect 3758 3236 3762 3292
rect 3762 3236 3818 3292
rect 3818 3236 3822 3292
rect 3758 3232 3822 3236
rect 3838 3292 3902 3296
rect 3838 3236 3842 3292
rect 3842 3236 3898 3292
rect 3898 3236 3902 3292
rect 3838 3232 3902 3236
rect 3918 3292 3982 3296
rect 3918 3236 3922 3292
rect 3922 3236 3978 3292
rect 3978 3236 3982 3292
rect 3918 3232 3982 3236
rect 3998 3292 4062 3296
rect 3998 3236 4002 3292
rect 4002 3236 4058 3292
rect 4058 3236 4062 3292
rect 3998 3232 4062 3236
rect 10474 3292 10538 3296
rect 10474 3236 10478 3292
rect 10478 3236 10534 3292
rect 10534 3236 10538 3292
rect 10474 3232 10538 3236
rect 10554 3292 10618 3296
rect 10554 3236 10558 3292
rect 10558 3236 10614 3292
rect 10614 3236 10618 3292
rect 10554 3232 10618 3236
rect 10634 3292 10698 3296
rect 10634 3236 10638 3292
rect 10638 3236 10694 3292
rect 10694 3236 10698 3292
rect 10634 3232 10698 3236
rect 10714 3292 10778 3296
rect 10714 3236 10718 3292
rect 10718 3236 10774 3292
rect 10774 3236 10778 3292
rect 10714 3232 10778 3236
rect 17190 3292 17254 3296
rect 17190 3236 17194 3292
rect 17194 3236 17250 3292
rect 17250 3236 17254 3292
rect 17190 3232 17254 3236
rect 17270 3292 17334 3296
rect 17270 3236 17274 3292
rect 17274 3236 17330 3292
rect 17330 3236 17334 3292
rect 17270 3232 17334 3236
rect 17350 3292 17414 3296
rect 17350 3236 17354 3292
rect 17354 3236 17410 3292
rect 17410 3236 17414 3292
rect 17350 3232 17414 3236
rect 17430 3292 17494 3296
rect 17430 3236 17434 3292
rect 17434 3236 17490 3292
rect 17490 3236 17494 3292
rect 17430 3232 17494 3236
rect 23906 3292 23970 3296
rect 23906 3236 23910 3292
rect 23910 3236 23966 3292
rect 23966 3236 23970 3292
rect 23906 3232 23970 3236
rect 23986 3292 24050 3296
rect 23986 3236 23990 3292
rect 23990 3236 24046 3292
rect 24046 3236 24050 3292
rect 23986 3232 24050 3236
rect 24066 3292 24130 3296
rect 24066 3236 24070 3292
rect 24070 3236 24126 3292
rect 24126 3236 24130 3292
rect 24066 3232 24130 3236
rect 24146 3292 24210 3296
rect 24146 3236 24150 3292
rect 24150 3236 24206 3292
rect 24206 3236 24210 3292
rect 24146 3232 24210 3236
rect 7116 2748 7180 2752
rect 7116 2692 7120 2748
rect 7120 2692 7176 2748
rect 7176 2692 7180 2748
rect 7116 2688 7180 2692
rect 7196 2748 7260 2752
rect 7196 2692 7200 2748
rect 7200 2692 7256 2748
rect 7256 2692 7260 2748
rect 7196 2688 7260 2692
rect 7276 2748 7340 2752
rect 7276 2692 7280 2748
rect 7280 2692 7336 2748
rect 7336 2692 7340 2748
rect 7276 2688 7340 2692
rect 7356 2748 7420 2752
rect 7356 2692 7360 2748
rect 7360 2692 7416 2748
rect 7416 2692 7420 2748
rect 7356 2688 7420 2692
rect 13832 2748 13896 2752
rect 13832 2692 13836 2748
rect 13836 2692 13892 2748
rect 13892 2692 13896 2748
rect 13832 2688 13896 2692
rect 13912 2748 13976 2752
rect 13912 2692 13916 2748
rect 13916 2692 13972 2748
rect 13972 2692 13976 2748
rect 13912 2688 13976 2692
rect 13992 2748 14056 2752
rect 13992 2692 13996 2748
rect 13996 2692 14052 2748
rect 14052 2692 14056 2748
rect 13992 2688 14056 2692
rect 14072 2748 14136 2752
rect 14072 2692 14076 2748
rect 14076 2692 14132 2748
rect 14132 2692 14136 2748
rect 14072 2688 14136 2692
rect 20548 2748 20612 2752
rect 20548 2692 20552 2748
rect 20552 2692 20608 2748
rect 20608 2692 20612 2748
rect 20548 2688 20612 2692
rect 20628 2748 20692 2752
rect 20628 2692 20632 2748
rect 20632 2692 20688 2748
rect 20688 2692 20692 2748
rect 20628 2688 20692 2692
rect 20708 2748 20772 2752
rect 20708 2692 20712 2748
rect 20712 2692 20768 2748
rect 20768 2692 20772 2748
rect 20708 2688 20772 2692
rect 20788 2748 20852 2752
rect 20788 2692 20792 2748
rect 20792 2692 20848 2748
rect 20848 2692 20852 2748
rect 20788 2688 20852 2692
rect 27264 2748 27328 2752
rect 27264 2692 27268 2748
rect 27268 2692 27324 2748
rect 27324 2692 27328 2748
rect 27264 2688 27328 2692
rect 27344 2748 27408 2752
rect 27344 2692 27348 2748
rect 27348 2692 27404 2748
rect 27404 2692 27408 2748
rect 27344 2688 27408 2692
rect 27424 2748 27488 2752
rect 27424 2692 27428 2748
rect 27428 2692 27484 2748
rect 27484 2692 27488 2748
rect 27424 2688 27488 2692
rect 27504 2748 27568 2752
rect 27504 2692 27508 2748
rect 27508 2692 27564 2748
rect 27564 2692 27568 2748
rect 27504 2688 27568 2692
rect 8524 2484 8588 2548
rect 3758 2204 3822 2208
rect 3758 2148 3762 2204
rect 3762 2148 3818 2204
rect 3818 2148 3822 2204
rect 3758 2144 3822 2148
rect 3838 2204 3902 2208
rect 3838 2148 3842 2204
rect 3842 2148 3898 2204
rect 3898 2148 3902 2204
rect 3838 2144 3902 2148
rect 3918 2204 3982 2208
rect 3918 2148 3922 2204
rect 3922 2148 3978 2204
rect 3978 2148 3982 2204
rect 3918 2144 3982 2148
rect 3998 2204 4062 2208
rect 3998 2148 4002 2204
rect 4002 2148 4058 2204
rect 4058 2148 4062 2204
rect 3998 2144 4062 2148
rect 10474 2204 10538 2208
rect 10474 2148 10478 2204
rect 10478 2148 10534 2204
rect 10534 2148 10538 2204
rect 10474 2144 10538 2148
rect 10554 2204 10618 2208
rect 10554 2148 10558 2204
rect 10558 2148 10614 2204
rect 10614 2148 10618 2204
rect 10554 2144 10618 2148
rect 10634 2204 10698 2208
rect 10634 2148 10638 2204
rect 10638 2148 10694 2204
rect 10694 2148 10698 2204
rect 10634 2144 10698 2148
rect 10714 2204 10778 2208
rect 10714 2148 10718 2204
rect 10718 2148 10774 2204
rect 10774 2148 10778 2204
rect 10714 2144 10778 2148
rect 17190 2204 17254 2208
rect 17190 2148 17194 2204
rect 17194 2148 17250 2204
rect 17250 2148 17254 2204
rect 17190 2144 17254 2148
rect 17270 2204 17334 2208
rect 17270 2148 17274 2204
rect 17274 2148 17330 2204
rect 17330 2148 17334 2204
rect 17270 2144 17334 2148
rect 17350 2204 17414 2208
rect 17350 2148 17354 2204
rect 17354 2148 17410 2204
rect 17410 2148 17414 2204
rect 17350 2144 17414 2148
rect 17430 2204 17494 2208
rect 17430 2148 17434 2204
rect 17434 2148 17490 2204
rect 17490 2148 17494 2204
rect 17430 2144 17494 2148
rect 23906 2204 23970 2208
rect 23906 2148 23910 2204
rect 23910 2148 23966 2204
rect 23966 2148 23970 2204
rect 23906 2144 23970 2148
rect 23986 2204 24050 2208
rect 23986 2148 23990 2204
rect 23990 2148 24046 2204
rect 24046 2148 24050 2204
rect 23986 2144 24050 2148
rect 24066 2204 24130 2208
rect 24066 2148 24070 2204
rect 24070 2148 24126 2204
rect 24126 2148 24130 2204
rect 24066 2144 24130 2148
rect 24146 2204 24210 2208
rect 24146 2148 24150 2204
rect 24150 2148 24206 2204
rect 24206 2148 24210 2204
rect 24146 2144 24210 2148
rect 16804 1940 16868 2004
rect 7116 1660 7180 1664
rect 7116 1604 7120 1660
rect 7120 1604 7176 1660
rect 7176 1604 7180 1660
rect 7116 1600 7180 1604
rect 7196 1660 7260 1664
rect 7196 1604 7200 1660
rect 7200 1604 7256 1660
rect 7256 1604 7260 1660
rect 7196 1600 7260 1604
rect 7276 1660 7340 1664
rect 7276 1604 7280 1660
rect 7280 1604 7336 1660
rect 7336 1604 7340 1660
rect 7276 1600 7340 1604
rect 7356 1660 7420 1664
rect 7356 1604 7360 1660
rect 7360 1604 7416 1660
rect 7416 1604 7420 1660
rect 7356 1600 7420 1604
rect 13832 1660 13896 1664
rect 13832 1604 13836 1660
rect 13836 1604 13892 1660
rect 13892 1604 13896 1660
rect 13832 1600 13896 1604
rect 13912 1660 13976 1664
rect 13912 1604 13916 1660
rect 13916 1604 13972 1660
rect 13972 1604 13976 1660
rect 13912 1600 13976 1604
rect 13992 1660 14056 1664
rect 13992 1604 13996 1660
rect 13996 1604 14052 1660
rect 14052 1604 14056 1660
rect 13992 1600 14056 1604
rect 14072 1660 14136 1664
rect 14072 1604 14076 1660
rect 14076 1604 14132 1660
rect 14132 1604 14136 1660
rect 14072 1600 14136 1604
rect 20548 1660 20612 1664
rect 20548 1604 20552 1660
rect 20552 1604 20608 1660
rect 20608 1604 20612 1660
rect 20548 1600 20612 1604
rect 20628 1660 20692 1664
rect 20628 1604 20632 1660
rect 20632 1604 20688 1660
rect 20688 1604 20692 1660
rect 20628 1600 20692 1604
rect 20708 1660 20772 1664
rect 20708 1604 20712 1660
rect 20712 1604 20768 1660
rect 20768 1604 20772 1660
rect 20708 1600 20772 1604
rect 20788 1660 20852 1664
rect 20788 1604 20792 1660
rect 20792 1604 20848 1660
rect 20848 1604 20852 1660
rect 20788 1600 20852 1604
rect 27264 1660 27328 1664
rect 27264 1604 27268 1660
rect 27268 1604 27324 1660
rect 27324 1604 27328 1660
rect 27264 1600 27328 1604
rect 27344 1660 27408 1664
rect 27344 1604 27348 1660
rect 27348 1604 27404 1660
rect 27404 1604 27408 1660
rect 27344 1600 27408 1604
rect 27424 1660 27488 1664
rect 27424 1604 27428 1660
rect 27428 1604 27484 1660
rect 27484 1604 27488 1660
rect 27424 1600 27488 1604
rect 27504 1660 27568 1664
rect 27504 1604 27508 1660
rect 27508 1604 27564 1660
rect 27564 1604 27568 1660
rect 27504 1600 27568 1604
rect 8524 1396 8588 1460
rect 3758 1116 3822 1120
rect 3758 1060 3762 1116
rect 3762 1060 3818 1116
rect 3818 1060 3822 1116
rect 3758 1056 3822 1060
rect 3838 1116 3902 1120
rect 3838 1060 3842 1116
rect 3842 1060 3898 1116
rect 3898 1060 3902 1116
rect 3838 1056 3902 1060
rect 3918 1116 3982 1120
rect 3918 1060 3922 1116
rect 3922 1060 3978 1116
rect 3978 1060 3982 1116
rect 3918 1056 3982 1060
rect 3998 1116 4062 1120
rect 3998 1060 4002 1116
rect 4002 1060 4058 1116
rect 4058 1060 4062 1116
rect 3998 1056 4062 1060
rect 10474 1116 10538 1120
rect 10474 1060 10478 1116
rect 10478 1060 10534 1116
rect 10534 1060 10538 1116
rect 10474 1056 10538 1060
rect 10554 1116 10618 1120
rect 10554 1060 10558 1116
rect 10558 1060 10614 1116
rect 10614 1060 10618 1116
rect 10554 1056 10618 1060
rect 10634 1116 10698 1120
rect 10634 1060 10638 1116
rect 10638 1060 10694 1116
rect 10694 1060 10698 1116
rect 10634 1056 10698 1060
rect 10714 1116 10778 1120
rect 10714 1060 10718 1116
rect 10718 1060 10774 1116
rect 10774 1060 10778 1116
rect 10714 1056 10778 1060
rect 17190 1116 17254 1120
rect 17190 1060 17194 1116
rect 17194 1060 17250 1116
rect 17250 1060 17254 1116
rect 17190 1056 17254 1060
rect 17270 1116 17334 1120
rect 17270 1060 17274 1116
rect 17274 1060 17330 1116
rect 17330 1060 17334 1116
rect 17270 1056 17334 1060
rect 17350 1116 17414 1120
rect 17350 1060 17354 1116
rect 17354 1060 17410 1116
rect 17410 1060 17414 1116
rect 17350 1056 17414 1060
rect 17430 1116 17494 1120
rect 17430 1060 17434 1116
rect 17434 1060 17490 1116
rect 17490 1060 17494 1116
rect 17430 1056 17494 1060
rect 23906 1116 23970 1120
rect 23906 1060 23910 1116
rect 23910 1060 23966 1116
rect 23966 1060 23970 1116
rect 23906 1056 23970 1060
rect 23986 1116 24050 1120
rect 23986 1060 23990 1116
rect 23990 1060 24046 1116
rect 24046 1060 24050 1116
rect 23986 1056 24050 1060
rect 24066 1116 24130 1120
rect 24066 1060 24070 1116
rect 24070 1060 24126 1116
rect 24126 1060 24130 1116
rect 24066 1056 24130 1060
rect 24146 1116 24210 1120
rect 24146 1060 24150 1116
rect 24150 1060 24206 1116
rect 24206 1060 24210 1116
rect 24146 1056 24210 1060
rect 7116 572 7180 576
rect 7116 516 7120 572
rect 7120 516 7176 572
rect 7176 516 7180 572
rect 7116 512 7180 516
rect 7196 572 7260 576
rect 7196 516 7200 572
rect 7200 516 7256 572
rect 7256 516 7260 572
rect 7196 512 7260 516
rect 7276 572 7340 576
rect 7276 516 7280 572
rect 7280 516 7336 572
rect 7336 516 7340 572
rect 7276 512 7340 516
rect 7356 572 7420 576
rect 7356 516 7360 572
rect 7360 516 7416 572
rect 7416 516 7420 572
rect 7356 512 7420 516
rect 13832 572 13896 576
rect 13832 516 13836 572
rect 13836 516 13892 572
rect 13892 516 13896 572
rect 13832 512 13896 516
rect 13912 572 13976 576
rect 13912 516 13916 572
rect 13916 516 13972 572
rect 13972 516 13976 572
rect 13912 512 13976 516
rect 13992 572 14056 576
rect 13992 516 13996 572
rect 13996 516 14052 572
rect 14052 516 14056 572
rect 13992 512 14056 516
rect 14072 572 14136 576
rect 14072 516 14076 572
rect 14076 516 14132 572
rect 14132 516 14136 572
rect 14072 512 14136 516
rect 20548 572 20612 576
rect 20548 516 20552 572
rect 20552 516 20608 572
rect 20608 516 20612 572
rect 20548 512 20612 516
rect 20628 572 20692 576
rect 20628 516 20632 572
rect 20632 516 20688 572
rect 20688 516 20692 572
rect 20628 512 20692 516
rect 20708 572 20772 576
rect 20708 516 20712 572
rect 20712 516 20768 572
rect 20768 516 20772 572
rect 20708 512 20772 516
rect 20788 572 20852 576
rect 20788 516 20792 572
rect 20792 516 20848 572
rect 20848 516 20852 572
rect 20788 512 20852 516
rect 27264 572 27328 576
rect 27264 516 27268 572
rect 27268 516 27324 572
rect 27324 516 27328 572
rect 27264 512 27328 516
rect 27344 572 27408 576
rect 27344 516 27348 572
rect 27348 516 27404 572
rect 27404 516 27408 572
rect 27344 512 27408 516
rect 27424 572 27488 576
rect 27424 516 27428 572
rect 27428 516 27484 572
rect 27484 516 27488 572
rect 27424 512 27488 516
rect 27504 572 27568 576
rect 27504 516 27508 572
rect 27508 516 27564 572
rect 27564 516 27568 572
rect 27504 512 27568 516
<< metal4 >>
rect 3750 17440 4070 17456
rect 3750 17376 3758 17440
rect 3822 17376 3838 17440
rect 3902 17376 3918 17440
rect 3982 17376 3998 17440
rect 4062 17376 4070 17440
rect 3750 16352 4070 17376
rect 3750 16288 3758 16352
rect 3822 16288 3838 16352
rect 3902 16288 3918 16352
rect 3982 16288 3998 16352
rect 4062 16288 4070 16352
rect 3750 15264 4070 16288
rect 3750 15200 3758 15264
rect 3822 15200 3838 15264
rect 3902 15200 3918 15264
rect 3982 15200 3998 15264
rect 4062 15200 4070 15264
rect 3750 14176 4070 15200
rect 3750 14112 3758 14176
rect 3822 14112 3838 14176
rect 3902 14112 3918 14176
rect 3982 14112 3998 14176
rect 4062 14112 4070 14176
rect 3750 13088 4070 14112
rect 3750 13024 3758 13088
rect 3822 13024 3838 13088
rect 3902 13024 3918 13088
rect 3982 13024 3998 13088
rect 4062 13024 4070 13088
rect 3750 12000 4070 13024
rect 3750 11936 3758 12000
rect 3822 11936 3838 12000
rect 3902 11936 3918 12000
rect 3982 11936 3998 12000
rect 4062 11936 4070 12000
rect 3750 10912 4070 11936
rect 3750 10848 3758 10912
rect 3822 10848 3838 10912
rect 3902 10848 3918 10912
rect 3982 10848 3998 10912
rect 4062 10848 4070 10912
rect 3750 9824 4070 10848
rect 3750 9760 3758 9824
rect 3822 9760 3838 9824
rect 3902 9760 3918 9824
rect 3982 9760 3998 9824
rect 4062 9760 4070 9824
rect 3750 8736 4070 9760
rect 3750 8672 3758 8736
rect 3822 8672 3838 8736
rect 3902 8672 3918 8736
rect 3982 8672 3998 8736
rect 4062 8672 4070 8736
rect 3750 7648 4070 8672
rect 3750 7584 3758 7648
rect 3822 7584 3838 7648
rect 3902 7584 3918 7648
rect 3982 7584 3998 7648
rect 4062 7584 4070 7648
rect 3750 6560 4070 7584
rect 3750 6496 3758 6560
rect 3822 6496 3838 6560
rect 3902 6496 3918 6560
rect 3982 6496 3998 6560
rect 4062 6496 4070 6560
rect 3750 5472 4070 6496
rect 3750 5408 3758 5472
rect 3822 5408 3838 5472
rect 3902 5408 3918 5472
rect 3982 5408 3998 5472
rect 4062 5408 4070 5472
rect 3750 4384 4070 5408
rect 3750 4320 3758 4384
rect 3822 4320 3838 4384
rect 3902 4320 3918 4384
rect 3982 4320 3998 4384
rect 4062 4320 4070 4384
rect 3750 3296 4070 4320
rect 3750 3232 3758 3296
rect 3822 3232 3838 3296
rect 3902 3232 3918 3296
rect 3982 3232 3998 3296
rect 4062 3232 4070 3296
rect 3750 2208 4070 3232
rect 3750 2144 3758 2208
rect 3822 2144 3838 2208
rect 3902 2144 3918 2208
rect 3982 2144 3998 2208
rect 4062 2144 4070 2208
rect 3750 1120 4070 2144
rect 3750 1056 3758 1120
rect 3822 1056 3838 1120
rect 3902 1056 3918 1120
rect 3982 1056 3998 1120
rect 4062 1056 4070 1120
rect 3750 496 4070 1056
rect 7108 16896 7428 17456
rect 7108 16832 7116 16896
rect 7180 16832 7196 16896
rect 7260 16832 7276 16896
rect 7340 16832 7356 16896
rect 7420 16832 7428 16896
rect 7108 15808 7428 16832
rect 7108 15744 7116 15808
rect 7180 15744 7196 15808
rect 7260 15744 7276 15808
rect 7340 15744 7356 15808
rect 7420 15744 7428 15808
rect 7108 14720 7428 15744
rect 7108 14656 7116 14720
rect 7180 14656 7196 14720
rect 7260 14656 7276 14720
rect 7340 14656 7356 14720
rect 7420 14656 7428 14720
rect 7108 13632 7428 14656
rect 7108 13568 7116 13632
rect 7180 13568 7196 13632
rect 7260 13568 7276 13632
rect 7340 13568 7356 13632
rect 7420 13568 7428 13632
rect 7108 12544 7428 13568
rect 7108 12480 7116 12544
rect 7180 12480 7196 12544
rect 7260 12480 7276 12544
rect 7340 12480 7356 12544
rect 7420 12480 7428 12544
rect 7108 11456 7428 12480
rect 7108 11392 7116 11456
rect 7180 11392 7196 11456
rect 7260 11392 7276 11456
rect 7340 11392 7356 11456
rect 7420 11392 7428 11456
rect 7108 10368 7428 11392
rect 7108 10304 7116 10368
rect 7180 10304 7196 10368
rect 7260 10304 7276 10368
rect 7340 10304 7356 10368
rect 7420 10304 7428 10368
rect 7108 9280 7428 10304
rect 7108 9216 7116 9280
rect 7180 9216 7196 9280
rect 7260 9216 7276 9280
rect 7340 9216 7356 9280
rect 7420 9216 7428 9280
rect 7108 8192 7428 9216
rect 10466 17440 10786 17456
rect 10466 17376 10474 17440
rect 10538 17376 10554 17440
rect 10618 17376 10634 17440
rect 10698 17376 10714 17440
rect 10778 17376 10786 17440
rect 10466 16352 10786 17376
rect 13824 16896 14144 17456
rect 13824 16832 13832 16896
rect 13896 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14144 16896
rect 12571 16692 12637 16693
rect 12571 16628 12572 16692
rect 12636 16628 12637 16692
rect 12571 16627 12637 16628
rect 10466 16288 10474 16352
rect 10538 16288 10554 16352
rect 10618 16288 10634 16352
rect 10698 16288 10714 16352
rect 10778 16288 10786 16352
rect 10466 15264 10786 16288
rect 10466 15200 10474 15264
rect 10538 15200 10554 15264
rect 10618 15200 10634 15264
rect 10698 15200 10714 15264
rect 10778 15200 10786 15264
rect 10466 14176 10786 15200
rect 10466 14112 10474 14176
rect 10538 14112 10554 14176
rect 10618 14112 10634 14176
rect 10698 14112 10714 14176
rect 10778 14112 10786 14176
rect 10466 13088 10786 14112
rect 10466 13024 10474 13088
rect 10538 13024 10554 13088
rect 10618 13024 10634 13088
rect 10698 13024 10714 13088
rect 10778 13024 10786 13088
rect 10466 12000 10786 13024
rect 10915 12340 10981 12341
rect 10915 12276 10916 12340
rect 10980 12276 10981 12340
rect 10915 12275 10981 12276
rect 10466 11936 10474 12000
rect 10538 11936 10554 12000
rect 10618 11936 10634 12000
rect 10698 11936 10714 12000
rect 10778 11936 10786 12000
rect 10466 10912 10786 11936
rect 10466 10848 10474 10912
rect 10538 10848 10554 10912
rect 10618 10848 10634 10912
rect 10698 10848 10714 10912
rect 10778 10848 10786 10912
rect 10466 9824 10786 10848
rect 10466 9760 10474 9824
rect 10538 9760 10554 9824
rect 10618 9760 10634 9824
rect 10698 9760 10714 9824
rect 10778 9760 10786 9824
rect 8339 8940 8405 8941
rect 8339 8876 8340 8940
rect 8404 8876 8405 8940
rect 8339 8875 8405 8876
rect 7108 8128 7116 8192
rect 7180 8128 7196 8192
rect 7260 8128 7276 8192
rect 7340 8128 7356 8192
rect 7420 8128 7428 8192
rect 7108 7104 7428 8128
rect 7108 7040 7116 7104
rect 7180 7040 7196 7104
rect 7260 7040 7276 7104
rect 7340 7040 7356 7104
rect 7420 7040 7428 7104
rect 7108 6016 7428 7040
rect 7108 5952 7116 6016
rect 7180 5952 7196 6016
rect 7260 5952 7276 6016
rect 7340 5952 7356 6016
rect 7420 5952 7428 6016
rect 7108 4928 7428 5952
rect 8342 5541 8402 8875
rect 10466 8736 10786 9760
rect 10918 9621 10978 12275
rect 10915 9620 10981 9621
rect 10915 9556 10916 9620
rect 10980 9556 10981 9620
rect 10915 9555 10981 9556
rect 10466 8672 10474 8736
rect 10538 8672 10554 8736
rect 10618 8672 10634 8736
rect 10698 8672 10714 8736
rect 10778 8672 10786 8736
rect 8523 8396 8589 8397
rect 8523 8332 8524 8396
rect 8588 8332 8589 8396
rect 8523 8331 8589 8332
rect 8339 5540 8405 5541
rect 8339 5476 8340 5540
rect 8404 5476 8405 5540
rect 8339 5475 8405 5476
rect 7108 4864 7116 4928
rect 7180 4864 7196 4928
rect 7260 4864 7276 4928
rect 7340 4864 7356 4928
rect 7420 4864 7428 4928
rect 7108 3840 7428 4864
rect 7108 3776 7116 3840
rect 7180 3776 7196 3840
rect 7260 3776 7276 3840
rect 7340 3776 7356 3840
rect 7420 3776 7428 3840
rect 7108 2752 7428 3776
rect 7108 2688 7116 2752
rect 7180 2688 7196 2752
rect 7260 2688 7276 2752
rect 7340 2688 7356 2752
rect 7420 2688 7428 2752
rect 7108 1664 7428 2688
rect 8526 2549 8586 8331
rect 10466 7648 10786 8672
rect 10466 7584 10474 7648
rect 10538 7584 10554 7648
rect 10618 7584 10634 7648
rect 10698 7584 10714 7648
rect 10778 7584 10786 7648
rect 10466 6560 10786 7584
rect 10918 6901 10978 9555
rect 10915 6900 10981 6901
rect 10915 6836 10916 6900
rect 10980 6836 10981 6900
rect 10915 6835 10981 6836
rect 10466 6496 10474 6560
rect 10538 6496 10554 6560
rect 10618 6496 10634 6560
rect 10698 6496 10714 6560
rect 10778 6496 10786 6560
rect 10466 5472 10786 6496
rect 12574 5949 12634 16627
rect 13824 15808 14144 16832
rect 17182 17440 17502 17456
rect 17182 17376 17190 17440
rect 17254 17376 17270 17440
rect 17334 17376 17350 17440
rect 17414 17376 17430 17440
rect 17494 17376 17502 17440
rect 16803 16692 16869 16693
rect 16803 16628 16804 16692
rect 16868 16628 16869 16692
rect 16803 16627 16869 16628
rect 13824 15744 13832 15808
rect 13896 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14144 15808
rect 13824 14720 14144 15744
rect 13824 14656 13832 14720
rect 13896 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14144 14720
rect 13824 13632 14144 14656
rect 13824 13568 13832 13632
rect 13896 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14144 13632
rect 13824 12544 14144 13568
rect 13824 12480 13832 12544
rect 13896 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14144 12544
rect 13824 11456 14144 12480
rect 13824 11392 13832 11456
rect 13896 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14144 11456
rect 13824 10368 14144 11392
rect 13824 10304 13832 10368
rect 13896 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14144 10368
rect 13824 9280 14144 10304
rect 13824 9216 13832 9280
rect 13896 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14144 9280
rect 13824 8192 14144 9216
rect 13824 8128 13832 8192
rect 13896 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14144 8192
rect 13824 7104 14144 8128
rect 13824 7040 13832 7104
rect 13896 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14144 7104
rect 13824 6016 14144 7040
rect 13824 5952 13832 6016
rect 13896 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14144 6016
rect 12571 5948 12637 5949
rect 12571 5884 12572 5948
rect 12636 5884 12637 5948
rect 12571 5883 12637 5884
rect 10466 5408 10474 5472
rect 10538 5408 10554 5472
rect 10618 5408 10634 5472
rect 10698 5408 10714 5472
rect 10778 5408 10786 5472
rect 10466 4384 10786 5408
rect 10466 4320 10474 4384
rect 10538 4320 10554 4384
rect 10618 4320 10634 4384
rect 10698 4320 10714 4384
rect 10778 4320 10786 4384
rect 10466 3296 10786 4320
rect 10466 3232 10474 3296
rect 10538 3232 10554 3296
rect 10618 3232 10634 3296
rect 10698 3232 10714 3296
rect 10778 3232 10786 3296
rect 8523 2548 8589 2549
rect 8523 2484 8524 2548
rect 8588 2484 8589 2548
rect 8523 2483 8589 2484
rect 7108 1600 7116 1664
rect 7180 1600 7196 1664
rect 7260 1600 7276 1664
rect 7340 1600 7356 1664
rect 7420 1600 7428 1664
rect 7108 576 7428 1600
rect 8526 1461 8586 2483
rect 10466 2208 10786 3232
rect 10466 2144 10474 2208
rect 10538 2144 10554 2208
rect 10618 2144 10634 2208
rect 10698 2144 10714 2208
rect 10778 2144 10786 2208
rect 8523 1460 8589 1461
rect 8523 1396 8524 1460
rect 8588 1396 8589 1460
rect 8523 1395 8589 1396
rect 7108 512 7116 576
rect 7180 512 7196 576
rect 7260 512 7276 576
rect 7340 512 7356 576
rect 7420 512 7428 576
rect 7108 496 7428 512
rect 10466 1120 10786 2144
rect 10466 1056 10474 1120
rect 10538 1056 10554 1120
rect 10618 1056 10634 1120
rect 10698 1056 10714 1120
rect 10778 1056 10786 1120
rect 10466 496 10786 1056
rect 13824 4928 14144 5952
rect 13824 4864 13832 4928
rect 13896 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14144 4928
rect 13824 3840 14144 4864
rect 13824 3776 13832 3840
rect 13896 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14144 3840
rect 13824 2752 14144 3776
rect 13824 2688 13832 2752
rect 13896 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14144 2752
rect 13824 1664 14144 2688
rect 16806 2005 16866 16627
rect 17182 16352 17502 17376
rect 17182 16288 17190 16352
rect 17254 16288 17270 16352
rect 17334 16288 17350 16352
rect 17414 16288 17430 16352
rect 17494 16288 17502 16352
rect 17182 15264 17502 16288
rect 17182 15200 17190 15264
rect 17254 15200 17270 15264
rect 17334 15200 17350 15264
rect 17414 15200 17430 15264
rect 17494 15200 17502 15264
rect 17182 14176 17502 15200
rect 17182 14112 17190 14176
rect 17254 14112 17270 14176
rect 17334 14112 17350 14176
rect 17414 14112 17430 14176
rect 17494 14112 17502 14176
rect 17182 13088 17502 14112
rect 17182 13024 17190 13088
rect 17254 13024 17270 13088
rect 17334 13024 17350 13088
rect 17414 13024 17430 13088
rect 17494 13024 17502 13088
rect 17182 12000 17502 13024
rect 17182 11936 17190 12000
rect 17254 11936 17270 12000
rect 17334 11936 17350 12000
rect 17414 11936 17430 12000
rect 17494 11936 17502 12000
rect 17182 10912 17502 11936
rect 17182 10848 17190 10912
rect 17254 10848 17270 10912
rect 17334 10848 17350 10912
rect 17414 10848 17430 10912
rect 17494 10848 17502 10912
rect 17182 9824 17502 10848
rect 17182 9760 17190 9824
rect 17254 9760 17270 9824
rect 17334 9760 17350 9824
rect 17414 9760 17430 9824
rect 17494 9760 17502 9824
rect 17182 8736 17502 9760
rect 17182 8672 17190 8736
rect 17254 8672 17270 8736
rect 17334 8672 17350 8736
rect 17414 8672 17430 8736
rect 17494 8672 17502 8736
rect 17182 7648 17502 8672
rect 17182 7584 17190 7648
rect 17254 7584 17270 7648
rect 17334 7584 17350 7648
rect 17414 7584 17430 7648
rect 17494 7584 17502 7648
rect 17182 6560 17502 7584
rect 17182 6496 17190 6560
rect 17254 6496 17270 6560
rect 17334 6496 17350 6560
rect 17414 6496 17430 6560
rect 17494 6496 17502 6560
rect 17182 5472 17502 6496
rect 17182 5408 17190 5472
rect 17254 5408 17270 5472
rect 17334 5408 17350 5472
rect 17414 5408 17430 5472
rect 17494 5408 17502 5472
rect 17182 4384 17502 5408
rect 17182 4320 17190 4384
rect 17254 4320 17270 4384
rect 17334 4320 17350 4384
rect 17414 4320 17430 4384
rect 17494 4320 17502 4384
rect 17182 3296 17502 4320
rect 17182 3232 17190 3296
rect 17254 3232 17270 3296
rect 17334 3232 17350 3296
rect 17414 3232 17430 3296
rect 17494 3232 17502 3296
rect 17182 2208 17502 3232
rect 17182 2144 17190 2208
rect 17254 2144 17270 2208
rect 17334 2144 17350 2208
rect 17414 2144 17430 2208
rect 17494 2144 17502 2208
rect 16803 2004 16869 2005
rect 16803 1940 16804 2004
rect 16868 1940 16869 2004
rect 16803 1939 16869 1940
rect 13824 1600 13832 1664
rect 13896 1600 13912 1664
rect 13976 1600 13992 1664
rect 14056 1600 14072 1664
rect 14136 1600 14144 1664
rect 13824 576 14144 1600
rect 13824 512 13832 576
rect 13896 512 13912 576
rect 13976 512 13992 576
rect 14056 512 14072 576
rect 14136 512 14144 576
rect 13824 496 14144 512
rect 17182 1120 17502 2144
rect 17182 1056 17190 1120
rect 17254 1056 17270 1120
rect 17334 1056 17350 1120
rect 17414 1056 17430 1120
rect 17494 1056 17502 1120
rect 17182 496 17502 1056
rect 20540 16896 20860 17456
rect 20540 16832 20548 16896
rect 20612 16832 20628 16896
rect 20692 16832 20708 16896
rect 20772 16832 20788 16896
rect 20852 16832 20860 16896
rect 20540 15808 20860 16832
rect 20540 15744 20548 15808
rect 20612 15744 20628 15808
rect 20692 15744 20708 15808
rect 20772 15744 20788 15808
rect 20852 15744 20860 15808
rect 20540 14720 20860 15744
rect 20540 14656 20548 14720
rect 20612 14656 20628 14720
rect 20692 14656 20708 14720
rect 20772 14656 20788 14720
rect 20852 14656 20860 14720
rect 20540 13632 20860 14656
rect 20540 13568 20548 13632
rect 20612 13568 20628 13632
rect 20692 13568 20708 13632
rect 20772 13568 20788 13632
rect 20852 13568 20860 13632
rect 20540 12544 20860 13568
rect 20540 12480 20548 12544
rect 20612 12480 20628 12544
rect 20692 12480 20708 12544
rect 20772 12480 20788 12544
rect 20852 12480 20860 12544
rect 20540 11456 20860 12480
rect 20540 11392 20548 11456
rect 20612 11392 20628 11456
rect 20692 11392 20708 11456
rect 20772 11392 20788 11456
rect 20852 11392 20860 11456
rect 20540 10368 20860 11392
rect 20540 10304 20548 10368
rect 20612 10304 20628 10368
rect 20692 10304 20708 10368
rect 20772 10304 20788 10368
rect 20852 10304 20860 10368
rect 20540 9280 20860 10304
rect 20540 9216 20548 9280
rect 20612 9216 20628 9280
rect 20692 9216 20708 9280
rect 20772 9216 20788 9280
rect 20852 9216 20860 9280
rect 20540 8192 20860 9216
rect 20540 8128 20548 8192
rect 20612 8128 20628 8192
rect 20692 8128 20708 8192
rect 20772 8128 20788 8192
rect 20852 8128 20860 8192
rect 20540 7104 20860 8128
rect 20540 7040 20548 7104
rect 20612 7040 20628 7104
rect 20692 7040 20708 7104
rect 20772 7040 20788 7104
rect 20852 7040 20860 7104
rect 20540 6016 20860 7040
rect 20540 5952 20548 6016
rect 20612 5952 20628 6016
rect 20692 5952 20708 6016
rect 20772 5952 20788 6016
rect 20852 5952 20860 6016
rect 20540 4928 20860 5952
rect 20540 4864 20548 4928
rect 20612 4864 20628 4928
rect 20692 4864 20708 4928
rect 20772 4864 20788 4928
rect 20852 4864 20860 4928
rect 20540 3840 20860 4864
rect 20540 3776 20548 3840
rect 20612 3776 20628 3840
rect 20692 3776 20708 3840
rect 20772 3776 20788 3840
rect 20852 3776 20860 3840
rect 20540 2752 20860 3776
rect 20540 2688 20548 2752
rect 20612 2688 20628 2752
rect 20692 2688 20708 2752
rect 20772 2688 20788 2752
rect 20852 2688 20860 2752
rect 20540 1664 20860 2688
rect 20540 1600 20548 1664
rect 20612 1600 20628 1664
rect 20692 1600 20708 1664
rect 20772 1600 20788 1664
rect 20852 1600 20860 1664
rect 20540 576 20860 1600
rect 20540 512 20548 576
rect 20612 512 20628 576
rect 20692 512 20708 576
rect 20772 512 20788 576
rect 20852 512 20860 576
rect 20540 496 20860 512
rect 23898 17440 24218 17456
rect 23898 17376 23906 17440
rect 23970 17376 23986 17440
rect 24050 17376 24066 17440
rect 24130 17376 24146 17440
rect 24210 17376 24218 17440
rect 23898 16352 24218 17376
rect 23898 16288 23906 16352
rect 23970 16288 23986 16352
rect 24050 16288 24066 16352
rect 24130 16288 24146 16352
rect 24210 16288 24218 16352
rect 23898 15264 24218 16288
rect 23898 15200 23906 15264
rect 23970 15200 23986 15264
rect 24050 15200 24066 15264
rect 24130 15200 24146 15264
rect 24210 15200 24218 15264
rect 23898 14176 24218 15200
rect 23898 14112 23906 14176
rect 23970 14112 23986 14176
rect 24050 14112 24066 14176
rect 24130 14112 24146 14176
rect 24210 14112 24218 14176
rect 23898 13088 24218 14112
rect 23898 13024 23906 13088
rect 23970 13024 23986 13088
rect 24050 13024 24066 13088
rect 24130 13024 24146 13088
rect 24210 13024 24218 13088
rect 23898 12000 24218 13024
rect 27256 16896 27576 17456
rect 27256 16832 27264 16896
rect 27328 16832 27344 16896
rect 27408 16832 27424 16896
rect 27488 16832 27504 16896
rect 27568 16832 27576 16896
rect 27256 15808 27576 16832
rect 27256 15744 27264 15808
rect 27328 15744 27344 15808
rect 27408 15744 27424 15808
rect 27488 15744 27504 15808
rect 27568 15744 27576 15808
rect 27256 14720 27576 15744
rect 27256 14656 27264 14720
rect 27328 14656 27344 14720
rect 27408 14656 27424 14720
rect 27488 14656 27504 14720
rect 27568 14656 27576 14720
rect 27256 13632 27576 14656
rect 27256 13568 27264 13632
rect 27328 13568 27344 13632
rect 27408 13568 27424 13632
rect 27488 13568 27504 13632
rect 27568 13568 27576 13632
rect 27256 12544 27576 13568
rect 27256 12480 27264 12544
rect 27328 12480 27344 12544
rect 27408 12480 27424 12544
rect 27488 12480 27504 12544
rect 27568 12480 27576 12544
rect 26187 12340 26253 12341
rect 26187 12276 26188 12340
rect 26252 12276 26253 12340
rect 26187 12275 26253 12276
rect 23898 11936 23906 12000
rect 23970 11936 23986 12000
rect 24050 11936 24066 12000
rect 24130 11936 24146 12000
rect 24210 11936 24218 12000
rect 23898 10912 24218 11936
rect 23898 10848 23906 10912
rect 23970 10848 23986 10912
rect 24050 10848 24066 10912
rect 24130 10848 24146 10912
rect 24210 10848 24218 10912
rect 23898 9824 24218 10848
rect 23898 9760 23906 9824
rect 23970 9760 23986 9824
rect 24050 9760 24066 9824
rect 24130 9760 24146 9824
rect 24210 9760 24218 9824
rect 23898 8736 24218 9760
rect 26190 9485 26250 12275
rect 27256 11456 27576 12480
rect 27256 11392 27264 11456
rect 27328 11392 27344 11456
rect 27408 11392 27424 11456
rect 27488 11392 27504 11456
rect 27568 11392 27576 11456
rect 27256 10368 27576 11392
rect 27256 10304 27264 10368
rect 27328 10304 27344 10368
rect 27408 10304 27424 10368
rect 27488 10304 27504 10368
rect 27568 10304 27576 10368
rect 26187 9484 26253 9485
rect 26187 9420 26188 9484
rect 26252 9420 26253 9484
rect 26187 9419 26253 9420
rect 23898 8672 23906 8736
rect 23970 8672 23986 8736
rect 24050 8672 24066 8736
rect 24130 8672 24146 8736
rect 24210 8672 24218 8736
rect 23898 7648 24218 8672
rect 23898 7584 23906 7648
rect 23970 7584 23986 7648
rect 24050 7584 24066 7648
rect 24130 7584 24146 7648
rect 24210 7584 24218 7648
rect 23898 6560 24218 7584
rect 23898 6496 23906 6560
rect 23970 6496 23986 6560
rect 24050 6496 24066 6560
rect 24130 6496 24146 6560
rect 24210 6496 24218 6560
rect 23898 5472 24218 6496
rect 23898 5408 23906 5472
rect 23970 5408 23986 5472
rect 24050 5408 24066 5472
rect 24130 5408 24146 5472
rect 24210 5408 24218 5472
rect 23898 4384 24218 5408
rect 23898 4320 23906 4384
rect 23970 4320 23986 4384
rect 24050 4320 24066 4384
rect 24130 4320 24146 4384
rect 24210 4320 24218 4384
rect 23898 3296 24218 4320
rect 23898 3232 23906 3296
rect 23970 3232 23986 3296
rect 24050 3232 24066 3296
rect 24130 3232 24146 3296
rect 24210 3232 24218 3296
rect 23898 2208 24218 3232
rect 23898 2144 23906 2208
rect 23970 2144 23986 2208
rect 24050 2144 24066 2208
rect 24130 2144 24146 2208
rect 24210 2144 24218 2208
rect 23898 1120 24218 2144
rect 23898 1056 23906 1120
rect 23970 1056 23986 1120
rect 24050 1056 24066 1120
rect 24130 1056 24146 1120
rect 24210 1056 24218 1120
rect 23898 496 24218 1056
rect 27256 9280 27576 10304
rect 27256 9216 27264 9280
rect 27328 9216 27344 9280
rect 27408 9216 27424 9280
rect 27488 9216 27504 9280
rect 27568 9216 27576 9280
rect 27256 8192 27576 9216
rect 27256 8128 27264 8192
rect 27328 8128 27344 8192
rect 27408 8128 27424 8192
rect 27488 8128 27504 8192
rect 27568 8128 27576 8192
rect 27256 7104 27576 8128
rect 27256 7040 27264 7104
rect 27328 7040 27344 7104
rect 27408 7040 27424 7104
rect 27488 7040 27504 7104
rect 27568 7040 27576 7104
rect 27256 6016 27576 7040
rect 27256 5952 27264 6016
rect 27328 5952 27344 6016
rect 27408 5952 27424 6016
rect 27488 5952 27504 6016
rect 27568 5952 27576 6016
rect 27256 4928 27576 5952
rect 27256 4864 27264 4928
rect 27328 4864 27344 4928
rect 27408 4864 27424 4928
rect 27488 4864 27504 4928
rect 27568 4864 27576 4928
rect 27256 3840 27576 4864
rect 27256 3776 27264 3840
rect 27328 3776 27344 3840
rect 27408 3776 27424 3840
rect 27488 3776 27504 3840
rect 27568 3776 27576 3840
rect 27256 2752 27576 3776
rect 27256 2688 27264 2752
rect 27328 2688 27344 2752
rect 27408 2688 27424 2752
rect 27488 2688 27504 2752
rect 27568 2688 27576 2752
rect 27256 1664 27576 2688
rect 27256 1600 27264 1664
rect 27328 1600 27344 1664
rect 27408 1600 27424 1664
rect 27488 1600 27504 1664
rect 27568 1600 27576 1664
rect 27256 576 27576 1600
rect 27256 512 27264 576
rect 27328 512 27344 576
rect 27408 512 27424 576
rect 27488 512 27504 576
rect 27568 512 27576 576
rect 27256 496 27576 512
use sky130_fd_sc_hd__clkbuf_2  _378_
timestamp -7200
transform 1 0 16100 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _379_
timestamp -7200
transform 1 0 17572 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _380_
timestamp -7200
transform -1 0 5704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _381_
timestamp -7200
transform 1 0 5796 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _382_
timestamp -7200
transform 1 0 5336 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _383_
timestamp -7200
transform 1 0 20056 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp -7200
transform -1 0 3128 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp -7200
transform -1 0 6256 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _386_
timestamp -7200
transform -1 0 6624 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _387_
timestamp -7200
transform -1 0 4692 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _388_
timestamp -7200
transform 1 0 4692 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _389_
timestamp -7200
transform 1 0 15088 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _390_
timestamp -7200
transform -1 0 11224 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _391_
timestamp -7200
transform -1 0 9384 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _392_
timestamp -7200
transform -1 0 6256 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _393_
timestamp -7200
transform 1 0 4968 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _394_
timestamp -7200
transform 1 0 4416 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _395_
timestamp -7200
transform 1 0 4416 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _396_
timestamp -7200
transform -1 0 9936 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _397_
timestamp -7200
transform 1 0 8740 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _398_
timestamp -7200
transform 1 0 6348 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _399_
timestamp -7200
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _400_
timestamp -7200
transform 1 0 8924 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _401_
timestamp -7200
transform 1 0 7544 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _402_
timestamp -7200
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _403_
timestamp -7200
transform -1 0 11868 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _404_
timestamp -7200
transform -1 0 8924 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _405_
timestamp -7200
transform 1 0 8004 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _406_
timestamp -7200
transform -1 0 8648 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _407_
timestamp -7200
transform 1 0 3864 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _408_
timestamp -7200
transform 1 0 3220 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp -7200
transform 1 0 3772 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _410_
timestamp -7200
transform -1 0 5428 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _411_
timestamp -7200
transform 1 0 5428 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _412_
timestamp -7200
transform -1 0 16192 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _413_
timestamp -7200
transform -1 0 15824 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _414_
timestamp -7200
transform -1 0 10396 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _415_
timestamp -7200
transform -1 0 14904 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _416_
timestamp -7200
transform 1 0 7912 0 -1 1632
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_2  _417_
timestamp -7200
transform -1 0 17664 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _418_
timestamp -7200
transform 1 0 6992 0 1 544
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_2  _419_
timestamp -7200
transform -1 0 18492 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _420_
timestamp -7200
transform 1 0 6900 0 1 1632
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_2  _421_
timestamp -7200
transform -1 0 19596 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _422_
timestamp -7200
transform 1 0 6808 0 -1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_2  _423_
timestamp -7200
transform 1 0 19596 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _424_
timestamp -7200
transform -1 0 9108 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _425_
timestamp -7200
transform 1 0 21252 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _426_
timestamp -7200
transform -1 0 10580 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _427_
timestamp -7200
transform 1 0 19596 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _428_
timestamp -7200
transform -1 0 11960 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _429_
timestamp -7200
transform -1 0 20884 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _430_
timestamp -7200
transform 1 0 12512 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp -7200
transform 1 0 15456 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _432_
timestamp -7200
transform 1 0 14260 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _433_
timestamp -7200
transform 1 0 15732 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _434_
timestamp -7200
transform 1 0 17756 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _435_
timestamp -7200
transform 1 0 19044 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _436_
timestamp -7200
transform -1 0 21068 0 -1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _437_
timestamp -7200
transform -1 0 21068 0 -1 1632
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _438_
timestamp -7200
transform -1 0 21528 0 1 1632
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _439_
timestamp -7200
transform -1 0 20240 0 1 1632
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _440_
timestamp -7200
transform -1 0 14720 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _441_
timestamp -7200
transform -1 0 14812 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _442_
timestamp -7200
transform 1 0 16100 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _443_
timestamp -7200
transform 1 0 16100 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _444_
timestamp -7200
transform 1 0 15088 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _445_
timestamp -7200
transform 1 0 15456 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _446_
timestamp -7200
transform 1 0 15180 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _447_
timestamp -7200
transform 1 0 14720 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _448_
timestamp -7200
transform -1 0 13432 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _449_
timestamp -7200
transform 1 0 14628 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _450_
timestamp -7200
transform 1 0 13892 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _451_
timestamp -7200
transform -1 0 13064 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _452_
timestamp -7200
transform 1 0 13800 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _453_
timestamp -7200
transform 1 0 13064 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _454_
timestamp -7200
transform -1 0 12696 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _455_
timestamp -7200
transform 1 0 13156 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _456_
timestamp -7200
transform 1 0 12236 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _457_
timestamp -7200
transform 1 0 12420 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _458_
timestamp -7200
transform 1 0 13524 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _459_
timestamp -7200
transform -1 0 7268 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _460_
timestamp -7200
transform 1 0 12604 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _461_
timestamp -7200
transform -1 0 12420 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp -7200
transform 1 0 13524 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _463_
timestamp -7200
transform 1 0 11776 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _464_
timestamp -7200
transform -1 0 12052 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _465_
timestamp -7200
transform 1 0 4784 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _466_
timestamp -7200
transform 1 0 5336 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _467_
timestamp -7200
transform -1 0 3220 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _468_
timestamp -7200
transform -1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _469_
timestamp -7200
transform 1 0 2484 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _470_
timestamp -7200
transform -1 0 4968 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _471_
timestamp -7200
transform -1 0 23000 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _472_
timestamp -7200
transform -1 0 3680 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _473_
timestamp -7200
transform 1 0 3956 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _474_
timestamp -7200
transform -1 0 4324 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _475_
timestamp -7200
transform 1 0 3312 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _476_
timestamp -7200
transform 1 0 2852 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _477_
timestamp -7200
transform -1 0 5612 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _478_
timestamp -7200
transform 1 0 5796 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _479_
timestamp -7200
transform 1 0 4968 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _480_
timestamp -7200
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _481_
timestamp -7200
transform -1 0 9016 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _482_
timestamp -7200
transform -1 0 24104 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _483_
timestamp -7200
transform 1 0 7452 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _484_
timestamp -7200
transform 1 0 8004 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _485_
timestamp -7200
transform -1 0 10028 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _486_
timestamp -7200
transform 1 0 10028 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _487_
timestamp -7200
transform -1 0 8740 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _488_
timestamp -7200
transform 1 0 10396 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _489_
timestamp -7200
transform -1 0 11408 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _490_
timestamp -7200
transform 1 0 11408 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _491_
timestamp -7200
transform 1 0 19872 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _492_
timestamp -7200
transform -1 0 20976 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _493_
timestamp -7200
transform -1 0 20148 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _494_
timestamp -7200
transform -1 0 24288 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _495_
timestamp -7200
transform -1 0 19688 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _496_
timestamp -7200
transform -1 0 20884 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _497_
timestamp -7200
transform 1 0 17480 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _498_
timestamp -7200
transform 1 0 18216 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _499_
timestamp -7200
transform 1 0 20240 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _500_
timestamp -7200
transform 1 0 19780 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_1  _501_
timestamp -7200
transform -1 0 18584 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _502_
timestamp -7200
transform -1 0 21160 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _503_
timestamp -7200
transform 1 0 22080 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _504_
timestamp -7200
transform 1 0 20332 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _505_
timestamp -7200
transform 1 0 22724 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _506_
timestamp -7200
transform 1 0 23920 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _507_
timestamp -7200
transform -1 0 23736 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _508_
timestamp -7200
transform -1 0 23368 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _509_
timestamp -7200
transform -1 0 25576 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _510_
timestamp -7200
transform 1 0 25576 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _511_
timestamp -7200
transform 1 0 24564 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _512_
timestamp -7200
transform -1 0 25300 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _513_
timestamp -7200
transform -1 0 26220 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _514_
timestamp -7200
transform -1 0 25392 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _515_
timestamp -7200
transform -1 0 24656 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _516_
timestamp -7200
transform -1 0 24472 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _517_
timestamp -7200
transform -1 0 24472 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _518_
timestamp -7200
transform -1 0 23736 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _519_
timestamp -7200
transform 1 0 23920 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _520_
timestamp -7200
transform 1 0 24748 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _521_
timestamp -7200
transform -1 0 24472 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _522_
timestamp -7200
transform 1 0 25208 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _523_
timestamp -7200
transform -1 0 25944 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _524_
timestamp -7200
transform -1 0 21712 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _525_
timestamp -7200
transform -1 0 22724 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _526_
timestamp -7200
transform -1 0 22080 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _527_
timestamp -7200
transform -1 0 23184 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _528_
timestamp -7200
transform 1 0 24012 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _529_
timestamp -7200
transform 1 0 23276 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _530_
timestamp -7200
transform 1 0 23828 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _531_
timestamp -7200
transform 1 0 23828 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _532_
timestamp -7200
transform 1 0 23828 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _533_
timestamp -7200
transform 1 0 24288 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _534_
timestamp -7200
transform -1 0 24932 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _535_
timestamp -7200
transform -1 0 22356 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _536_
timestamp -7200
transform -1 0 21896 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _537_
timestamp -7200
transform 1 0 20516 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _538_
timestamp -7200
transform -1 0 19964 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _539_
timestamp -7200
transform 1 0 19228 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _540_
timestamp -7200
transform 1 0 17940 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _541_
timestamp -7200
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _542_
timestamp -7200
transform -1 0 16836 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _543_
timestamp -7200
transform -1 0 16008 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _544_
timestamp -7200
transform -1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _545_
timestamp -7200
transform 1 0 17572 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _546_
timestamp -7200
transform -1 0 16008 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _547_
timestamp -7200
transform -1 0 4784 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _548_
timestamp -7200
transform 1 0 3220 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _549_
timestamp -7200
transform 1 0 9936 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _550_
timestamp -7200
transform 1 0 6440 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _551_
timestamp -7200
transform 1 0 11224 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _552_
timestamp -7200
transform 1 0 7084 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _553_
timestamp -7200
transform 1 0 6348 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _554_
timestamp -7200
transform -1 0 4968 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _555_
timestamp -7200
transform 1 0 3404 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _556_
timestamp -7200
transform 1 0 3956 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _557_
timestamp -7200
transform 1 0 6624 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _558_
timestamp -7200
transform -1 0 7820 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _559_
timestamp -7200
transform -1 0 4048 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _560_
timestamp -7200
transform 1 0 4232 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _561_
timestamp -7200
transform 1 0 3864 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _562_
timestamp -7200
transform -1 0 6900 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _563_
timestamp -7200
transform -1 0 6532 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _564_
timestamp -7200
transform -1 0 5520 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _565_
timestamp -7200
transform -1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _566_
timestamp -7200
transform 1 0 5060 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _567_
timestamp -7200
transform 1 0 5060 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _568_
timestamp -7200
transform 1 0 6256 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _569_
timestamp -7200
transform -1 0 12328 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _570_
timestamp -7200
transform -1 0 14168 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _571_
timestamp -7200
transform -1 0 13064 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _572_
timestamp -7200
transform 1 0 12328 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _573_
timestamp -7200
transform 1 0 10396 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _574_
timestamp -7200
transform -1 0 11776 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _575_
timestamp -7200
transform 1 0 11776 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _576_
timestamp -7200
transform -1 0 14536 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _577_
timestamp -7200
transform 1 0 12880 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _578_
timestamp -7200
transform -1 0 15088 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _579_
timestamp -7200
transform 1 0 10948 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _580_
timestamp -7200
transform 1 0 9476 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _581_
timestamp -7200
transform 1 0 10028 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _582_
timestamp -7200
transform 1 0 9752 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _583_
timestamp -7200
transform 1 0 10120 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _584_
timestamp -7200
transform 1 0 9384 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _585_
timestamp -7200
transform 1 0 8464 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _586_
timestamp -7200
transform 1 0 8924 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _587_
timestamp -7200
transform 1 0 6532 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _588_
timestamp -7200
transform 1 0 7912 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _589_
timestamp -7200
transform 1 0 9936 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _590_
timestamp -7200
transform 1 0 6072 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _591_
timestamp -7200
transform 1 0 7176 0 1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _592_
timestamp -7200
transform 1 0 9660 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _593_
timestamp -7200
transform -1 0 16928 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _594_
timestamp -7200
transform -1 0 12144 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _595_
timestamp -7200
transform 1 0 9844 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _596_
timestamp -7200
transform -1 0 9752 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _597_
timestamp -7200
transform -1 0 9016 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _598_
timestamp -7200
transform -1 0 9292 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _599_
timestamp -7200
transform -1 0 10120 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _600_
timestamp -7200
transform -1 0 9660 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _601_
timestamp -7200
transform -1 0 9844 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _602_
timestamp -7200
transform -1 0 9660 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _603_
timestamp -7200
transform 1 0 8188 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _604_
timestamp -7200
transform -1 0 9476 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _605_
timestamp -7200
transform -1 0 8924 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _606_
timestamp -7200
transform 1 0 8096 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _607_
timestamp -7200
transform 1 0 12696 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _608_
timestamp -7200
transform -1 0 15180 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _609_
timestamp -7200
transform 1 0 12972 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _610_
timestamp -7200
transform -1 0 15916 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _611_
timestamp -7200
transform 1 0 11316 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _612_
timestamp -7200
transform 1 0 12052 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _613_
timestamp -7200
transform -1 0 13432 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _614_
timestamp -7200
transform -1 0 13156 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _615_
timestamp -7200
transform 1 0 14628 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _616_
timestamp -7200
transform -1 0 16008 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _617_
timestamp -7200
transform 1 0 20148 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _618_
timestamp -7200
transform 1 0 17572 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _619_
timestamp -7200
transform -1 0 19044 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _620_
timestamp -7200
transform 1 0 17296 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _621_
timestamp -7200
transform 1 0 18216 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _622_
timestamp -7200
transform 1 0 20608 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _623_
timestamp -7200
transform 1 0 19504 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _624_
timestamp -7200
transform 1 0 16100 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _625_
timestamp -7200
transform 1 0 16836 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _626_
timestamp -7200
transform 1 0 23828 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _627_
timestamp -7200
transform -1 0 26036 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _628_
timestamp -7200
transform -1 0 26772 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _629_
timestamp -7200
transform 1 0 24564 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _630_
timestamp -7200
transform -1 0 26036 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _631_
timestamp -7200
transform -1 0 26036 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _632_
timestamp -7200
transform 1 0 26404 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _633_
timestamp -7200
transform -1 0 25208 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _634_
timestamp -7200
transform 1 0 26404 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _635_
timestamp -7200
transform -1 0 24564 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _636_
timestamp -7200
transform -1 0 23460 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _637_
timestamp -7200
transform 1 0 22264 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _638_
timestamp -7200
transform -1 0 23460 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _639_
timestamp -7200
transform -1 0 21068 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _640_
timestamp -7200
transform -1 0 21988 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _641_
timestamp -7200
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _642_
timestamp -7200
transform -1 0 20884 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _643_
timestamp -7200
transform 1 0 18676 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _644_
timestamp -7200
transform -1 0 18584 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _645_
timestamp -7200
transform 1 0 6808 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _646_
timestamp -7200
transform -1 0 16008 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _647_
timestamp -7200
transform -1 0 16836 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _648_
timestamp -7200
transform 1 0 13800 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _649_
timestamp -7200
transform -1 0 14720 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _650_
timestamp -7200
transform 1 0 11868 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _651_
timestamp -7200
transform -1 0 7544 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _652_
timestamp -7200
transform 1 0 10120 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _653_
timestamp -7200
transform -1 0 11684 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _654_
timestamp -7200
transform 1 0 8372 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _655_
timestamp -7200
transform 1 0 6164 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _656_
timestamp -7200
transform -1 0 7636 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _657_
timestamp -7200
transform 1 0 6256 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _658_
timestamp -7200
transform -1 0 7544 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _659_
timestamp -7200
transform 1 0 8924 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _660_
timestamp -7200
transform 1 0 6900 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _661_
timestamp -7200
transform 1 0 8924 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _662_
timestamp -7200
transform 1 0 5704 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _663_
timestamp -7200
transform -1 0 11592 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _664_
timestamp -7200
transform -1 0 11960 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _665_
timestamp -7200
transform -1 0 11224 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _666_
timestamp -7200
transform -1 0 14260 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _667_
timestamp -7200
transform 1 0 10672 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _668_
timestamp -7200
transform 1 0 19872 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _669_
timestamp -7200
transform 1 0 12696 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _670_
timestamp -7200
transform 1 0 19504 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _671_
timestamp -7200
transform 1 0 11960 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _672_
timestamp -7200
transform 1 0 13892 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _673_
timestamp -7200
transform 1 0 18400 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _674_
timestamp -7200
transform 1 0 13524 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _675_
timestamp -7200
transform 1 0 16928 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _676_
timestamp -7200
transform 1 0 18952 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _677_
timestamp -7200
transform -1 0 18400 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _678_
timestamp -7200
transform -1 0 20884 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _679_
timestamp -7200
transform -1 0 20976 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _680_
timestamp -7200
transform 1 0 23092 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _681_
timestamp -7200
transform -1 0 23460 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _682_
timestamp -7200
transform -1 0 24840 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _683_
timestamp -7200
transform -1 0 25024 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _684_
timestamp -7200
transform -1 0 24288 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _685_
timestamp -7200
transform -1 0 27140 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _686_
timestamp -7200
transform -1 0 26956 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _687_
timestamp -7200
transform -1 0 25576 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _688_
timestamp -7200
transform 1 0 24656 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _689_
timestamp -7200
transform -1 0 25300 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _690_
timestamp -7200
transform 1 0 21252 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _691_
timestamp -7200
transform 1 0 20056 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _692_
timestamp -7200
transform -1 0 21620 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _693_
timestamp -7200
transform -1 0 21160 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _694_
timestamp -7200
transform -1 0 22816 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _695_
timestamp -7200
transform 1 0 18768 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _696_
timestamp -7200
transform 1 0 20332 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _697_
timestamp -7200
transform -1 0 20608 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _698_
timestamp -7200
transform 1 0 19412 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _699_
timestamp -7200
transform -1 0 19688 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _700_
timestamp -7200
transform 1 0 18676 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _701_
timestamp -7200
transform -1 0 18216 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _702_
timestamp -7200
transform -1 0 16652 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _703_
timestamp -7200
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _704_
timestamp -7200
transform 1 0 15180 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _705_
timestamp -7200
transform 1 0 14628 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _706_
timestamp -7200
transform -1 0 5704 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _707_
timestamp -7200
transform -1 0 5428 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _708_
timestamp -7200
transform 1 0 5428 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _709_
timestamp -7200
transform 1 0 5796 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _710_
timestamp -7200
transform -1 0 4692 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _711_
timestamp -7200
transform -1 0 5612 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _712_
timestamp -7200
transform -1 0 6256 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _713_
timestamp -7200
transform -1 0 4784 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _714_
timestamp -7200
transform -1 0 8924 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _715_
timestamp -7200
transform 1 0 9108 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _716_
timestamp -7200
transform 1 0 8096 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _717_
timestamp -7200
transform 1 0 6348 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _718_
timestamp -7200
transform 1 0 7544 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _719_
timestamp -7200
transform 1 0 6624 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _720_
timestamp -7200
transform 1 0 6992 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _721_
timestamp -7200
transform 1 0 3680 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _722_
timestamp -7200
transform 1 0 7544 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _723_
timestamp -7200
transform 1 0 4692 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _724_
timestamp -7200
transform 1 0 13524 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _725_
timestamp -7200
transform 1 0 10120 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _726_
timestamp -7200
transform 1 0 12420 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _727_
timestamp -7200
transform -1 0 11500 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _728_
timestamp -7200
transform 1 0 11684 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _729_
timestamp -7200
transform -1 0 12236 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _730_
timestamp -7200
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _731_
timestamp -7200
transform 1 0 3864 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _732_
timestamp -7200
transform -1 0 8280 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _733_
timestamp -7200
transform -1 0 10304 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _734_
timestamp -7200
transform 1 0 8464 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _735_
timestamp -7200
transform -1 0 5520 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _736_
timestamp -7200
transform -1 0 6808 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _737_
timestamp -7200
transform 1 0 6164 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _738_
timestamp -7200
transform 1 0 6624 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _739_
timestamp -7200
transform -1 0 5796 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _740_
timestamp -7200
transform -1 0 5428 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _741_
timestamp -7200
transform 1 0 4876 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _742_
timestamp -7200
transform -1 0 4508 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _743_
timestamp -7200
transform -1 0 3864 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _744_
timestamp -7200
transform 1 0 2760 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _745_
timestamp -7200
transform -1 0 5152 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _746_
timestamp -7200
transform -1 0 4232 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _747_
timestamp -7200
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _748_
timestamp -7200
transform 1 0 14352 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _749_
timestamp -7200
transform -1 0 11316 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _750_
timestamp -7200
transform -1 0 10764 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _751_
timestamp -7200
transform 1 0 10212 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _752_
timestamp -7200
transform 1 0 11868 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _753_
timestamp -7200
transform 1 0 12236 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _754_
timestamp -7200
transform -1 0 12880 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _755_
timestamp -7200
transform -1 0 13064 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _756_
timestamp -7200
transform -1 0 11868 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _757_
timestamp -7200
transform 1 0 11316 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _758_
timestamp -7200
transform 1 0 13800 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _759_
timestamp -7200
transform 1 0 14444 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _760_
timestamp -7200
transform -1 0 15180 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _761_
timestamp -7200
transform 1 0 16468 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _762_
timestamp -7200
transform 1 0 16744 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _763_
timestamp -7200
transform -1 0 17480 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _764_
timestamp -7200
transform 1 0 15824 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _765_
timestamp -7200
transform 1 0 16284 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _766_
timestamp -7200
transform -1 0 17756 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _767_
timestamp -7200
transform 1 0 16192 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _768_
timestamp -7200
transform 1 0 17296 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _769_
timestamp -7200
transform -1 0 18124 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _770_
timestamp -7200
transform 1 0 16836 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _771_
timestamp -7200
transform 1 0 18584 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _772_
timestamp -7200
transform -1 0 19596 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _773_
timestamp -7200
transform 1 0 16652 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _774_
timestamp -7200
transform 1 0 18676 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _775_
timestamp -7200
transform -1 0 20516 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _776_
timestamp -7200
transform 1 0 16928 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _777_
timestamp -7200
transform 1 0 17664 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _778_
timestamp -7200
transform -1 0 18584 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _779_
timestamp -7200
transform 1 0 13708 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _780_
timestamp -7200
transform 1 0 16100 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _781_
timestamp -7200
transform -1 0 16836 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _782_
timestamp -7200
transform 1 0 1564 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _783_
timestamp -7200
transform 1 0 1840 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _784_
timestamp -7200
transform 1 0 2484 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _785_
timestamp -7200
transform 1 0 4140 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _786_
timestamp -7200
transform 1 0 6532 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _787_
timestamp -7200
transform 1 0 8464 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _788_
timestamp -7200
transform -1 0 11500 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _789_
timestamp -7200
transform 1 0 20424 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _790_
timestamp -7200
transform 1 0 17756 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _791_
timestamp -7200
transform 1 0 17572 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _792_
timestamp -7200
transform -1 0 22448 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _793_
timestamp -7200
transform 1 0 23828 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _794_
timestamp -7200
transform 1 0 25300 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _795_
timestamp -7200
transform 1 0 24472 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _796_
timestamp -7200
transform 1 0 24472 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _797_
timestamp -7200
transform 1 0 25484 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _798_
timestamp -7200
transform 1 0 21436 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _799_
timestamp -7200
transform -1 0 23736 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _800_
timestamp -7200
transform 1 0 24840 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _801_
timestamp -7200
transform -1 0 21620 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _802_
timestamp -7200
transform 1 0 18676 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _803_
timestamp -7200
transform 1 0 16100 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _804_
timestamp -7200
transform -1 0 17572 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _805_
timestamp -7200
transform 1 0 4784 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _806_
timestamp -7200
transform 1 0 1656 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _807_
timestamp -7200
transform 1 0 8372 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _808_
timestamp -7200
transform 1 0 8556 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _809_
timestamp -7200
transform 1 0 1656 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _810_
timestamp -7200
transform 1 0 1748 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _811_
timestamp -7200
transform 1 0 6072 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _812_
timestamp -7200
transform 1 0 3128 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _813_
timestamp -7200
transform 1 0 1380 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _814_
timestamp -7200
transform 1 0 13064 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _815_
timestamp -7200
transform 1 0 12788 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _816_
timestamp -7200
transform -1 0 16008 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _817_
timestamp -7200
transform 1 0 9292 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _818_
timestamp -7200
transform 1 0 7728 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _819_
timestamp -7200
transform 1 0 11500 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _820_
timestamp -7200
transform 1 0 8556 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _821_
timestamp -7200
transform 1 0 9108 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _822_
timestamp -7200
transform 1 0 8832 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _823_
timestamp -7200
transform 1 0 8832 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _824_
timestamp -7200
transform 1 0 15088 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _825_
timestamp -7200
transform 1 0 16100 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _826_
timestamp -7200
transform 1 0 11960 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _827_
timestamp -7200
transform 1 0 13524 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _828_
timestamp -7200
transform 1 0 15180 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _829_
timestamp -7200
transform 1 0 16928 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _830_
timestamp -7200
transform 1 0 19228 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _831_
timestamp -7200
transform 1 0 23000 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _832_
timestamp -7200
transform 1 0 24564 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _833_
timestamp -7200
transform 1 0 25484 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _834_
timestamp -7200
transform 1 0 24288 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _835_
timestamp -7200
transform -1 0 25944 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _836_
timestamp -7200
transform 1 0 21068 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _837_
timestamp -7200
transform -1 0 22724 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _838_
timestamp -7200
transform 1 0 18860 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _839_
timestamp -7200
transform 1 0 17388 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _840_
timestamp -7200
transform 1 0 14904 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _841_
timestamp -7200
transform 1 0 13524 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _842_
timestamp -7200
transform 1 0 11408 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _843_
timestamp -7200
transform -1 0 11500 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _844_
timestamp -7200
transform 1 0 6900 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _845_
timestamp -7200
transform 1 0 7268 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _846_
timestamp -7200
transform 1 0 5428 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _847_
timestamp -7200
transform 1 0 6164 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _848_
timestamp -7200
transform 1 0 11500 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _849_
timestamp -7200
transform -1 0 14996 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _850_
timestamp -7200
transform -1 0 11960 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _851_
timestamp -7200
transform 1 0 11132 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _852_
timestamp -7200
transform 1 0 13156 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _853_
timestamp -7200
transform -1 0 18768 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _854_
timestamp -7200
transform -1 0 21344 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _855_
timestamp -7200
transform 1 0 22172 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _856_
timestamp -7200
transform 1 0 24104 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _857_
timestamp -7200
transform 1 0 25024 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _858_
timestamp -7200
transform 1 0 25484 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _859_
timestamp -7200
transform 1 0 24840 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _860_
timestamp -7200
transform 1 0 21252 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _861_
timestamp -7200
transform 1 0 20608 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _862_
timestamp -7200
transform -1 0 22724 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _863_
timestamp -7200
transform 1 0 17848 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _864_
timestamp -7200
transform 1 0 17112 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _865_
timestamp -7200
transform 1 0 15088 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _866_
timestamp -7200
transform -1 0 15272 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _867_
timestamp -7200
transform 1 0 2944 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _868_
timestamp -7200
transform -1 0 9200 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _869_
timestamp -7200
transform 1 0 5888 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _870_
timestamp -7200
transform 1 0 4232 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _871_
timestamp -7200
transform 1 0 3036 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _872_
timestamp -7200
transform 1 0 4140 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _873_
timestamp -7200
transform 1 0 9384 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _874_
timestamp -7200
transform 1 0 10948 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _875_
timestamp -7200
transform 1 0 10948 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _876_
timestamp -7200
transform 1 0 2576 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _877_
timestamp -7200
transform 1 0 8372 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _878_
timestamp -7200
transform 1 0 5796 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _879_
timestamp -7200
transform 1 0 4508 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _880_
timestamp -7200
transform 1 0 1656 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _881_
timestamp -7200
transform 1 0 3220 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _882_
timestamp -7200
transform 1 0 9384 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _883_
timestamp -7200
transform 1 0 12512 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _884_
timestamp -7200
transform 1 0 10948 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _885_
timestamp -7200
transform -1 0 15456 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _886_
timestamp -7200
transform -1 0 17756 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _887_
timestamp -7200
transform -1 0 18124 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _888_
timestamp -7200
transform 1 0 18124 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _889_
timestamp -7200
transform -1 0 21068 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _890_
timestamp -7200
transform -1 0 21068 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _891_
timestamp -7200
transform 1 0 18768 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _892_
timestamp -7200
transform 1 0 16560 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  _903_
timestamp -7200
transform 1 0 4416 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _904_
timestamp -7200
transform 1 0 8372 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _905_
timestamp -7200
transform 1 0 5888 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _906_
timestamp -7200
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -7200
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -7200
transform -1 0 16100 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp -7200
transform -1 0 7912 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp -7200
transform -1 0 10856 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp -7200
transform 1 0 6624 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp -7200
transform 1 0 10948 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp -7200
transform -1 0 20516 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp -7200
transform 1 0 21712 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp -7200
transform -1 0 20516 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp -7200
transform 1 0 21988 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  digital_top_14
timestamp -7200
transform -1 0 4324 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_15
timestamp -7200
transform -1 0 1748 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_16
timestamp -7200
transform -1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_17
timestamp -7200
transform -1 0 9476 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_18
timestamp -7200
transform -1 0 7084 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_19
timestamp -7200
transform 1 0 5428 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_20
timestamp -7200
transform -1 0 5428 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_21
timestamp -7200
transform 1 0 4692 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_22
timestamp -7200
transform 1 0 3404 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_23
timestamp -7200
transform 1 0 2760 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp -7200
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp -7200
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp -7200
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp -7200
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp -7200
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp -7200
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp -7200
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_69
timestamp -7200
transform 1 0 6900 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_93
timestamp -7200
transform 1 0 9108 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp -7200
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113
timestamp -7200
transform 1 0 10948 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_124
timestamp -7200
transform 1 0 11960 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138
timestamp -7200
transform 1 0 13248 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp -7200
transform 1 0 13524 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_157
timestamp -7200
transform 1 0 14996 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp -7200
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp -7200
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp -7200
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp -7200
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp -7200
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp -7200
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp -7200
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp -7200
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp -7200
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp -7200
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp -7200
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp -7200
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp -7200
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_281
timestamp -7200
transform 1 0 26404 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp -7200
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp -7200
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp -7200
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_39
timestamp -7200
transform 1 0 4140 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_50
timestamp -7200
transform 1 0 5152 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_73
timestamp -7200
transform 1 0 7268 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_79
timestamp -7200
transform 1 0 7820 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_94
timestamp -7200
transform 1 0 9200 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_129
timestamp -7200
transform 1 0 12420 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_165
timestamp -7200
transform 1 0 15732 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp -7200
transform 1 0 16100 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_195
timestamp -7200
transform 1 0 18492 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp -7200
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp -7200
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp -7200
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp -7200
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp -7200
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp -7200
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp -7200
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_281
timestamp -7200
transform 1 0 26404 0 -1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp -7200
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp -7200
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp -7200
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp -7200
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_41
timestamp -7200
transform 1 0 4324 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_59
timestamp -7200
transform 1 0 5980 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp -7200
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_101
timestamp -7200
transform 1 0 9844 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_108
timestamp -7200
transform 1 0 10488 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_116
timestamp -7200
transform 1 0 11224 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_120
timestamp -7200
transform 1 0 11592 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_128
timestamp -7200
transform 1 0 12328 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_134
timestamp -7200
transform 1 0 12880 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_141
timestamp -7200
transform 1 0 13524 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_159
timestamp -7200
transform 1 0 15180 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_173
timestamp -7200
transform 1 0 16468 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_191
timestamp -7200
transform 1 0 18124 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp -7200
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_197
timestamp -7200
transform 1 0 18676 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_228
timestamp -7200
transform 1 0 21528 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_240
timestamp -7200
transform 1 0 22632 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp -7200
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp -7200
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp -7200
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp -7200
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp -7200
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_27
timestamp -7200
transform 1 0 3036 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_33
timestamp -7200
transform 1 0 3588 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_37
timestamp -7200
transform 1 0 3956 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_45
timestamp -7200
transform 1 0 4692 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_53
timestamp -7200
transform 1 0 5428 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_57
timestamp -7200
transform 1 0 5796 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_82
timestamp -7200
transform 1 0 8096 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_89
timestamp -7200
transform 1 0 8740 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_101
timestamp -7200
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_105
timestamp -7200
transform 1 0 10212 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp -7200
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_113
timestamp -7200
transform 1 0 10948 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_117
timestamp -7200
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_123
timestamp -7200
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_132
timestamp -7200
transform 1 0 12696 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_144
timestamp -7200
transform 1 0 13800 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_154
timestamp -7200
transform 1 0 14720 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp -7200
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_169
timestamp -7200
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_187
timestamp -7200
transform 1 0 17756 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_199
timestamp -7200
transform 1 0 18860 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_207
timestamp -7200
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp -7200
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp -7200
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp -7200
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp -7200
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp -7200
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp -7200
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp -7200
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_281
timestamp -7200
transform 1 0 26404 0 -1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp -7200
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp -7200
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp -7200
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_45
timestamp -7200
transform 1 0 4692 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_49
timestamp -7200
transform 1 0 5060 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_57
timestamp -7200
transform 1 0 5796 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_74
timestamp -7200
transform 1 0 7360 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_106
timestamp -7200
transform 1 0 10304 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_117
timestamp -7200
transform 1 0 11316 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_130
timestamp -7200
transform 1 0 12512 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp -7200
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_156
timestamp -7200
transform 1 0 14904 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_164
timestamp -7200
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_180
timestamp -7200
transform 1 0 17112 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_192
timestamp -7200
transform 1 0 18216 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_197
timestamp -7200
transform 1 0 18676 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_217
timestamp -7200
transform 1 0 20516 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_229
timestamp -7200
transform 1 0 21620 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_241
timestamp -7200
transform 1 0 22724 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_249
timestamp -7200
transform 1 0 23460 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp -7200
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp -7200
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp -7200
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp -7200
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_15
timestamp -7200
transform 1 0 1932 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_23
timestamp -7200
transform 1 0 2668 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_27
timestamp -7200
transform 1 0 3036 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp -7200
transform 1 0 5796 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_74
timestamp -7200
transform 1 0 7360 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_94
timestamp -7200
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_136
timestamp -7200
transform 1 0 13064 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_155
timestamp -7200
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_185
timestamp -7200
transform 1 0 17572 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp -7200
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp -7200
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp -7200
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp -7200
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp -7200
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp -7200
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp -7200
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_281
timestamp -7200
transform 1 0 26404 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_3
timestamp -7200
transform 1 0 828 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_11
timestamp -7200
transform 1 0 1564 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp -7200
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_54
timestamp -7200
transform 1 0 5520 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_62
timestamp -7200
transform 1 0 6256 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_79
timestamp -7200
transform 1 0 7820 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp -7200
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_91
timestamp -7200
transform 1 0 8924 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_135
timestamp -7200
transform 1 0 12972 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp -7200
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_147
timestamp -7200
transform 1 0 14076 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_159
timestamp -7200
transform 1 0 15180 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_171
timestamp -7200
transform 1 0 16284 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_187
timestamp -7200
transform 1 0 17756 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_191
timestamp -7200
transform 1 0 18124 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp -7200
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_202
timestamp -7200
transform 1 0 19136 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_223
timestamp -7200
transform 1 0 21068 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_235
timestamp -7200
transform 1 0 22172 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_247
timestamp -7200
transform 1 0 23276 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp -7200
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_253
timestamp -7200
transform 1 0 23828 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_258
timestamp -7200
transform 1 0 24288 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_270
timestamp -7200
transform 1 0 25392 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_282
timestamp -7200
transform 1 0 26496 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_288
timestamp -7200
transform 1 0 27048 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp -7200
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp -7200
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_43
timestamp -7200
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp -7200
transform 1 0 5428 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp -7200
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_69
timestamp -7200
transform 1 0 6900 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_75
timestamp -7200
transform 1 0 7452 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_88
timestamp -7200
transform 1 0 8648 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_100
timestamp -7200
transform 1 0 9752 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_135
timestamp -7200
transform 1 0 12972 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_143
timestamp -7200
transform 1 0 13708 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_162
timestamp -7200
transform 1 0 15456 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_169
timestamp -7200
transform 1 0 16100 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_184
timestamp -7200
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_201
timestamp -7200
transform 1 0 19044 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_213
timestamp -7200
transform 1 0 20148 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_221
timestamp -7200
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp -7200
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp -7200
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_249
timestamp -7200
transform 1 0 23460 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_260
timestamp -7200
transform 1 0 24472 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_269
timestamp -7200
transform 1 0 25300 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_277
timestamp -7200
transform 1 0 26036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_281
timestamp -7200
transform 1 0 26404 0 -1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp -7200
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp -7200
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp -7200
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp -7200
transform 1 0 3220 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_37
timestamp -7200
transform 1 0 3956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_63
timestamp -7200
transform 1 0 6348 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_69
timestamp -7200
transform 1 0 6900 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp -7200
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp -7200
transform 1 0 8372 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_102
timestamp -7200
transform 1 0 9936 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_119
timestamp -7200
transform 1 0 11500 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_125
timestamp -7200
transform 1 0 12052 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_134
timestamp -7200
transform 1 0 12880 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_154
timestamp -7200
transform 1 0 14720 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_167
timestamp -7200
transform 1 0 15916 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_173
timestamp -7200
transform 1 0 16468 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_190
timestamp -7200
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp -7200
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp -7200
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_209
timestamp -7200
transform 1 0 19780 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_213
timestamp -7200
transform 1 0 20148 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_232
timestamp -7200
transform 1 0 21896 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_244
timestamp -7200
transform 1 0 23000 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_285
timestamp -7200
transform 1 0 26772 0 1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp -7200
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp -7200
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_27
timestamp -7200
transform 1 0 3036 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_33
timestamp -7200
transform 1 0 3588 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_50
timestamp -7200
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_60
timestamp -7200
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_72
timestamp -7200
transform 1 0 7176 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_163
timestamp -7200
transform 1 0 15548 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp -7200
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_177
timestamp -7200
transform 1 0 16836 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_185
timestamp -7200
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_208
timestamp -7200
transform 1 0 19688 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp -7200
transform 1 0 20976 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_225
timestamp -7200
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_244
timestamp -7200
transform 1 0 23000 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_252
timestamp -7200
transform 1 0 23736 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_275
timestamp -7200
transform 1 0 25852 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp -7200
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_281
timestamp -7200
transform 1 0 26404 0 -1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp -7200
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp -7200
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp -7200
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp -7200
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_41
timestamp -7200
transform 1 0 4324 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_47
timestamp -7200
transform 1 0 4876 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_55
timestamp -7200
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_64
timestamp -7200
transform 1 0 6440 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp -7200
transform 1 0 8372 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_97
timestamp -7200
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp -7200
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp -7200
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp -7200
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp -7200
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_150
timestamp -7200
transform 1 0 14352 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_162
timestamp -7200
transform 1 0 15456 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_170
timestamp -7200
transform 1 0 16192 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_182
timestamp -7200
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_217
timestamp -7200
transform 1 0 20516 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_238
timestamp -7200
transform 1 0 22448 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_246
timestamp -7200
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_253
timestamp -7200
transform 1 0 23828 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_276
timestamp -7200
transform 1 0 25944 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_288
timestamp -7200
transform 1 0 27048 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp -7200
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_15
timestamp -7200
transform 1 0 1932 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_37
timestamp -7200
transform 1 0 3956 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp -7200
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_57
timestamp -7200
transform 1 0 5796 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_80
timestamp -7200
transform 1 0 7912 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_107
timestamp -7200
transform 1 0 10396 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp -7200
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_120
timestamp -7200
transform 1 0 11592 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_140
timestamp -7200
transform 1 0 13432 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_152
timestamp -7200
transform 1 0 14536 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_164
timestamp -7200
transform 1 0 15640 0 -1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp -7200
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_181
timestamp -7200
transform 1 0 17204 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_225
timestamp -7200
transform 1 0 21252 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_229
timestamp -7200
transform 1 0 21620 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_250
timestamp -7200
transform 1 0 23552 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp -7200
transform 1 0 26220 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp -7200
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_15
timestamp -7200
transform 1 0 1932 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_23
timestamp -7200
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp -7200
transform 1 0 3220 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_45
timestamp -7200
transform 1 0 4692 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_55
timestamp -7200
transform 1 0 5612 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp -7200
transform 1 0 7912 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_85
timestamp -7200
transform 1 0 8372 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_89
timestamp -7200
transform 1 0 8740 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_106
timestamp -7200
transform 1 0 10304 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_124
timestamp -7200
transform 1 0 11960 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_157
timestamp -7200
transform 1 0 14996 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_178
timestamp -7200
transform 1 0 16928 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_184
timestamp -7200
transform 1 0 17480 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_191
timestamp -7200
transform 1 0 18124 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp -7200
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_197
timestamp -7200
transform 1 0 18676 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_202
timestamp -7200
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_221
timestamp -7200
transform 1 0 20884 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_246
timestamp -7200
transform 1 0 23184 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_253
timestamp -7200
transform 1 0 23828 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_262
timestamp -7200
transform 1 0 24656 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_287
timestamp -7200
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp -7200
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_15
timestamp -7200
transform 1 0 1932 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_33
timestamp -7200
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_41
timestamp -7200
transform 1 0 4324 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp -7200
transform 1 0 5428 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_57
timestamp -7200
transform 1 0 5796 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_77
timestamp -7200
transform 1 0 7636 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_81
timestamp -7200
transform 1 0 8004 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_106
timestamp -7200
transform 1 0 10304 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_113
timestamp -7200
transform 1 0 10948 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp -7200
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_185
timestamp -7200
transform 1 0 17572 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_193
timestamp -7200
transform 1 0 18308 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_199
timestamp -7200
transform 1 0 18860 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_210
timestamp -7200
transform 1 0 19872 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_216
timestamp -7200
transform 1 0 20424 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_260
timestamp -7200
transform 1 0 24472 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_270
timestamp -7200
transform 1 0 25392 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_278
timestamp -7200
transform 1 0 26128 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_281
timestamp -7200
transform 1 0 26404 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp -7200
transform 1 0 828 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp -7200
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_48
timestamp -7200
transform 1 0 4968 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_52
timestamp -7200
transform 1 0 5336 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_69
timestamp -7200
transform 1 0 6900 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_78
timestamp -7200
transform 1 0 7728 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp -7200
transform 1 0 8372 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp -7200
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_109
timestamp -7200
transform 1 0 10580 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_125
timestamp -7200
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_136
timestamp -7200
transform 1 0 13064 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_149
timestamp -7200
transform 1 0 14260 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_161
timestamp -7200
transform 1 0 15364 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp -7200
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_241
timestamp -7200
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp -7200
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_276
timestamp -7200
transform 1 0 25944 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_288
timestamp -7200
transform 1 0 27048 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp -7200
transform 1 0 828 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_11
timestamp -7200
transform 1 0 1564 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_30
timestamp -7200
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_40
timestamp -7200
transform 1 0 4232 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_52
timestamp -7200
transform 1 0 5336 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_57
timestamp -7200
transform 1 0 5796 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_61
timestamp -7200
transform 1 0 6164 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_77
timestamp -7200
transform 1 0 7636 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_98
timestamp -7200
transform 1 0 9568 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp -7200
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp -7200
transform 1 0 10948 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_122
timestamp -7200
transform 1 0 11776 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_133
timestamp -7200
transform 1 0 12788 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_145
timestamp -7200
transform 1 0 13892 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_153
timestamp -7200
transform 1 0 14628 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_160
timestamp -7200
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_192
timestamp -7200
transform 1 0 18216 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_211
timestamp -7200
transform 1 0 19964 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp -7200
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_225
timestamp -7200
transform 1 0 21252 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_262
timestamp -7200
transform 1 0 24656 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_287
timestamp -7200
transform 1 0 26956 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp -7200
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp -7200
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp -7200
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_29
timestamp -7200
transform 1 0 3220 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_34
timestamp -7200
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_40
timestamp -7200
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_57
timestamp -7200
transform 1 0 5796 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_89
timestamp -7200
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_99
timestamp -7200
transform 1 0 9660 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_107
timestamp -7200
transform 1 0 10396 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_141
timestamp -7200
transform 1 0 13524 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_193
timestamp -7200
transform 1 0 18308 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_203
timestamp -7200
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_211
timestamp -7200
transform 1 0 19964 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_221
timestamp -7200
transform 1 0 20884 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_232
timestamp -7200
transform 1 0 21896 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_256
timestamp -7200
transform 1 0 24104 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_268
timestamp -7200
transform 1 0 25208 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_287
timestamp -7200
transform 1 0 26956 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp -7200
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_15
timestamp -7200
transform 1 0 1932 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_21
timestamp -7200
transform 1 0 2484 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp -7200
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_62
timestamp -7200
transform 1 0 6256 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_68
timestamp -7200
transform 1 0 6808 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_89
timestamp -7200
transform 1 0 8740 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp -7200
transform 1 0 10580 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_113
timestamp -7200
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_140
timestamp -7200
transform 1 0 13432 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_149
timestamp -7200
transform 1 0 14260 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_157
timestamp -7200
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_169
timestamp -7200
transform 1 0 16100 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_231
timestamp -7200
transform 1 0 21804 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_243
timestamp -7200
transform 1 0 22908 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_251
timestamp -7200
transform 1 0 23644 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp -7200
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp -7200
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp -7200
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_29
timestamp -7200
transform 1 0 3220 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_66
timestamp -7200
transform 1 0 6624 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp -7200
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp -7200
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_107
timestamp -7200
transform 1 0 10396 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp -7200
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_141
timestamp -7200
transform 1 0 13524 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_147
timestamp -7200
transform 1 0 14076 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_156
timestamp -7200
transform 1 0 14904 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_168
timestamp -7200
transform 1 0 16008 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_175
timestamp -7200
transform 1 0 16652 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_183
timestamp -7200
transform 1 0 17388 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp -7200
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_205
timestamp -7200
transform 1 0 19412 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_209
timestamp -7200
transform 1 0 19780 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_214
timestamp -7200
transform 1 0 20240 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_237
timestamp -7200
transform 1 0 22356 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp -7200
transform 1 0 23460 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_253
timestamp -7200
transform 1 0 23828 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_257
timestamp -7200
transform 1 0 24196 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_274
timestamp -7200
transform 1 0 25760 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_286
timestamp -7200
transform 1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp -7200
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_15
timestamp -7200
transform 1 0 1932 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_23
timestamp -7200
transform 1 0 2668 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_45
timestamp -7200
transform 1 0 4692 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_61
timestamp -7200
transform 1 0 6164 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_93
timestamp -7200
transform 1 0 9108 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_101
timestamp -7200
transform 1 0 9844 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp -7200
transform 1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_121
timestamp -7200
transform 1 0 11684 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp -7200
transform 1 0 15364 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp -7200
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp -7200
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_181
timestamp -7200
transform 1 0 17204 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_222
timestamp -7200
transform 1 0 20976 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_249
timestamp -7200
transform 1 0 23460 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_255
timestamp -7200
transform 1 0 24012 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp -7200
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp -7200
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp -7200
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_29
timestamp -7200
transform 1 0 3220 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_38
timestamp -7200
transform 1 0 4048 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_44
timestamp -7200
transform 1 0 4600 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_48
timestamp -7200
transform 1 0 4968 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_52
timestamp -7200
transform 1 0 5336 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_56
timestamp -7200
transform 1 0 5704 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_64
timestamp -7200
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_71
timestamp -7200
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_79
timestamp -7200
transform 1 0 7820 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp -7200
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp -7200
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_135
timestamp -7200
transform 1 0 12972 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp -7200
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_157
timestamp -7200
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_175
timestamp -7200
transform 1 0 16652 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp -7200
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_205
timestamp -7200
transform 1 0 19412 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_209
timestamp -7200
transform 1 0 19780 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_234
timestamp -7200
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp -7200
transform 1 0 23644 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_261
timestamp -7200
transform 1 0 24564 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_265
timestamp -7200
transform 1 0 24932 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_282
timestamp -7200
transform 1 0 26496 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_288
timestamp -7200
transform 1 0 27048 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp -7200
transform 1 0 828 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_11
timestamp -7200
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_44
timestamp -7200
transform 1 0 4600 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_50
timestamp -7200
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_133
timestamp -7200
transform 1 0 12788 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp -7200
transform 1 0 15364 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp -7200
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_201
timestamp -7200
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_219
timestamp -7200
transform 1 0 20700 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp -7200
transform 1 0 21068 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_261
timestamp -7200
transform 1 0 24564 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_3
timestamp -7200
transform 1 0 828 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_29
timestamp -7200
transform 1 0 3220 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_62
timestamp -7200
transform 1 0 6256 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_92
timestamp -7200
transform 1 0 9016 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_100
timestamp -7200
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_126
timestamp -7200
transform 1 0 12144 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_141
timestamp -7200
transform 1 0 13524 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_176
timestamp -7200
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp -7200
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_217
timestamp -7200
transform 1 0 20516 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp -7200
transform 1 0 23552 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_285
timestamp -7200
transform 1 0 26772 0 1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp -7200
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_15
timestamp -7200
transform 1 0 1932 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_48
timestamp -7200
transform 1 0 4968 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp -7200
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_65
timestamp -7200
transform 1 0 6532 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_72
timestamp -7200
transform 1 0 7176 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_80
timestamp -7200
transform 1 0 7912 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_98
timestamp -7200
transform 1 0 9568 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_104
timestamp -7200
transform 1 0 10120 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_113
timestamp -7200
transform 1 0 10948 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_139
timestamp -7200
transform 1 0 13340 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_145
timestamp -7200
transform 1 0 13892 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_162
timestamp -7200
transform 1 0 15456 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_181
timestamp -7200
transform 1 0 17204 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_208
timestamp -7200
transform 1 0 19688 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp -7200
transform 1 0 20976 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_260
timestamp -7200
transform 1 0 24472 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_277
timestamp -7200
transform 1 0 26036 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp -7200
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp -7200
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp -7200
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_46
timestamp -7200
transform 1 0 4784 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_59
timestamp -7200
transform 1 0 5980 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_70
timestamp -7200
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp -7200
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_107
timestamp -7200
transform 1 0 10396 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_115
timestamp -7200
transform 1 0 11132 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_134
timestamp -7200
transform 1 0 12880 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_157
timestamp -7200
transform 1 0 14996 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_174
timestamp -7200
transform 1 0 16560 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_217
timestamp -7200
transform 1 0 20516 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_269
timestamp -7200
transform 1 0 25300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_287
timestamp -7200
transform 1 0 26956 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_3
timestamp -7200
transform 1 0 828 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_11
timestamp -7200
transform 1 0 1564 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_40
timestamp -7200
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_48
timestamp -7200
transform 1 0 4968 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp -7200
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp -7200
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp -7200
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_86
timestamp -7200
transform 1 0 8464 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_103
timestamp -7200
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp -7200
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_113
timestamp -7200
transform 1 0 10948 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_125
timestamp -7200
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_135
timestamp -7200
transform 1 0 12972 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_143
timestamp -7200
transform 1 0 13708 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_181
timestamp -7200
transform 1 0 17204 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_187
timestamp -7200
transform 1 0 17756 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_220
timestamp -7200
transform 1 0 20792 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_249
timestamp -7200
transform 1 0 23460 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_277
timestamp -7200
transform 1 0 26036 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_3
timestamp -7200
transform 1 0 828 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_11
timestamp -7200
transform 1 0 1564 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp -7200
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_41
timestamp -7200
transform 1 0 4324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_48
timestamp -7200
transform 1 0 4968 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_69
timestamp -7200
transform 1 0 6900 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp -7200
transform 1 0 8004 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_85
timestamp -7200
transform 1 0 8372 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_95
timestamp -7200
transform 1 0 9292 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_112
timestamp -7200
transform 1 0 10856 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_124
timestamp -7200
transform 1 0 11960 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_136
timestamp -7200
transform 1 0 13064 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_148
timestamp -7200
transform 1 0 14168 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_221
timestamp -7200
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_247
timestamp -7200
transform 1 0 23276 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp -7200
transform 1 0 23644 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_253
timestamp -7200
transform 1 0 23828 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_259
timestamp -7200
transform 1 0 24380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_284
timestamp -7200
transform 1 0 26680 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_288
timestamp -7200
transform 1 0 27048 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp -7200
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp -7200
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_27
timestamp -7200
transform 1 0 3036 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_44
timestamp -7200
transform 1 0 4600 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp -7200
transform 1 0 5336 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_57
timestamp -7200
transform 1 0 5796 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_63
timestamp -7200
transform 1 0 6348 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_67
timestamp -7200
transform 1 0 6716 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_77
timestamp -7200
transform 1 0 7636 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_85
timestamp -7200
transform 1 0 8372 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_91
timestamp -7200
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_110
timestamp -7200
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp -7200
transform 1 0 10948 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_152
timestamp -7200
transform 1 0 14536 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_164
timestamp -7200
transform 1 0 15640 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_177
timestamp -7200
transform 1 0 16836 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp -7200
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_249
timestamp -7200
transform 1 0 23460 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_256
timestamp -7200
transform 1 0 24104 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_274
timestamp -7200
transform 1 0 25760 0 -1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp -7200
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp -7200
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp -7200
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp -7200
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp -7200
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_53
timestamp -7200
transform 1 0 5428 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_71
timestamp -7200
transform 1 0 7084 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp -7200
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_94
timestamp -7200
transform 1 0 9200 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_116
timestamp -7200
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp -7200
transform 1 0 13524 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_163
timestamp -7200
transform 1 0 15548 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_175
timestamp -7200
transform 1 0 16652 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_187
timestamp -7200
transform 1 0 17756 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp -7200
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_221
timestamp -7200
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_231
timestamp -7200
transform 1 0 21804 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_243
timestamp -7200
transform 1 0 22908 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp -7200
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_253
timestamp -7200
transform 1 0 23828 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_267
timestamp -7200
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_277
timestamp -7200
transform 1 0 26036 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_288
timestamp -7200
transform 1 0 27048 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp -7200
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp -7200
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp -7200
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_39
timestamp -7200
transform 1 0 4140 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_48
timestamp -7200
transform 1 0 4968 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_57
timestamp -7200
transform 1 0 5796 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_76
timestamp -7200
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_94
timestamp -7200
transform 1 0 9200 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp -7200
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_117
timestamp -7200
transform 1 0 11316 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_173
timestamp -7200
transform 1 0 16468 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_186
timestamp -7200
transform 1 0 17664 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_195
timestamp -7200
transform 1 0 18492 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_199
timestamp -7200
transform 1 0 18860 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp -7200
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_232
timestamp -7200
transform 1 0 21896 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_244
timestamp -7200
transform 1 0 23000 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_256
timestamp -7200
transform 1 0 24104 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp -7200
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_6
timestamp -7200
transform 1 0 1104 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_13
timestamp -7200
transform 1 0 1748 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_21
timestamp -7200
transform 1 0 2484 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp -7200
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_29
timestamp -7200
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_34
timestamp -7200
transform 1 0 3680 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_41
timestamp -7200
transform 1 0 4324 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_48
timestamp -7200
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_57
timestamp -7200
transform 1 0 5796 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_71
timestamp -7200
transform 1 0 7084 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp -7200
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_85
timestamp -7200
transform 1 0 8372 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_93
timestamp -7200
transform 1 0 9108 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_97
timestamp -7200
transform 1 0 9476 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_108
timestamp -7200
transform 1 0 10488 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_121
timestamp -7200
transform 1 0 11684 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_127
timestamp -7200
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_141
timestamp -7200
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_151
timestamp -7200
transform 1 0 14444 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_166
timestamp -7200
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_177
timestamp -7200
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_182
timestamp -7200
transform 1 0 17296 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_188
timestamp -7200
transform 1 0 17848 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_197
timestamp -7200
transform 1 0 18676 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_205
timestamp -7200
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_217
timestamp -7200
transform 1 0 20516 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_223
timestamp -7200
transform 1 0 21068 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_225
timestamp -7200
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_230
timestamp -7200
transform 1 0 21712 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_237
timestamp -7200
transform 1 0 22356 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_244
timestamp -7200
transform 1 0 23000 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp -7200
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_253
timestamp -7200
transform 1 0 23828 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_258
timestamp -7200
transform 1 0 24288 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_265
timestamp -7200
transform 1 0 24932 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_279
timestamp -7200
transform 1 0 26220 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_281
timestamp -7200
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_287
timestamp -7200
transform 1 0 26956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp -7200
transform -1 0 13340 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp -7200
transform -1 0 12972 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp -7200
transform 1 0 8372 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp -7200
transform -1 0 17204 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp -7200
transform 1 0 19412 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp -7200
transform -1 0 20056 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp -7200
transform -1 0 10764 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp -7200
transform 1 0 20148 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp -7200
transform -1 0 20148 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp -7200
transform -1 0 12972 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp -7200
transform -1 0 19412 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp -7200
transform -1 0 18400 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp -7200
transform -1 0 17848 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp -7200
transform -1 0 17112 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp -7200
transform -1 0 16744 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp -7200
transform 1 0 14720 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp -7200
transform -1 0 7820 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp -7200
transform -1 0 19412 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp -7200
transform -1 0 20148 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp -7200
transform -1 0 6348 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp -7200
transform 1 0 11224 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp -7200
transform -1 0 11776 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp -7200
transform -1 0 13064 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp -7200
transform -1 0 17572 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp -7200
transform -1 0 16836 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp -7200
transform 1 0 24564 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp -7200
transform -1 0 24564 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp -7200
transform -1 0 14904 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp -7200
transform 1 0 18676 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp -7200
transform 1 0 8372 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp -7200
transform -1 0 8280 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp -7200
transform 1 0 13708 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp -7200
transform -1 0 15272 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp -7200
transform 1 0 5888 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp -7200
transform -1 0 19504 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp -7200
transform -1 0 19412 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp -7200
transform 1 0 26404 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp -7200
transform -1 0 26312 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp -7200
transform -1 0 24564 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp -7200
transform -1 0 24564 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp -7200
transform -1 0 12880 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp -7200
transform -1 0 27140 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp -7200
transform 1 0 24380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp -7200
transform -1 0 7912 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp -7200
transform -1 0 7176 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp -7200
transform 1 0 22540 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp -7200
transform -1 0 22724 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp -7200
transform -1 0 26680 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp -7200
transform 1 0 23000 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp -7200
transform -1 0 25944 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp -7200
transform -1 0 25944 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp -7200
transform -1 0 27048 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp -7200
transform 1 0 6992 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp -7200
transform 1 0 10672 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp -7200
transform -1 0 25116 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp -7200
transform -1 0 27140 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp -7200
transform 1 0 22816 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp -7200
transform -1 0 22080 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp -7200
transform -1 0 22356 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp -7200
transform -1 0 5152 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp -7200
transform -1 0 14628 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp -7200
transform 1 0 13156 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp -7200
transform -1 0 26312 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp -7200
transform -1 0 25760 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp -7200
transform 1 0 3496 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp -7200
transform -1 0 13340 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp -7200
transform 1 0 8372 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp -7200
transform -1 0 21804 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp -7200
transform -1 0 21528 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp -7200
transform 1 0 21528 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp -7200
transform 1 0 21620 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp -7200
transform -1 0 21988 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp -7200
transform 1 0 19320 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp -7200
transform -1 0 19780 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp -7200
transform -1 0 27140 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp -7200
transform -1 0 18308 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp -7200
transform -1 0 11684 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp -7200
transform -1 0 23460 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp -7200
transform -1 0 3956 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp -7200
transform -1 0 26864 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp -7200
transform -1 0 27140 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp -7200
transform 1 0 16928 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp -7200
transform 1 0 16192 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp -7200
transform -1 0 23092 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp -7200
transform 1 0 10948 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp -7200
transform -1 0 25484 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp -7200
transform -1 0 4048 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp -7200
transform -1 0 3404 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp -7200
transform -1 0 4784 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp -7200
transform -1 0 14352 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp -7200
transform -1 0 8188 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp -7200
transform 1 0 8740 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp -7200
transform -1 0 4692 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp -7200
transform -1 0 3956 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp -7200
transform -1 0 14444 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp -7200
transform -1 0 8556 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp -7200
transform -1 0 24472 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp -7200
transform -1 0 16468 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp -7200
transform -1 0 15456 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp -7200
transform -1 0 22080 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp -7200
transform -1 0 4784 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp -7200
transform -1 0 23828 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp -7200
transform 1 0 22908 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp -7200
transform 1 0 22540 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp -7200
transform -1 0 18400 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp -7200
transform -1 0 10856 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp -7200
transform -1 0 22540 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp -7200
transform 1 0 9660 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp -7200
transform 1 0 26588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp -7200
transform -1 0 26220 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp -7200
transform 1 0 25944 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -7200
transform 1 0 24656 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp -7200
transform 1 0 24012 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp -7200
transform 1 0 23368 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp -7200
transform 1 0 22724 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp -7200
transform 1 0 22080 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp -7200
transform 1 0 21436 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp -7200
transform -1 0 20516 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp -7200
transform -1 0 17848 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input12
timestamp -7200
transform 1 0 16928 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp -7200
transform 1 0 16468 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_31
timestamp -7200
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -7200
transform -1 0 27416 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_32
timestamp -7200
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -7200
transform -1 0 27416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_33
timestamp -7200
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -7200
transform -1 0 27416 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_34
timestamp -7200
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -7200
transform -1 0 27416 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_35
timestamp -7200
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -7200
transform -1 0 27416 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_36
timestamp -7200
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -7200
transform -1 0 27416 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_37
timestamp -7200
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -7200
transform -1 0 27416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_38
timestamp -7200
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -7200
transform -1 0 27416 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_39
timestamp -7200
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -7200
transform -1 0 27416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_40
timestamp -7200
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -7200
transform -1 0 27416 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_41
timestamp -7200
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -7200
transform -1 0 27416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_42
timestamp -7200
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -7200
transform -1 0 27416 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_43
timestamp -7200
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -7200
transform -1 0 27416 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_44
timestamp -7200
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -7200
transform -1 0 27416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_45
timestamp -7200
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -7200
transform -1 0 27416 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_46
timestamp -7200
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -7200
transform -1 0 27416 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_47
timestamp -7200
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -7200
transform -1 0 27416 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_48
timestamp -7200
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -7200
transform -1 0 27416 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_49
timestamp -7200
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -7200
transform -1 0 27416 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_50
timestamp -7200
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -7200
transform -1 0 27416 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_51
timestamp -7200
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -7200
transform -1 0 27416 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_52
timestamp -7200
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -7200
transform -1 0 27416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_53
timestamp -7200
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -7200
transform -1 0 27416 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_54
timestamp -7200
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -7200
transform -1 0 27416 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_55
timestamp -7200
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -7200
transform -1 0 27416 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_56
timestamp -7200
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -7200
transform -1 0 27416 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_57
timestamp -7200
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -7200
transform -1 0 27416 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_58
timestamp -7200
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -7200
transform -1 0 27416 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_59
timestamp -7200
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -7200
transform -1 0 27416 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_60
timestamp -7200
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -7200
transform -1 0 27416 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_61
timestamp -7200
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -7200
transform -1 0 27416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp -7200
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp -7200
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp -7200
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp -7200
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp -7200
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp -7200
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68
timestamp -7200
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp -7200
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp -7200
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp -7200
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_72
timestamp -7200
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_73
timestamp -7200
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_74
timestamp -7200
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_75
timestamp -7200
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_76
timestamp -7200
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_77
timestamp -7200
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_78
timestamp -7200
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_79
timestamp -7200
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_80
timestamp -7200
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_81
timestamp -7200
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_82
timestamp -7200
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_83
timestamp -7200
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_84
timestamp -7200
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_85
timestamp -7200
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_86
timestamp -7200
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_87
timestamp -7200
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_88
timestamp -7200
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_89
timestamp -7200
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_90
timestamp -7200
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_91
timestamp -7200
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_92
timestamp -7200
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_93
timestamp -7200
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_94
timestamp -7200
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_95
timestamp -7200
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_96
timestamp -7200
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_97
timestamp -7200
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_98
timestamp -7200
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_99
timestamp -7200
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_100
timestamp -7200
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_101
timestamp -7200
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_102
timestamp -7200
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_103
timestamp -7200
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_104
timestamp -7200
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_105
timestamp -7200
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_106
timestamp -7200
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_107
timestamp -7200
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_108
timestamp -7200
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_109
timestamp -7200
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_110
timestamp -7200
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_111
timestamp -7200
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_112
timestamp -7200
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_113
timestamp -7200
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_114
timestamp -7200
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_115
timestamp -7200
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_116
timestamp -7200
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_117
timestamp -7200
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_118
timestamp -7200
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_119
timestamp -7200
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_120
timestamp -7200
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_121
timestamp -7200
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_122
timestamp -7200
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_123
timestamp -7200
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_124
timestamp -7200
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_125
timestamp -7200
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_126
timestamp -7200
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_127
timestamp -7200
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_128
timestamp -7200
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_129
timestamp -7200
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_130
timestamp -7200
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_131
timestamp -7200
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_132
timestamp -7200
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_133
timestamp -7200
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_134
timestamp -7200
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_135
timestamp -7200
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_136
timestamp -7200
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_137
timestamp -7200
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_138
timestamp -7200
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_139
timestamp -7200
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_140
timestamp -7200
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_141
timestamp -7200
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_142
timestamp -7200
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_143
timestamp -7200
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_144
timestamp -7200
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_145
timestamp -7200
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_146
timestamp -7200
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_147
timestamp -7200
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_148
timestamp -7200
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_149
timestamp -7200
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_150
timestamp -7200
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_151
timestamp -7200
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_152
timestamp -7200
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_153
timestamp -7200
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_154
timestamp -7200
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_155
timestamp -7200
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_156
timestamp -7200
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_157
timestamp -7200
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_158
timestamp -7200
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_159
timestamp -7200
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_160
timestamp -7200
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp -7200
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_162
timestamp -7200
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_163
timestamp -7200
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp -7200
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp -7200
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_166
timestamp -7200
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_167
timestamp -7200
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp -7200
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp -7200
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_170
timestamp -7200
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_171
timestamp -7200
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_172
timestamp -7200
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_173
timestamp -7200
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_174
timestamp -7200
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_175
timestamp -7200
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_176
timestamp -7200
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_177
timestamp -7200
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_178
timestamp -7200
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_179
timestamp -7200
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_180
timestamp -7200
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_181
timestamp -7200
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_182
timestamp -7200
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_183
timestamp -7200
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_184
timestamp -7200
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_185
timestamp -7200
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_186
timestamp -7200
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_187
timestamp -7200
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_188
timestamp -7200
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_189
timestamp -7200
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_190
timestamp -7200
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_191
timestamp -7200
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_192
timestamp -7200
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_193
timestamp -7200
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_194
timestamp -7200
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_195
timestamp -7200
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_196
timestamp -7200
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_197
timestamp -7200
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_198
timestamp -7200
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_199
timestamp -7200
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_200
timestamp -7200
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_201
timestamp -7200
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_202
timestamp -7200
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_203
timestamp -7200
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_204
timestamp -7200
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_205
timestamp -7200
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_206
timestamp -7200
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_207
timestamp -7200
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_208
timestamp -7200
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_209
timestamp -7200
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_210
timestamp -7200
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_211
timestamp -7200
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_212
timestamp -7200
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_213
timestamp -7200
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_214
timestamp -7200
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_215
timestamp -7200
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_216
timestamp -7200
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_217
timestamp -7200
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_218
timestamp -7200
transform 1 0 5704 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_219
timestamp -7200
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_220
timestamp -7200
transform 1 0 10856 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_221
timestamp -7200
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_222
timestamp -7200
transform 1 0 16008 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_223
timestamp -7200
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_224
timestamp -7200
transform 1 0 21160 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_225
timestamp -7200
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_226
timestamp -7200
transform 1 0 26312 0 1 16864
box -38 -48 130 592
<< labels >>
rlabel metal2 s 14064 16864 14064 16864 4 VGND
rlabel metal1 s 13984 17408 13984 17408 4 VPWR
rlabel metal1 s 4998 12682 4998 12682 4 _000_
rlabel metal2 s 3266 14246 3266 14246 4 _001_
rlabel metal1 s 8648 13498 8648 13498 4 _002_
rlabel metal1 s 8924 13498 8924 13498 4 _003_
rlabel metal1 s 4416 14586 4416 14586 4 _004_
rlabel metal2 s 2622 8194 2622 8194 4 _005_
rlabel metal1 s 3818 8602 3818 8602 4 _006_
rlabel metal2 s 2801 6834 2801 6834 4 _007_
rlabel metal1 s 5796 5882 5796 5882 4 _008_
rlabel metal1 s 7493 6154 7493 6154 4 _009_
rlabel metal1 s 8678 5066 8678 5066 4 _010_
rlabel metal1 s 11377 5066 11377 5066 4 _011_
rlabel metal1 s 20362 5066 20362 5066 4 _012_
rlabel metal1 s 18170 5338 18170 5338 4 _013_
rlabel metal2 s 19642 6596 19642 6596 4 _014_
rlabel metal2 s 22770 6018 22770 6018 4 _015_
rlabel metal1 s 23904 5066 23904 5066 4 _016_
rlabel metal1 s 25346 4794 25346 4794 4 _017_
rlabel metal1 s 24334 5746 24334 5746 4 _018_
rlabel metal2 s 24789 6834 24789 6834 4 _019_
rlabel metal2 s 25801 7310 25801 7310 4 _020_
rlabel metal1 s 21891 7310 21891 7310 4 _021_
rlabel metal1 s 23000 8942 23000 8942 4 _022_
rlabel metal1 s 24932 8058 24932 8058 4 _023_
rlabel metal2 s 21114 8092 21114 8092 4 _024_
rlabel metal2 s 18814 8194 18814 8194 4 _025_
rlabel metal1 s 16320 9010 16320 9010 4 _026_
rlabel metal1 s 16054 10030 16054 10030 4 _027_
rlabel metal2 s 3266 12750 3266 12750 4 _028_
rlabel metal2 s 6394 16422 6394 16422 4 _029_
rlabel metal1 s 3726 14586 3726 14586 4 _030_
rlabel metal1 s 2893 12682 2893 12682 4 _031_
rlabel metal1 s 13186 15606 13186 15606 4 _032_
rlabel metal1 s 12236 16218 12236 16218 4 _033_
rlabel metal1 s 15134 16218 15134 16218 4 _034_
rlabel metal1 s 9701 16694 9701 16694 4 _035_
rlabel metal1 s 8740 16218 8740 16218 4 _036_
rlabel metal1 s 11955 11594 11955 11594 4 _037_
rlabel metal1 s 8678 11594 8678 11594 4 _038_
rlabel metal1 s 9522 9690 9522 9690 4 _039_
rlabel metal1 s 9287 7922 9287 7922 4 _040_
rlabel metal1 s 8638 7310 8638 7310 4 _041_
rlabel metal2 s 15405 7242 15405 7242 4 _042_
rlabel metal1 s 16320 7922 16320 7922 4 _043_
rlabel metal2 s 12098 9282 12098 9282 4 _044_
rlabel metal2 s 13110 11764 13110 11764 4 _045_
rlabel metal1 s 16330 12682 16330 12682 4 _046_
rlabel metal1 s 18676 12410 18676 12410 4 _047_
rlabel metal2 s 19550 11798 19550 11798 4 _048_
rlabel metal1 s 25944 12886 25944 12886 4 _049_
rlabel metal1 s 23138 13940 23138 13940 4 _050_
rlabel metal1 s 25939 13838 25939 13838 4 _051_
rlabel metal1 s 25806 16660 25806 16660 4 _052_
rlabel metal1 s 24702 14586 24702 14586 4 _053_
rlabel metal2 s 22310 14212 22310 14212 4 _054_
rlabel metal1 s 21551 15674 21551 15674 4 _055_
rlabel metal2 s 20102 15300 20102 15300 4 _056_
rlabel metal2 s 18722 15334 18722 15334 4 _057_
rlabel metal2 s 15962 14756 15962 14756 4 _058_
rlabel metal2 s 13841 13838 13841 13838 4 _059_
rlabel metal2 s 11914 13940 11914 13940 4 _060_
rlabel metal2 s 11638 11458 11638 11458 4 _061_
rlabel metal2 s 7590 10812 7590 10812 4 _062_
rlabel metal1 s 7820 9554 7820 9554 4 _063_
rlabel metal1 s 6343 8398 6343 8398 4 _064_
rlabel metal1 s 6716 7378 6716 7378 4 _065_
rlabel metal1 s 11868 7514 11868 7514 4 _066_
rlabel metal1 s 14448 7310 14448 7310 4 _067_
rlabel metal2 s 12742 9520 12742 9520 4 _068_
rlabel metal2 s 12006 10370 12006 10370 4 _069_
rlabel metal1 s 13524 10234 13524 10234 4 _070_
rlabel metal1 s 18814 10642 18814 10642 4 _071_
rlabel metal2 s 22218 10948 22218 10948 4 _072_
rlabel metal1 s 23920 10778 23920 10778 4 _073_
rlabel metal1 s 25300 10642 25300 10642 4 _074_
rlabel metal1 s 26680 10098 26680 10098 4 _075_
rlabel metal1 s 27002 9996 27002 9996 4 _076_
rlabel metal1 s 25203 12342 25203 12342 4 _077_
rlabel metal2 s 21574 10982 21574 10982 4 _078_
rlabel metal1 s 21845 12682 21845 12682 4 _079_
rlabel metal1 s 20838 13498 20838 13498 4 _080_
rlabel metal1 s 19780 13498 19780 13498 4 _081_
rlabel metal2 s 19734 13770 19734 13770 4 _082_
rlabel metal2 s 16146 13634 16146 13634 4 _083_
rlabel metal1 s 14720 12410 14720 12410 4 _084_
rlabel metal1 s 3905 11254 3905 11254 4 _085_
rlabel metal1 s 9108 3162 9108 3162 4 _086_
rlabel metal1 s 6297 3638 6297 3638 4 _087_
rlabel metal1 s 6256 3162 6256 3162 4 _088_
rlabel metal2 s 3353 4658 3353 4658 4 _089_
rlabel metal2 s 4738 4930 4738 4930 4 _090_
rlabel metal1 s 9931 3570 9931 3570 4 _091_
rlabel metal1 s 11357 3638 11357 3638 4 _092_
rlabel metal2 s 12190 4454 12190 4454 4 _093_
rlabel metal2 s 2893 10098 2893 10098 4 _094_
rlabel metal1 s 8586 1802 8586 1802 4 _095_
rlabel metal1 s 6389 1462 6389 1462 4 _096_
rlabel metal2 s 4922 1666 4922 1666 4 _097_
rlabel metal2 s 2806 3842 2806 3842 4 _098_
rlabel metal1 s 3629 2890 3629 2890 4 _099_
rlabel metal1 s 9977 1462 9977 1462 4 _100_
rlabel metal2 s 12829 1462 12829 1462 4 _101_
rlabel metal1 s 11311 1462 11311 1462 4 _102_
rlabel metal2 s 15138 1462 15138 1462 4 _103_
rlabel metal1 s 17541 1462 17541 1462 4 _104_
rlabel metal2 s 17806 1870 17806 1870 4 _105_
rlabel metal1 s 18246 3638 18246 3638 4 _106_
rlabel metal1 s 20152 3978 20152 3978 4 _107_
rlabel metal2 s 20470 3366 20470 3366 4 _108_
rlabel metal1 s 18798 2890 18798 2890 4 _109_
rlabel metal2 s 16877 5134 16877 5134 4 _110_
rlabel metal1 s 16652 16626 16652 16626 4 _111_
rlabel metal2 s 18172 1394 18172 1394 4 _112_
rlabel metal1 s 5796 11866 5796 11866 4 _113_
rlabel metal2 s 20654 13107 20654 13107 4 _114_
rlabel metal1 s 4646 14518 4646 14518 4 _115_
rlabel metal1 s 4416 13498 4416 13498 4 _116_
rlabel metal1 s 4186 13361 4186 13361 4 _117_
rlabel metal1 s 6578 12070 6578 12070 4 _118_
rlabel metal1 s 4968 13498 4968 13498 4 _119_
rlabel metal2 s 13202 16235 13202 16235 4 _120_
rlabel metal2 s 10534 15776 10534 15776 4 _121_
rlabel metal2 s 9798 15436 9798 15436 4 _122_
rlabel metal2 s 5566 14722 5566 14722 4 _123_
rlabel metal2 s 3542 13634 3542 13634 4 _124_
rlabel metal1 s 5060 15130 5060 15130 4 _125_
rlabel metal1 s 9752 13838 9752 13838 4 _126_
rlabel metal2 s 9246 14076 9246 14076 4 _127_
rlabel metal1 s 6854 12682 6854 12682 4 _128_
rlabel metal1 s 7314 12750 7314 12750 4 _129_
rlabel metal2 s 10810 3978 10810 3978 4 _130_
rlabel metal1 s 14165 13362 14165 13362 4 _131_
rlabel metal2 s 13204 7310 13204 7310 4 _132_
rlabel metal1 s 8648 13430 8648 13430 4 _133_
rlabel metal1 s 8280 13362 8280 13362 4 _134_
rlabel metal2 s 4538 13770 4538 13770 4 _135_
rlabel metal2 s 4140 10098 4140 10098 4 _136_
rlabel metal1 s 4462 10098 4462 10098 4 _137_
rlabel metal1 s 15502 2550 15502 2550 4 _138_
rlabel metal2 s 16148 1870 16148 1870 4 _139_
rlabel metal1 s 13754 1360 13754 1360 4 _140_
rlabel metal1 s 14306 2414 14306 2414 4 _141_
rlabel metal2 s 15962 1921 15962 1921 4 _142_
rlabel metal2 s 17986 1462 17986 1462 4 _143_
rlabel metal1 s 19136 16762 19136 16762 4 _144_
rlabel metal1 s 20240 2482 20240 2482 4 _145_
rlabel metal1 s 20424 1394 20424 1394 4 _146_
rlabel metal1 s 20746 1870 20746 1870 4 _147_
rlabel metal1 s 19642 1870 19642 1870 4 _148_
rlabel metal1 s 20562 1428 20562 1428 4 _149_
rlabel metal1 s 14490 2618 14490 2618 4 _150_
rlabel metal1 s 15870 17034 15870 17034 4 _151_
rlabel metal1 s 16100 3706 16100 3706 4 _152_
rlabel metal1 s 15686 17102 15686 17102 4 _153_
rlabel metal2 s 15226 4692 15226 4692 4 _154_
rlabel metal2 s 13662 14756 13662 14756 4 _155_
rlabel metal1 s 14536 4794 14536 4794 4 _156_
rlabel metal2 s 13340 14620 13340 14620 4 _157_
rlabel metal1 s 14030 4794 14030 4794 4 _158_
rlabel metal1 s 12788 17102 12788 17102 4 _159_
rlabel metal1 s 12972 3706 12972 3706 4 _160_
rlabel metal3 s 12535 16660 12535 16660 4 _161_
rlabel metal1 s 13340 3162 13340 3162 4 _162_
rlabel metal1 s 13386 6766 13386 6766 4 _163_
rlabel metal1 s 12282 8398 12282 8398 4 _164_
rlabel metal1 s 13248 5338 13248 5338 4 _165_
rlabel metal2 s 11822 16626 11822 16626 4 _166_
rlabel metal1 s 14352 5134 14352 5134 4 _167_
rlabel metal1 s 6118 2482 6118 2482 4 _168_
rlabel metal2 s 2806 8262 2806 8262 4 _169_
rlabel metal1 s 2530 7956 2530 7956 4 _170_
rlabel metal1 s 3956 8534 3956 8534 4 _171_
rlabel metal2 s 18078 8993 18078 8993 4 _172_
rlabel metal2 s 4186 9010 4186 9010 4 _173_
rlabel metal1 s 3266 7310 3266 7310 4 _174_
rlabel metal1 s 2898 7344 2898 7344 4 _175_
rlabel metal2 s 5014 6868 5014 6868 4 _176_
rlabel metal2 s 5842 6834 5842 6834 4 _177_
rlabel metal2 s 6026 6460 6026 6460 4 _178_
rlabel metal1 s 9384 5814 9384 5814 4 _179_
rlabel metal2 s 18032 13396 18032 13396 4 _180_
rlabel metal2 s 7774 6052 7774 6052 4 _181_
rlabel metal1 s 10442 6698 10442 6698 4 _182_
rlabel metal1 s 8694 6256 8694 6256 4 _183_
rlabel metal1 s 20056 5746 20056 5746 4 _184_
rlabel metal1 s 11454 6188 11454 6188 4 _185_
rlabel metal1 s 20332 5882 20332 5882 4 _186_
rlabel metal1 s 20240 5134 20240 5134 4 _187_
rlabel metal1 s 19458 4080 19458 4080 4 _188_
rlabel metal1 s 18492 5882 18492 5882 4 _189_
rlabel metal2 s 18078 6834 18078 6834 4 _190_
rlabel metal1 s 18446 5168 18446 5168 4 _191_
rlabel metal1 s 18170 6188 18170 6188 4 _192_
rlabel metal1 s 20884 6902 20884 6902 4 _193_
rlabel metal1 s 20884 6630 20884 6630 4 _194_
rlabel metal1 s 22126 5848 22126 5848 4 _195_
rlabel metal1 s 20930 5678 20930 5678 4 _196_
rlabel metal1 s 24058 5542 24058 5542 4 _197_
rlabel metal1 s 23322 5100 23322 5100 4 _198_
rlabel metal1 s 24978 4454 24978 4454 4 _199_
rlabel metal1 s 25162 5814 25162 5814 4 _200_
rlabel metal1 s 25024 4658 25024 4658 4 _201_
rlabel metal2 s 24334 6426 24334 6426 4 _202_
rlabel metal2 s 24418 7242 24418 7242 4 _203_
rlabel metal1 s 23966 6426 23966 6426 4 _204_
rlabel metal2 s 19550 8466 19550 8466 4 _205_
rlabel metal2 s 23506 6868 23506 6868 4 _206_
rlabel metal1 s 25300 8602 25300 8602 4 _207_
rlabel metal1 s 23966 8568 23966 8568 4 _208_
rlabel metal1 s 25668 8398 25668 8398 4 _209_
rlabel metal1 s 21758 7854 21758 7854 4 _210_
rlabel metal2 s 22034 8160 22034 8160 4 _211_
rlabel metal1 s 23276 8398 23276 8398 4 _212_
rlabel metal1 s 23782 8976 23782 8976 4 _213_
rlabel metal1 s 23874 8466 23874 8466 4 _214_
rlabel metal1 s 24334 8058 24334 8058 4 _215_
rlabel metal1 s 23828 8262 23828 8262 4 _216_
rlabel metal2 s 24702 8075 24702 8075 4 _217_
rlabel metal1 s 20930 8024 20930 8024 4 _218_
rlabel metal2 s 20884 7990 20884 7990 4 _219_
rlabel metal1 s 17802 9044 17802 9044 4 _220_
rlabel metal1 s 18814 7854 18814 7854 4 _221_
rlabel metal2 s 18630 8092 18630 8092 4 _222_
rlabel metal1 s 16284 8602 16284 8602 4 _223_
rlabel metal1 s 15502 8874 15502 8874 4 _224_
rlabel metal1 s 17388 8942 17388 8942 4 _225_
rlabel metal1 s 3680 12274 3680 12274 4 _226_
rlabel metal2 s 6854 14722 6854 14722 4 _227_
rlabel metal2 s 6670 15844 6670 15844 4 _228_
rlabel metal1 s 11178 14586 11178 14586 4 _229_
rlabel metal1 s 6992 15674 6992 15674 4 _230_
rlabel metal3 s 4830 13413 4830 13413 4 _231_
rlabel metal1 s 4140 13498 4140 13498 4 _232_
rlabel metal1 s 7360 11594 7360 11594 4 _233_
rlabel metal1 s 19734 10166 19734 10166 4 _234_
rlabel metal1 s 3818 11866 3818 11866 4 _235_
rlabel metal1 s 4140 12070 4140 12070 4 _236_
rlabel metal1 s 13156 14926 13156 14926 4 _237_
rlabel metal2 s 6302 14144 6302 14144 4 _238_
rlabel metal2 s 5382 14756 5382 14756 4 _239_
rlabel metal1 s 5704 13974 5704 13974 4 _240_
rlabel metal2 s 5106 14382 5106 14382 4 _241_
rlabel metal1 s 6072 14926 6072 14926 4 _242_
rlabel metal2 s 6486 14688 6486 14688 4 _243_
rlabel metal1 s 9614 15572 9614 15572 4 _244_
rlabel metal1 s 13064 15130 13064 15130 4 _245_
rlabel metal1 s 12328 16014 12328 16014 4 _246_
rlabel metal1 s 11086 16082 11086 16082 4 _247_
rlabel metal3 s 12190 16133 12190 16133 4 _248_
rlabel metal1 s 13498 16014 13498 16014 4 _249_
rlabel metal1 s 14582 16048 14582 16048 4 _250_
rlabel metal2 s 10182 16014 10182 16014 4 _251_
rlabel metal1 s 10258 15912 10258 15912 4 _252_
rlabel metal1 s 10166 16218 10166 16218 4 _253_
rlabel metal1 s 10051 15538 10051 15538 4 _254_
rlabel metal1 s 8694 15572 8694 15572 4 _255_
rlabel metal2 s 8878 15844 8878 15844 4 _256_
rlabel metal1 s 14674 13260 14674 13260 4 _257_
rlabel metal1 s 13386 12784 13386 12784 4 _258_
rlabel metal1 s 11730 12784 11730 12784 4 _259_
rlabel metal1 s 6854 13906 6854 13906 4 _260_
rlabel metal1 s 14214 14518 14214 14518 4 _261_
rlabel metal1 s 10856 12342 10856 12342 4 _262_
rlabel metal2 s 15318 12852 15318 12852 4 _263_
rlabel metal2 s 9522 13226 9522 13226 4 _264_
rlabel metal1 s 9200 12614 9200 12614 4 _265_
rlabel metal2 s 8970 12444 8970 12444 4 _266_
rlabel metal1 s 19918 11152 19918 11152 4 _267_
rlabel metal2 s 8556 9010 8556 9010 4 _268_
rlabel metal2 s 9154 9690 9154 9690 4 _269_
rlabel metal1 s 8924 8398 8924 8398 4 _270_
rlabel metal2 s 8234 7412 8234 7412 4 _271_
rlabel metal2 s 13386 7650 13386 7650 4 _272_
rlabel metal1 s 15410 7990 15410 7990 4 _273_
rlabel metal2 s 12558 8738 12558 8738 4 _274_
rlabel metal1 s 12650 11220 12650 11220 4 _275_
rlabel metal1 s 15410 11322 15410 11322 4 _276_
rlabel metal2 s 18724 13362 18724 13362 4 _277_
rlabel metal1 s 18538 12240 18538 12240 4 _278_
rlabel metal3 s 20838 14909 20838 14909 4 _279_
rlabel metal1 s 19458 13158 19458 13158 4 _280_
rlabel metal1 s 20148 15538 20148 15538 4 _281_
rlabel metal1 s 15870 14246 15870 14246 4 _282_
rlabel metal1 s 18262 14824 18262 14824 4 _283_
rlabel metal1 s 25530 12784 25530 12784 4 _284_
rlabel metal1 s 25576 12954 25576 12954 4 _285_
rlabel metal1 s 25438 14586 25438 14586 4 _286_
rlabel metal1 s 26680 14586 26680 14586 4 _287_
rlabel metal2 s 24058 14756 24058 14756 4 _288_
rlabel metal2 s 22770 14586 22770 14586 4 _289_
rlabel metal1 s 21298 15572 21298 15572 4 _290_
rlabel metal1 s 20562 14416 20562 14416 4 _291_
rlabel metal1 s 19182 14892 19182 14892 4 _292_
rlabel metal1 s 15502 14416 15502 14416 4 _293_
rlabel metal1 s 13570 8364 13570 8364 4 _294_
rlabel metal1 s 14306 14484 14306 14484 4 _295_
rlabel metal1 s 12374 13294 12374 13294 4 _296_
rlabel metal1 s 7406 12614 7406 12614 4 _297_
rlabel metal1 s 11178 11152 11178 11152 4 _298_
rlabel metal2 s 15410 9758 15410 9758 4 _299_
rlabel metal1 s 6624 9690 6624 9690 4 _300_
rlabel metal1 s 6670 9146 6670 9146 4 _301_
rlabel metal1 s 7406 9044 7406 9044 4 _302_
rlabel metal1 s 8004 6698 8004 6698 4 _303_
rlabel metal1 s 11500 6970 11500 6970 4 _304_
rlabel metal2 s 13662 7922 13662 7922 4 _305_
rlabel metal1 s 13202 10030 13202 10030 4 _306_
rlabel metal1 s 20286 11152 20286 11152 4 _307_
rlabel metal1 s 12512 10098 12512 10098 4 _308_
rlabel metal1 s 17296 9418 17296 9418 4 _309_
rlabel metal1 s 14950 9996 14950 9996 4 _310_
rlabel metal1 s 17710 12682 17710 12682 4 _311_
rlabel metal1 s 18446 10234 18446 10234 4 _312_
rlabel metal2 s 20838 10948 20838 10948 4 _313_
rlabel metal1 s 23046 10234 23046 10234 4 _314_
rlabel metal1 s 24656 10234 24656 10234 4 _315_
rlabel metal1 s 24794 10166 24794 10166 4 _316_
rlabel metal2 s 26910 9588 26910 9588 4 _317_
rlabel metal1 s 24748 12750 24748 12750 4 _318_
rlabel metal1 s 21206 10234 21206 10234 4 _319_
rlabel metal1 s 21528 12614 21528 12614 4 _320_
rlabel metal1 s 21344 10030 21344 10030 4 _321_
rlabel metal1 s 15686 10064 15686 10064 4 _322_
rlabel metal1 s 20240 9622 20240 9622 4 _323_
rlabel metal1 s 19274 13294 19274 13294 4 _324_
rlabel metal1 s 18262 9622 18262 9622 4 _325_
rlabel metal2 s 16606 12070 16606 12070 4 _326_
rlabel metal2 s 15226 10778 15226 10778 4 _327_
rlabel metal1 s 5244 9622 5244 9622 4 _328_
rlabel metal1 s 5428 9486 5428 9486 4 _329_
rlabel metal1 s 5796 11186 5796 11186 4 _330_
rlabel metal1 s 4646 11152 4646 11152 4 _331_
rlabel metal1 s 4416 9894 4416 9894 4 _332_
rlabel metal1 s 4738 9520 4738 9520 4 _333_
rlabel metal1 s 13754 4114 13754 4114 4 _334_
rlabel metal2 s 9614 3434 9614 3434 4 _335_
rlabel metal1 s 6900 4046 6900 4046 4 _336_
rlabel metal1 s 7176 2958 7176 2958 4 _337_
rlabel metal1 s 6900 5338 6900 5338 4 _338_
rlabel metal2 s 5198 4930 5198 4930 4 _339_
rlabel metal2 s 12374 4131 12374 4131 4 _340_
rlabel metal2 s 10994 4250 10994 4250 4 _341_
rlabel metal2 s 11730 4794 11730 4794 4 _342_
rlabel metal1 s 4232 9486 4232 9486 4 _343_
rlabel metal3 s 9338 3077 9338 3077 4 _344_
rlabel metal1 s 9292 2482 9292 2482 4 _345_
rlabel metal2 s 14490 2108 14490 2108 4 _346_
rlabel metal2 s 6394 2074 6394 2074 4 _347_
rlabel metal1 s 6716 1870 6716 1870 4 _348_
rlabel metal2 s 5198 2652 5198 2652 4 _349_
rlabel metal2 s 5106 1836 5106 1836 4 _350_
rlabel metal1 s 3634 4012 3634 4012 4 _351_
rlabel metal1 s 3220 3570 3220 3570 4 _352_
rlabel metal2 s 4002 3740 4002 3740 4 _353_
rlabel metal1 s 3772 2482 3772 2482 4 _354_
rlabel metal1 s 12466 3570 12466 3570 4 _355_
rlabel metal1 s 10626 2822 10626 2822 4 _356_
rlabel metal1 s 10396 1870 10396 1870 4 _357_
rlabel metal2 s 12466 2822 12466 2822 4 _358_
rlabel metal1 s 12696 1870 12696 1870 4 _359_
rlabel metal1 s 11642 2482 11642 2482 4 _360_
rlabel metal2 s 11546 2074 11546 2074 4 _361_
rlabel metal1 s 14674 1904 14674 1904 4 _362_
rlabel metal1 s 14904 1870 14904 1870 4 _363_
rlabel metal1 s 17020 2822 17020 2822 4 _364_
rlabel metal1 s 17204 2482 17204 2482 4 _365_
rlabel metal1 s 16468 2822 16468 2822 4 _366_
rlabel metal1 s 17526 2516 17526 2516 4 _367_
rlabel metal1 s 17480 4046 17480 4046 4 _368_
rlabel metal1 s 17802 4046 17802 4046 4 _369_
rlabel metal1 s 18814 4590 18814 4590 4 _370_
rlabel metal2 s 19366 4250 19366 4250 4 _371_
rlabel metal1 s 18906 4012 18906 4012 4 _372_
rlabel metal1 s 19872 2958 19872 2958 4 _373_
rlabel metal1 s 17710 3570 17710 3570 4 _374_
rlabel metal2 s 18354 3162 18354 3162 4 _375_
rlabel metal1 s 16100 5746 16100 5746 4 _376_
rlabel metal1 s 16560 5746 16560 5746 4 _377_
rlabel metal3 s 16054 9435 16054 9435 4 clk
rlabel metal3 s 14306 9571 14306 9571 4 clknet_0_clk
rlabel metal1 s 2070 6834 2070 6834 4 clknet_3_0__leaf_clk
rlabel metal1 s 12558 1258 12558 1258 4 clknet_3_1__leaf_clk
rlabel metal2 s 2714 11798 2714 11798 4 clknet_3_2__leaf_clk
rlabel metal2 s 8602 15538 8602 15538 4 clknet_3_3__leaf_clk
rlabel metal1 s 17710 1258 17710 1258 4 clknet_3_4__leaf_clk
rlabel metal2 s 21022 3842 21022 3842 4 clknet_3_5__leaf_clk
rlabel metal1 s 19918 12886 19918 12886 4 clknet_3_6__leaf_clk
rlabel metal2 s 21298 11458 21298 11458 4 clknet_3_7__leaf_clk
rlabel metal1 s 14490 12172 14490 12172 4 net1
rlabel metal2 s 20378 15181 20378 15181 4 net10
rlabel metal1 s 10074 17068 10074 17068 4 net100
rlabel metal2 s 22402 10778 22402 10778 4 net101
rlabel metal2 s 3450 14076 3450 14076 4 net102
rlabel metal2 s 25254 10268 25254 10268 4 net103
rlabel metal2 s 25801 9486 25801 9486 4 net104
rlabel metal1 s 17848 8942 17848 8942 4 net105
rlabel metal1 s 17070 9486 17070 9486 4 net106
rlabel metal1 s 21850 7888 21850 7888 4 net107
rlabel metal1 s 11500 5882 11500 5882 4 net108
rlabel metal2 s 23690 6732 23690 6732 4 net109
rlabel metal2 s 16468 12852 16468 12852 4 net11
rlabel metal1 s 3450 12274 3450 12274 4 net110
rlabel metal2 s 2065 12274 2065 12274 4 net111
rlabel metal1 s 4140 12954 4140 12954 4 net112
rlabel metal1 s 13202 15538 13202 15538 4 net113
rlabel metal1 s 7314 15537 7314 15537 4 net114
rlabel metal1 s 9752 6426 9752 6426 4 net115
rlabel metal1 s 4140 7514 4140 7514 4 net116
rlabel metal2 s 3542 8092 3542 8092 4 net117
rlabel metal2 s 12558 16490 12558 16490 4 net118
rlabel metal1 s 7682 5746 7682 5746 4 net119
rlabel metal1 s 17112 16966 17112 16966 4 net12
rlabel metal2 s 23782 4964 23782 4964 4 net120
rlabel metal2 s 14858 8092 14858 8092 4 net121
rlabel metal2 s 14766 16490 14766 16490 4 net122
rlabel metal2 s 21390 6052 21390 6052 4 net123
rlabel metal2 s 4370 10234 4370 10234 4 net124
rlabel metal2 s 23138 7514 23138 7514 4 net125
rlabel metal1 s 23644 8602 23644 8602 4 net126
rlabel metal2 s 23230 9282 23230 9282 4 net127
rlabel metal2 s 17710 10336 17710 10336 4 net128
rlabel metal2 s 10148 12750 10148 12750 4 net129
rlabel metal1 s 7222 10132 7222 10132 4 net13
rlabel metal1 s 21758 9146 21758 9146 4 net130
rlabel metal2 s 10350 6834 10350 6834 4 net131
rlabel metal1 s 3864 17306 3864 17306 4 net14
rlabel metal2 s 1518 17527 1518 17527 4 net15
rlabel metal2 s 874 17527 874 17527 4 net16
rlabel metal1 s 9200 17306 9200 17306 4 net17
rlabel metal1 s 6716 17306 6716 17306 4 net18
rlabel metal1 s 5796 17306 5796 17306 4 net19
rlabel metal1 s 25714 16422 25714 16422 4 net2
rlabel metal1 s 5336 17170 5336 17170 4 net20
rlabel metal2 s 4738 17459 4738 17459 4 net21
rlabel metal2 s 3450 17459 3450 17459 4 net22
rlabel metal2 s 2714 17452 2714 17452 4 net23
rlabel metal2 s 12190 13906 12190 13906 4 net24
rlabel metal1 s 12001 13838 12001 13838 4 net25
rlabel metal1 s 9246 2958 9246 2958 4 net26
rlabel metal1 s 16468 14586 16468 14586 4 net27
rlabel metal1 s 19734 14790 19734 14790 4 net28
rlabel metal1 s 18763 14450 18763 14450 4 net29
rlabel metal1 s 17526 16490 17526 16490 4 net3
rlabel metal1 s 10258 4658 10258 4658 4 net30
rlabel metal1 s 20745 14926 20745 14926 4 net31
rlabel metal1 s 19315 15606 19315 15606 4 net32
rlabel metal1 s 11339 4046 11339 4046 4 net33
rlabel metal2 s 18428 13362 18428 13362 4 net34
rlabel metal1 s 17475 11662 17475 11662 4 net35
rlabel metal1 s 16422 14790 16422 14790 4 net36
rlabel metal1 s 15221 14858 15221 14858 4 net37
rlabel metal2 s 14881 12274 14881 12274 4 net38
rlabel metal1 s 15052 12750 15052 12750 4 net39
rlabel metal2 s 18170 16354 18170 16354 4 net4
rlabel metal1 s 6670 4012 6670 4012 4 net40
rlabel metal1 s 17894 13328 17894 13328 4 net41
rlabel metal1 s 17705 13770 17705 13770 4 net42
rlabel metal1 s 5014 4692 5014 4692 4 net43
rlabel metal1 s 13018 10064 13018 10064 4 net44
rlabel metal1 s 11132 9146 11132 9146 4 net45
rlabel metal1 s 13110 7344 13110 7344 4 net46
rlabel metal1 s 16100 12750 16100 12750 4 net47
rlabel metal1 s 15819 11594 15819 11594 4 net48
rlabel metal2 s 25714 13226 25714 13226 4 net49
rlabel metal1 s 19274 16456 19274 16456 4 net5
rlabel metal1 s 23593 13362 23593 13362 4 net50
rlabel metal2 s 13836 10098 13836 10098 4 net51
rlabel metal1 s 18998 14960 18998 14960 4 net52
rlabel metal1 s 8694 10438 8694 10438 4 net53
rlabel metal2 s 7590 9894 7590 9894 4 net54
rlabel metal1 s 14168 8398 14168 8398 4 net55
rlabel metal1 s 14122 14416 14122 14416 4 net56
rlabel metal1 s 6762 2958 6762 2958 4 net57
rlabel metal2 s 18078 10778 18078 10778 4 net58
rlabel metal1 s 18676 10778 18676 10778 4 net59
rlabel metal1 s 20010 17272 20010 17272 4 net6
rlabel metal2 s 26312 13396 26312 13396 4 net60
rlabel metal2 s 25622 10914 25622 10914 4 net61
rlabel metal1 s 23322 10574 23322 10574 4 net62
rlabel metal1 s 23179 11594 23179 11594 4 net63
rlabel metal2 s 11914 4522 11914 4522 4 net64
rlabel metal1 s 26312 6834 26312 6834 4 net65
rlabel metal1 s 24932 5882 24932 5882 4 net66
rlabel metal1 s 7360 7174 7360 7174 4 net67
rlabel metal2 s 6486 7718 6486 7718 4 net68
rlabel metal2 s 23248 14450 23248 14450 4 net69
rlabel metal2 s 22770 16728 22770 16728 4 net7
rlabel metal2 s 22034 14620 22034 14620 4 net70
rlabel metal1 s 24886 14416 24886 14416 4 net71
rlabel metal2 s 24881 13430 24881 13430 4 net72
rlabel metal2 s 24886 16796 24886 16796 4 net73
rlabel metal1 s 24927 15606 24927 15606 4 net74
rlabel metal1 s 26036 16014 26036 16014 4 net75
rlabel metal1 s 7222 8976 7222 8976 4 net76
rlabel metal2 s 11362 11900 11362 11900 4 net77
rlabel metal1 s 24334 14450 24334 14450 4 net78
rlabel metal1 s 25729 14858 25729 14858 4 net79
rlabel metal1 s 20010 16524 20010 16524 4 net8
rlabel metal1 s 23276 12954 23276 12954 4 net80
rlabel metal1 s 19504 12954 19504 12954 4 net81
rlabel metal2 s 21666 11186 21666 11186 4 net82
rlabel metal1 s 4002 5712 4002 5712 4 net83
rlabel metal2 s 12834 11662 12834 11662 4 net84
rlabel metal2 s 13841 11662 13841 11662 4 net85
rlabel metal1 s 24932 10574 24932 10574 4 net86
rlabel metal1 s 25024 10778 25024 10778 4 net87
rlabel metal2 s 4462 8636 4462 8636 4 net88
rlabel metal2 s 12282 10302 12282 10302 4 net89
rlabel metal1 s 21022 16490 21022 16490 4 net9
rlabel metal2 s 8694 11186 8694 11186 4 net90
rlabel metal1 s 20930 15538 20930 15538 4 net91
rlabel metal1 s 20286 13396 20286 13396 4 net92
rlabel metal1 s 22314 13430 22314 13430 4 net93
rlabel metal1 s 22448 7922 22448 7922 4 net94
rlabel metal2 s 19826 11764 19826 11764 4 net95
rlabel metal1 s 20194 6834 20194 6834 4 net96
rlabel metal1 s 18487 6834 18487 6834 4 net97
rlabel metal2 s 24978 12954 24978 12954 4 net98
rlabel metal2 s 16790 8874 16790 8874 4 net99
rlabel metal2 s 874 908 874 908 4 o_digital[0]
rlabel metal2 s 18354 772 18354 772 4 o_digital[10]
rlabel metal2 s 20102 772 20102 772 4 o_digital[11]
rlabel metal2 s 21850 1384 21850 1384 4 o_digital[12]
rlabel metal2 s 23598 874 23598 874 4 o_digital[13]
rlabel metal2 s 25346 1044 25346 1044 4 o_digital[14]
rlabel metal2 s 27094 1078 27094 1078 4 o_digital[15]
rlabel metal2 s 2622 534 2622 534 4 o_digital[1]
rlabel metal2 s 4370 1044 4370 1044 4 o_digital[2]
rlabel metal2 s 6118 1384 6118 1384 4 o_digital[3]
rlabel metal2 s 7866 636 7866 636 4 o_digital[4]
rlabel metal2 s 9614 636 9614 636 4 o_digital[5]
rlabel metal2 s 11362 636 11362 636 4 o_digital[6]
rlabel metal2 s 13110 636 13110 636 4 o_digital[7]
rlabel metal2 s 14858 636 14858 636 4 o_digital[8]
rlabel metal2 s 16606 1180 16606 1180 4 o_digital[9]
rlabel metal1 s 26588 17102 26588 17102 4 rst_n
rlabel metal1 s 26036 16626 26036 16626 4 ui_in[0]
rlabel metal1 s 26174 17136 26174 17136 4 ui_in[1]
rlabel metal1 s 24748 17102 24748 17102 4 ui_in[2]
rlabel metal1 s 24012 17102 24012 17102 4 ui_in[3]
rlabel metal1 s 23460 17102 23460 17102 4 ui_in[4]
rlabel metal1 s 22816 17102 22816 17102 4 ui_in[5]
rlabel metal2 s 22034 17418 22034 17418 4 ui_in[6]
rlabel metal2 s 21666 17425 21666 17425 4 ui_in[7]
rlabel metal1 s 19964 17102 19964 17102 4 uio_in[2]
rlabel metal2 s 17802 17306 17802 17306 4 uio_in[5]
rlabel metal1 s 16928 17102 16928 17102 4 uio_in[6]
rlabel metal1 s 16376 17102 16376 17102 4 uio_in[7]
rlabel metal2 s 2070 17112 2070 17112 4 uio_oe[5]
rlabel metal1 s 5106 16626 5106 16626 4 uio_out[0]
rlabel metal1 s 9246 16150 9246 16150 4 uio_out[1]
rlabel metal1 s 7406 17170 7406 17170 4 uio_out[3]
rlabel metal1 s 7130 10778 7130 10778 4 uio_out[4]
rlabel metal1 s 6946 17238 6946 17238 4 uio_out[5]
rlabel metal1 s 15962 17306 15962 17306 4 uo_out[0]
rlabel metal1 s 15318 17238 15318 17238 4 uo_out[1]
rlabel metal1 s 13754 17306 13754 17306 4 uo_out[2]
rlabel metal1 s 13248 17238 13248 17238 4 uo_out[3]
rlabel metal1 s 12742 17306 12742 17306 4 uo_out[4]
rlabel metal2 s 12374 17248 12374 17248 4 uo_out[5]
rlabel metal1 s 11960 16762 11960 16762 4 uo_out[6]
rlabel metal1 s 11822 16558 11822 16558 4 uo_out[7]
rlabel metal2 s 5198 11764 5198 11764 4 wrapped.o_busy
rlabel metal2 s 8050 16252 8050 16252 4 wrapped.o_copi
rlabel metal2 s 4646 14722 4646 14722 4 wrapped.o_cs_n
rlabel metal1 s 12834 11798 12834 11798 4 wrapped.o_data\[0\]
rlabel metal2 s 8510 4896 8510 4896 4 wrapped.o_data\[1\]
rlabel metal2 s 15134 7123 15134 7123 4 wrapped.o_data\[2\]
rlabel metal2 s 8712 6834 8712 6834 4 wrapped.o_data\[3\]
rlabel metal1 s 8372 7922 8372 7922 4 wrapped.o_data\[4\]
rlabel metal1 s 15456 3910 15456 3910 4 wrapped.o_data\[5\]
rlabel metal1 s 17664 7718 17664 7718 4 wrapped.o_data\[6\]
rlabel metal2 s 13293 12750 13293 12750 4 wrapped.o_data\[7\]
rlabel metal1 s 3542 12750 3542 12750 4 wrapped.o_data_valid
rlabel metal1 s 9706 2074 9706 2074 4 wrapped.o_digital$17\[0\]
rlabel metal1 s 17296 1734 17296 1734 4 wrapped.o_digital$17\[10\]
rlabel metal2 s 19366 1411 19366 1411 4 wrapped.o_digital$17\[11\]
rlabel metal2 s 19642 4522 19642 4522 4 wrapped.o_digital$17\[12\]
rlabel metal1 s 19964 1394 19964 1394 4 wrapped.o_digital$17\[13\]
rlabel metal2 s 20424 3026 20424 3026 4 wrapped.o_digital$17\[14\]
rlabel metal1 s 18584 4998 18584 4998 4 wrapped.o_digital$17\[15\]
rlabel metal1 s 7084 2482 7084 2482 4 wrapped.o_digital$17\[1\]
rlabel metal2 s 15686 2788 15686 2788 4 wrapped.o_digital$17\[2\]
rlabel metal2 s 14398 4318 14398 4318 4 wrapped.o_digital$17\[3\]
rlabel metal2 s 14306 4097 14306 4097 4 wrapped.o_digital$17\[4\]
rlabel metal1 s 11408 2958 11408 2958 4 wrapped.o_digital$17\[5\]
rlabel metal1 s 14076 1530 14076 1530 4 wrapped.o_digital$17\[6\]
rlabel metal1 s 12834 816 12834 816 4 wrapped.o_digital$17\[7\]
rlabel metal1 s 14214 1190 14214 1190 4 wrapped.o_digital$17\[8\]
rlabel metal1 s 16376 1530 16376 1530 4 wrapped.o_digital$17\[9\]
rlabel metal2 s 6026 16082 6026 16082 4 wrapped.o_sclk
rlabel metal2 s 19366 8738 19366 8738 4 wrapped.o_spi_address\[10\]
rlabel metal1 s 21114 6902 21114 6902 4 wrapped.o_spi_address\[11\]
rlabel metal1 s 23966 10234 23966 10234 4 wrapped.o_spi_address\[12\]
rlabel metal2 s 25162 8908 25162 8908 4 wrapped.o_spi_address\[13\]
rlabel metal2 s 25254 8806 25254 8806 4 wrapped.o_spi_address\[14\]
rlabel metal2 s 25898 8024 25898 8024 4 wrapped.o_spi_address\[15\]
rlabel metal1 s 25254 8398 25254 8398 4 wrapped.o_spi_address\[16\]
rlabel metal2 s 21482 9180 21482 9180 4 wrapped.o_spi_address\[17\]
rlabel metal1 s 21482 9486 21482 9486 4 wrapped.o_spi_address\[18\]
rlabel metal1 s 21666 9486 21666 9486 4 wrapped.o_spi_address\[19\]
rlabel metal1 s 4876 8398 4876 8398 4 wrapped.o_spi_address\[1\]
rlabel metal2 s 21758 8942 21758 8942 4 wrapped.o_spi_address\[20\]
rlabel metal1 s 19688 9078 19688 9078 4 wrapped.o_spi_address\[21\]
rlabel metal2 s 18262 9792 18262 9792 4 wrapped.o_spi_address\[22\]
rlabel metal1 s 16238 9690 16238 9690 4 wrapped.o_spi_address\[23\]
rlabel metal2 s 4922 8704 4922 8704 4 wrapped.o_spi_address\[2\]
rlabel metal1 s 6900 6222 6900 6222 4 wrapped.o_spi_address\[3\]
rlabel metal1 s 7314 6630 7314 6630 4 wrapped.o_spi_address\[4\]
rlabel metal1 s 10810 6154 10810 6154 4 wrapped.o_spi_address\[5\]
rlabel metal1 s 9292 6222 9292 6222 4 wrapped.o_spi_address\[6\]
rlabel metal1 s 10718 6222 10718 6222 4 wrapped.o_spi_address\[7\]
rlabel metal2 s 20930 6919 20930 6919 4 wrapped.o_spi_address\[8\]
rlabel metal1 s 20010 6868 20010 6868 4 wrapped.o_spi_address\[9\]
rlabel metal2 s 7958 3162 7958 3162 4 wrapped.player.buffer\[0\]
rlabel metal1 s 7084 2618 7084 2618 4 wrapped.player.buffer\[1\]
rlabel metal1 s 5566 2958 5566 2958 4 wrapped.player.buffer\[2\]
rlabel metal1 s 4508 4794 4508 4794 4 wrapped.player.buffer\[3\]
rlabel metal2 s 5566 4624 5566 4624 4 wrapped.player.buffer\[4\]
rlabel metal1 s 10764 3706 10764 3706 4 wrapped.player.buffer\[5\]
rlabel metal1 s 12328 3706 12328 3706 4 wrapped.player.buffer\[6\]
rlabel metal1 s 12696 5134 12696 5134 4 wrapped.player.buffer\[7\]
rlabel metal2 s 4646 10404 4646 10404 4 wrapped.player.received_samples
rlabel metal1 s 10488 12206 10488 12206 4 wrapped.spi_flash.address\[0\]
rlabel metal1 s 18354 11322 18354 11322 4 wrapped.spi_flash.address\[10\]
rlabel metal1 s 20930 11662 20930 11662 4 wrapped.spi_flash.address\[11\]
rlabel metal1 s 24426 12648 24426 12648 4 wrapped.spi_flash.address\[12\]
rlabel metal2 s 26266 11339 26266 11339 4 wrapped.spi_flash.address\[13\]
rlabel metal2 s 26450 12036 26450 12036 4 wrapped.spi_flash.address\[14\]
rlabel metal1 s 26864 9690 26864 9690 4 wrapped.spi_flash.address\[15\]
rlabel metal2 s 27094 15028 27094 15028 4 wrapped.spi_flash.address\[16\]
rlabel metal1 s 22862 15606 22862 15606 4 wrapped.spi_flash.address\[17\]
rlabel metal1 s 22862 12852 22862 12852 4 wrapped.spi_flash.address\[18\]
rlabel metal1 s 21482 13940 21482 13940 4 wrapped.spi_flash.address\[19\]
rlabel metal1 s 8418 11084 8418 11084 4 wrapped.spi_flash.address\[1\]
rlabel metal1 s 19412 14586 19412 14586 4 wrapped.spi_flash.address\[20\]
rlabel metal1 s 18354 13974 18354 13974 4 wrapped.spi_flash.address\[21\]
rlabel metal2 s 16514 14212 16514 14212 4 wrapped.spi_flash.address\[22\]
rlabel metal1 s 13846 12648 13846 12648 4 wrapped.spi_flash.address\[23\]
rlabel metal2 s 8694 10404 8694 10404 4 wrapped.spi_flash.address\[2\]
rlabel metal1 s 7038 8500 7038 8500 4 wrapped.spi_flash.address\[3\]
rlabel metal2 s 7774 7548 7774 7548 4 wrapped.spi_flash.address\[4\]
rlabel metal2 s 12926 8228 12926 8228 4 wrapped.spi_flash.address\[5\]
rlabel metal1 s 13662 7514 13662 7514 4 wrapped.spi_flash.address\[6\]
rlabel metal1 s 10764 9622 10764 9622 4 wrapped.spi_flash.address\[7\]
rlabel metal1 s 13110 10642 13110 10642 4 wrapped.spi_flash.address\[8\]
rlabel metal1 s 14950 11186 14950 11186 4 wrapped.spi_flash.address\[9\]
rlabel metal1 s 6716 12818 6716 12818 4 wrapped.spi_flash.fsm_state\[0\]
rlabel metal1 s 10212 13838 10212 13838 4 wrapped.spi_flash.fsm_state\[1\]
rlabel metal2 s 8234 14552 8234 14552 4 wrapped.spi_flash.fsm_state\[2\]
rlabel metal1 s 9706 14960 9706 14960 4 wrapped.spi_flash.fsm_state\[3\]
rlabel metal2 s 3818 14620 3818 14620 4 wrapped.spi_flash.fsm_state\[4\]
rlabel metal1 s 19274 11764 19274 11764 4 wrapped.spi_flash.shift_reg\[10\]
rlabel metal1 s 21850 12172 21850 12172 4 wrapped.spi_flash.shift_reg\[11\]
rlabel metal1 s 24518 13498 24518 13498 4 wrapped.spi_flash.shift_reg\[12\]
rlabel metal2 s 25990 14212 25990 14212 4 wrapped.spi_flash.shift_reg\[13\]
rlabel metal2 s 26616 14450 26616 14450 4 wrapped.spi_flash.shift_reg\[14\]
rlabel metal2 s 25806 16388 25806 16388 4 wrapped.spi_flash.shift_reg\[15\]
rlabel metal2 s 24518 15572 24518 15572 4 wrapped.spi_flash.shift_reg\[16\]
rlabel metal1 s 22586 14892 22586 14892 4 wrapped.spi_flash.shift_reg\[17\]
rlabel metal1 s 21528 15334 21528 15334 4 wrapped.spi_flash.shift_reg\[18\]
rlabel metal2 s 20286 15844 20286 15844 4 wrapped.spi_flash.shift_reg\[19\]
rlabel metal2 s 18814 15844 18814 15844 4 wrapped.spi_flash.shift_reg\[20\]
rlabel metal1 s 17710 15028 17710 15028 4 wrapped.spi_flash.shift_reg\[21\]
rlabel metal1 s 15042 14042 15042 14042 4 wrapped.spi_flash.shift_reg\[22\]
rlabel metal2 s 13202 13532 13202 13532 4 wrapped.spi_flash.shift_reg\[23\]
rlabel metal1 s 14766 11866 14766 11866 4 wrapped.spi_flash.shift_reg\[8\]
rlabel metal1 s 17204 12206 17204 12206 4 wrapped.spi_flash.shift_reg\[9\]
rlabel metal3 s 14214 15997 14214 15997 4 wrapped.spi_flash.timer\[0\]
rlabel metal1 s 14812 16762 14812 16762 4 wrapped.spi_flash.timer\[1\]
rlabel metal1 s 11224 16694 11224 16694 4 wrapped.spi_flash.timer\[2\]
rlabel metal2 s 10718 16796 10718 16796 4 wrapped.spi_flash.timer\[3\]
rlabel metal2 s 9522 16218 9522 16218 4 wrapped.spi_flash.timer\[4\]
flabel metal4 s 27256 496 27576 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 20540 496 20860 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 13824 496 14144 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7108 496 7428 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 23898 496 24218 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 17182 496 17502 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 10466 496 10786 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3750 496 4070 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 27158 17600 27214 18000 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal2 s 846 0 902 400 0 FreeSans 280 90 0 0 o_digital[0]
port 4 nsew
flabel metal2 s 18326 0 18382 400 0 FreeSans 280 90 0 0 o_digital[10]
port 5 nsew
flabel metal2 s 20074 0 20130 400 0 FreeSans 280 90 0 0 o_digital[11]
port 6 nsew
flabel metal2 s 21822 0 21878 400 0 FreeSans 280 90 0 0 o_digital[12]
port 7 nsew
flabel metal2 s 23570 0 23626 400 0 FreeSans 280 90 0 0 o_digital[13]
port 8 nsew
flabel metal2 s 25318 0 25374 400 0 FreeSans 280 90 0 0 o_digital[14]
port 9 nsew
flabel metal2 s 27066 0 27122 400 0 FreeSans 280 90 0 0 o_digital[15]
port 10 nsew
flabel metal2 s 2594 0 2650 400 0 FreeSans 280 90 0 0 o_digital[1]
port 11 nsew
flabel metal2 s 4342 0 4398 400 0 FreeSans 280 90 0 0 o_digital[2]
port 12 nsew
flabel metal2 s 6090 0 6146 400 0 FreeSans 280 90 0 0 o_digital[3]
port 13 nsew
flabel metal2 s 7838 0 7894 400 0 FreeSans 280 90 0 0 o_digital[4]
port 14 nsew
flabel metal2 s 9586 0 9642 400 0 FreeSans 280 90 0 0 o_digital[5]
port 15 nsew
flabel metal2 s 11334 0 11390 400 0 FreeSans 280 90 0 0 o_digital[6]
port 16 nsew
flabel metal2 s 13082 0 13138 400 0 FreeSans 280 90 0 0 o_digital[7]
port 17 nsew
flabel metal2 s 14830 0 14886 400 0 FreeSans 280 90 0 0 o_digital[8]
port 18 nsew
flabel metal2 s 16578 0 16634 400 0 FreeSans 280 90 0 0 o_digital[9]
port 19 nsew
flabel metal2 s 26514 17600 26570 18000 0 FreeSans 280 90 0 0 rst_n
port 20 nsew
flabel metal2 s 25870 17600 25926 18000 0 FreeSans 280 90 0 0 ui_in[0]
port 21 nsew
flabel metal2 s 25226 17600 25282 18000 0 FreeSans 280 90 0 0 ui_in[1]
port 22 nsew
flabel metal2 s 24582 17600 24638 18000 0 FreeSans 280 90 0 0 ui_in[2]
port 23 nsew
flabel metal2 s 23938 17600 23994 18000 0 FreeSans 280 90 0 0 ui_in[3]
port 24 nsew
flabel metal2 s 23294 17600 23350 18000 0 FreeSans 280 90 0 0 ui_in[4]
port 25 nsew
flabel metal2 s 22650 17600 22706 18000 0 FreeSans 280 90 0 0 ui_in[5]
port 26 nsew
flabel metal2 s 22006 17600 22062 18000 0 FreeSans 280 90 0 0 ui_in[6]
port 27 nsew
flabel metal2 s 21362 17600 21418 18000 0 FreeSans 280 90 0 0 ui_in[7]
port 28 nsew
flabel metal2 s 20718 17600 20774 18000 0 FreeSans 280 90 0 0 uio_in[0]
port 29 nsew
flabel metal2 s 20074 17600 20130 18000 0 FreeSans 280 90 0 0 uio_in[1]
port 30 nsew
flabel metal2 s 19430 17600 19486 18000 0 FreeSans 280 90 0 0 uio_in[2]
port 31 nsew
flabel metal2 s 18786 17600 18842 18000 0 FreeSans 280 90 0 0 uio_in[3]
port 32 nsew
flabel metal2 s 18142 17600 18198 18000 0 FreeSans 280 90 0 0 uio_in[4]
port 33 nsew
flabel metal2 s 17498 17600 17554 18000 0 FreeSans 280 90 0 0 uio_in[5]
port 34 nsew
flabel metal2 s 16854 17600 16910 18000 0 FreeSans 280 90 0 0 uio_in[6]
port 35 nsew
flabel metal2 s 16210 17600 16266 18000 0 FreeSans 280 90 0 0 uio_in[7]
port 36 nsew
flabel metal2 s 5262 17600 5318 18000 0 FreeSans 280 90 0 0 uio_oe[0]
port 37 nsew
flabel metal2 s 4618 17600 4674 18000 0 FreeSans 280 90 0 0 uio_oe[1]
port 38 nsew
flabel metal2 s 3974 17600 4030 18000 0 FreeSans 280 90 0 0 uio_oe[2]
port 39 nsew
flabel metal2 s 3330 17600 3386 18000 0 FreeSans 280 90 0 0 uio_oe[3]
port 40 nsew
flabel metal2 s 2686 17600 2742 18000 0 FreeSans 280 90 0 0 uio_oe[4]
port 41 nsew
flabel metal2 s 2042 17600 2098 18000 0 FreeSans 280 90 0 0 uio_oe[5]
port 42 nsew
flabel metal2 s 1398 17600 1454 18000 0 FreeSans 280 90 0 0 uio_oe[6]
port 43 nsew
flabel metal2 s 754 17600 810 18000 0 FreeSans 280 90 0 0 uio_oe[7]
port 44 nsew
flabel metal2 s 10414 17600 10470 18000 0 FreeSans 280 90 0 0 uio_out[0]
port 45 nsew
flabel metal2 s 9770 17600 9826 18000 0 FreeSans 280 90 0 0 uio_out[1]
port 46 nsew
flabel metal2 s 9126 17600 9182 18000 0 FreeSans 280 90 0 0 uio_out[2]
port 47 nsew
flabel metal2 s 8482 17600 8538 18000 0 FreeSans 280 90 0 0 uio_out[3]
port 48 nsew
flabel metal2 s 7838 17600 7894 18000 0 FreeSans 280 90 0 0 uio_out[4]
port 49 nsew
flabel metal2 s 7194 17600 7250 18000 0 FreeSans 280 90 0 0 uio_out[5]
port 50 nsew
flabel metal2 s 6550 17600 6606 18000 0 FreeSans 280 90 0 0 uio_out[6]
port 51 nsew
flabel metal2 s 5906 17600 5962 18000 0 FreeSans 280 90 0 0 uio_out[7]
port 52 nsew
flabel metal2 s 15566 17600 15622 18000 0 FreeSans 280 90 0 0 uo_out[0]
port 53 nsew
flabel metal2 s 14922 17600 14978 18000 0 FreeSans 280 90 0 0 uo_out[1]
port 54 nsew
flabel metal2 s 14278 17600 14334 18000 0 FreeSans 280 90 0 0 uo_out[2]
port 55 nsew
flabel metal2 s 13634 17600 13690 18000 0 FreeSans 280 90 0 0 uo_out[3]
port 56 nsew
flabel metal2 s 12990 17600 13046 18000 0 FreeSans 280 90 0 0 uo_out[4]
port 57 nsew
flabel metal2 s 12346 17600 12402 18000 0 FreeSans 280 90 0 0 uo_out[5]
port 58 nsew
flabel metal2 s 11702 17600 11758 18000 0 FreeSans 280 90 0 0 uo_out[6]
port 59 nsew
flabel metal2 s 11058 17600 11114 18000 0 FreeSans 280 90 0 0 uo_out[7]
port 60 nsew
<< properties >>
string FIXED_BBOX 0 0 28000 18000
string GDS_END 1940272
string GDS_FILE ../gds/digital_top.gds
string GDS_START 369032
<< end >>
