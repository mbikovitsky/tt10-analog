magic
tech sky130A
magscale 1 2
timestamp 1740246064
<< pwell >>
rect -201 -2582 201 2582
<< psubdiff >>
rect -165 2512 -69 2546
rect 69 2512 165 2546
rect -165 2450 -131 2512
rect 131 2450 165 2512
rect -165 -2512 -131 -2450
rect 131 -2512 165 -2450
rect -165 -2546 -69 -2512
rect 69 -2546 165 -2512
<< psubdiffcont >>
rect -69 2512 69 2546
rect -165 -2450 -131 2450
rect 131 -2450 165 2450
rect -69 -2546 69 -2512
<< xpolycontact >>
rect -35 1984 35 2416
rect -35 -2416 35 -1984
<< ppolyres >>
rect -35 -1984 35 1984
<< locali >>
rect -165 2512 -69 2546
rect 69 2512 165 2546
rect -165 2450 -131 2512
rect 131 2450 165 2512
rect -165 -2512 -131 -2450
rect 131 -2512 165 -2450
rect -165 -2546 -69 -2512
rect 69 -2546 165 -2512
<< viali >>
rect -19 2001 19 2398
rect -19 -2398 19 -2001
<< metal1 >>
rect -25 2398 25 2410
rect -25 2001 -19 2398
rect 19 2001 25 2398
rect -25 1989 25 2001
rect -25 -2001 25 -1989
rect -25 -2398 -19 -2001
rect 19 -2398 25 -2001
rect -25 -2410 25 -2398
<< properties >>
string FIXED_BBOX -148 -2529 148 2529
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 20.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 19.387k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
