magic
tech sky130A
magscale 1 2
timestamp 1740343563
<< viali >>
rect 4774 2046 4874 2080
rect 4650 188 4684 262
rect 890 -390 948 -220
rect 2460 -392 2534 -226
<< metal1 >>
rect 1818 7850 2742 8050
rect 438 3908 1164 4108
rect 438 200 638 3908
rect 964 3212 1164 3908
rect 14 0 638 200
rect 1818 -200 2018 7850
rect 2542 7112 2742 7850
rect 3654 4320 3854 8200
rect 3654 4120 4918 4320
rect 3654 2188 3854 4120
rect 4718 3652 4918 4120
rect 4052 2994 4808 3594
rect 4838 2994 6984 3594
rect 4052 2246 4808 2846
rect 4838 2334 6178 2846
rect 4838 2246 6180 2334
rect 3654 2142 4856 2188
rect 3654 2054 3854 2142
rect 4724 2080 4924 2104
rect 4724 2046 4774 2080
rect 4874 2046 4924 2080
rect 4724 1898 4924 2046
rect 3130 1698 4924 1898
rect 3130 -200 3330 1698
rect 16 -220 3330 -200
rect 16 -390 890 -220
rect 948 -226 3330 -220
rect 948 -390 2460 -226
rect 16 -392 2460 -390
rect 2534 -392 3330 -226
rect 16 -400 3330 -392
rect 3691 1433 4905 1595
rect 992 -1517 1154 -894
rect 2563 -1517 2725 -983
rect 3691 -1517 3853 1433
rect 4743 1311 4905 1433
rect 5580 1256 6180 2246
rect 4054 656 4810 1256
rect 4840 656 6180 1256
rect 6384 508 6984 2994
rect 4054 262 4810 508
rect 4054 188 4650 262
rect 4684 188 4810 262
rect 4054 -92 4810 188
rect 4840 -92 6984 508
rect 4739 -1517 4901 -149
rect 992 -1679 4901 -1517
rect 5904 -2066 6104 -92
use sky130_fd_pr__nfet_01v8_lvt_KBNS5F  XM1
timestamp 1740246064
transform 1 0 4825 0 1 582
box -211 -910 211 910
use sky130_fd_pr__nfet_01v8_lvt_KBNS5F  XM3
timestamp 1740246064
transform 1 0 4823 0 1 2920
box -211 -910 211 910
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR5
timestamp 1740246064
transform 1 0 2641 0 1 3090
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR6
timestamp 1740246064
transform 1 0 1065 0 1 1158
box -201 -2582 201 2582
<< labels >>
flabel metal1 3654 8000 3854 8200 0 FreeSans 256 0 0 0 in
port 3 nsew
flabel metal1 14 0 214 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 4052 2246 4252 2446 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 4052 2994 4252 3194 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 16 -400 216 -200 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 5904 -2066 6104 -1866 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 4054 -92 4254 108 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 4054 656 4254 856 0 FreeSans 256 0 0 0 VSS
port 1 nsew
<< end >>
