magic
tech sky130A
magscale 1 2
timestamp 1740253518
<< viali >>
rect -5990 1020 -5932 1196
rect -5498 1020 -5438 1198
rect -4220 1014 -4170 1198
rect -3666 1018 -3618 1196
rect -2636 1128 -2572 1306
rect -2116 1132 -2056 1302
rect -998 1054 -946 1218
rect -520 1048 -466 1208
rect 540 1020 612 1182
rect 1042 1018 1104 1186
rect 2080 1056 2142 1222
rect 2468 1060 2532 1222
rect 3432 1016 3496 1184
rect 3780 1020 3852 1178
rect 4826 1006 4880 1184
rect 5142 1012 5202 1182
rect 6216 902 6274 1072
rect 6542 906 6600 1066
<< metal1 >>
rect -6918 8236 -6010 8436
rect -6918 670 -6718 8236
rect -6210 7624 -6010 8236
rect -5416 7660 -5216 8620
rect -3598 7602 -3398 8626
rect -2040 7754 -1840 8744
rect -430 7766 -230 8746
rect 1114 7756 1314 8746
rect 2562 7890 2762 8748
rect 3864 7926 4064 8748
rect 5226 7898 5426 8748
rect 6608 7948 6808 8872
rect -4902 4312 -4280 4456
rect -6022 1196 -5826 1212
rect -6022 1020 -5990 1196
rect -5932 1020 -5826 1196
rect -6022 1012 -5826 1020
rect -5626 1198 -5408 1212
rect -5626 1020 -5498 1198
rect -5438 1020 -5408 1198
rect -5626 1012 -5408 1020
rect -6918 470 -6600 670
rect -6400 470 -6394 670
rect -6184 -1060 -6044 -476
rect -5386 -1040 -5246 -400
rect -4902 -1040 -4758 4312
rect -4424 3660 -4280 4312
rect -3176 4350 -2688 4494
rect -4252 1198 -4042 1208
rect -4252 1014 -4220 1198
rect -4170 1014 -4042 1198
rect -4252 1008 -4042 1014
rect -3842 1196 -3592 1208
rect -3842 1018 -3666 1196
rect -3618 1018 -3592 1196
rect -3842 1008 -3592 1018
rect -5386 -1060 -4758 -1040
rect -6184 -1184 -4758 -1060
rect -4413 -1107 -4279 -589
rect -3572 -1096 -3438 -460
rect -3176 -1096 -3032 4350
rect -2832 3680 -2688 4350
rect -1634 4396 -1054 4552
rect -2664 1306 -2458 1320
rect -2664 1128 -2636 1306
rect -2572 1128 -2458 1306
rect -2664 1120 -2458 1128
rect -2258 1302 -2024 1320
rect -2258 1132 -2116 1302
rect -2056 1132 -2024 1302
rect -2258 1120 -2024 1132
rect -3572 -1107 -3032 -1096
rect -6184 -1200 -5246 -1184
rect -4413 -1240 -3032 -1107
rect -2836 -1000 -2676 -592
rect -2024 -988 -1864 -292
rect -1634 -988 -1478 4396
rect -1210 3740 -1054 4396
rect -41 4413 494 4563
rect -830 1236 -630 1242
rect -1034 1218 -830 1236
rect -1034 1054 -998 1218
rect -946 1054 -830 1218
rect -1034 1036 -830 1054
rect -630 1208 -430 1236
rect -630 1048 -520 1208
rect -466 1048 -430 1208
rect -630 1036 -430 1048
rect -830 1030 -630 1036
rect -2024 -1000 -1478 -988
rect -2836 -1144 -1478 -1000
rect -1191 -993 -1053 -315
rect -420 -969 -282 -272
rect -41 -969 109 4413
rect 344 3720 494 4413
rect 1554 4532 2026 4680
rect 510 1182 720 1208
rect 510 1020 540 1182
rect 612 1020 720 1182
rect 510 1008 720 1020
rect 920 1186 1144 1208
rect 920 1018 1042 1186
rect 1104 1018 1144 1186
rect 920 1008 1144 1018
rect -420 -993 109 -969
rect -1191 -1119 109 -993
rect 353 -935 499 -315
rect 1142 -922 1288 -260
rect 1554 -922 1702 4532
rect 1878 3844 2026 4532
rect 2922 4632 3390 4796
rect 2058 1222 2188 1244
rect 2058 1056 2080 1222
rect 2142 1056 2188 1222
rect 2058 1044 2188 1056
rect 2388 1222 2570 1244
rect 2388 1060 2468 1222
rect 2532 1060 2570 1222
rect 2388 1044 2570 1060
rect 1142 -935 1702 -922
rect 353 -1070 1702 -935
rect 1896 -904 2032 -220
rect 2572 -874 2708 -162
rect 2922 -874 3086 4632
rect 3226 3948 3390 4632
rect 4283 4623 4778 4773
rect 3396 1184 3526 1206
rect 3396 1016 3432 1184
rect 3496 1016 3526 1184
rect 3396 1006 3526 1016
rect 3726 1178 3898 1206
rect 3726 1020 3780 1178
rect 3852 1020 3898 1178
rect 3726 1006 3898 1020
rect 2572 -904 3086 -874
rect 1896 -1038 3086 -904
rect 3247 -841 3389 -121
rect 3900 -817 4042 -88
rect 4283 -817 4433 4623
rect 4628 3880 4778 4623
rect 5622 4504 6160 4652
rect 4800 1184 4908 1198
rect 4800 1006 4826 1184
rect 4880 1006 4908 1184
rect 4800 998 4908 1006
rect 5108 1182 5244 1198
rect 5108 1012 5142 1182
rect 5202 1012 5244 1182
rect 5108 998 5244 1012
rect 3900 -841 4433 -817
rect 3247 -967 4433 -841
rect 4633 -815 4787 -163
rect 5244 -815 5398 -146
rect 4633 -824 5398 -815
rect 5622 -824 5770 4504
rect 6012 3918 6160 4504
rect 6172 1072 6298 1086
rect 6172 902 6216 1072
rect 6274 902 6298 1072
rect 6172 886 6298 902
rect 6498 1066 6654 1086
rect 6498 906 6542 1066
rect 6600 906 6654 1066
rect 6498 886 6654 906
rect 3247 -983 4042 -967
rect 4633 -969 5770 -824
rect 6016 -698 6172 -118
rect 6632 -698 6788 -80
rect 6016 -854 6788 -698
rect 5252 -972 5770 -969
rect 1896 -1040 2708 -1038
rect 353 -1081 1288 -1070
rect -1191 -1131 -282 -1119
rect -2836 -1160 -1864 -1144
rect -4413 -1241 -3438 -1240
rect 6328 -1472 6528 -854
<< via1 >>
rect -5826 1012 -5626 1212
rect -6600 470 -6400 670
rect -4042 1008 -3842 1208
rect -2458 1120 -2258 1320
rect -830 1036 -630 1236
rect 720 1008 920 1208
rect 2188 1044 2388 1244
rect 3526 1006 3726 1206
rect 4908 998 5108 1198
rect 6298 886 6498 1086
<< metal2 >>
rect -2458 1320 -2258 1326
rect -5826 1212 -5626 1218
rect -6600 670 -6400 676
rect -5826 670 -5626 1012
rect -4042 1208 -3842 1214
rect -4042 670 -3842 1008
rect 2188 1244 2388 1250
rect -2458 670 -2258 1120
rect -836 1036 -830 1236
rect -630 1036 -624 1236
rect 720 1208 920 1214
rect -830 670 -630 1036
rect 720 670 920 1008
rect 2188 670 2388 1044
rect 3526 1206 3726 1212
rect 3526 670 3726 1006
rect 4908 1198 5108 1204
rect 4908 670 5108 998
rect 6298 1086 6498 1092
rect 6298 670 6498 886
rect -6400 470 7384 670
rect -6600 464 -6400 470
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR1
timestamp 1740251180
transform 1 0 -5321 0 1 3636
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR2
timestamp 1740251180
transform 1 0 -3493 0 1 3568
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR3
timestamp 1740251180
transform 1 0 -6111 0 1 3618
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR4
timestamp 1740251180
transform 1 0 -4343 0 1 1610
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR5
timestamp 1740251180
transform 1 0 -1937 0 1 3732
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR6
timestamp 1740251180
transform 1 0 -2753 0 1 1648
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR7
timestamp 1740251180
transform 1 0 -345 0 1 3746
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR8
timestamp 1740251180
transform 1 0 -1121 0 1 1718
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR9
timestamp 1740251180
transform 1 0 1221 0 1 3748
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR10
timestamp 1740251180
transform 1 0 425 0 1 1720
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR11
timestamp 1740251180
transform 1 0 2647 0 1 3866
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR12
timestamp 1740251180
transform 1 0 1963 0 1 1824
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR13
timestamp 1740251180
transform 1 0 3965 0 1 3928
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR14
timestamp 1740251180
transform 1 0 3319 0 1 1928
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR15
timestamp 1740251180
transform 1 0 6717 0 1 3934
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR16
timestamp 1740251180
transform 1 0 6097 0 1 1918
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR17
timestamp 1740251180
transform 1 0 5321 0 1 3880
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR18
timestamp 1740251180
transform 1 0 4709 0 1 1866
box -201 -2582 201 2582
<< labels >>
flabel metal1 -5416 8420 -5216 8620 0 FreeSans 256 0 0 0 a0
port 9 nsew
flabel metal1 -3598 8426 -3398 8626 0 FreeSans 256 0 0 0 a1
port 2 nsew
flabel metal1 -2040 8544 -1840 8744 0 FreeSans 256 0 0 0 a2
port 7 nsew
flabel metal1 -430 8546 -230 8746 0 FreeSans 256 0 0 0 a3
port 3 nsew
flabel metal1 1114 8546 1314 8746 0 FreeSans 256 0 0 0 a4
port 4 nsew
flabel metal1 2562 8548 2762 8748 0 FreeSans 256 0 0 0 a5
port 5 nsew
flabel metal1 3864 8548 4064 8748 0 FreeSans 256 0 0 0 a6
port 6 nsew
flabel metal1 5226 8548 5426 8748 0 FreeSans 256 0 0 0 a7
port 8 nsew
flabel metal1 6328 -1472 6528 -1272 0 FreeSans 256 0 0 0 out
port 10 nsew
flabel metal1 -6918 470 -6718 670 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 6608 8672 6808 8872 0 FreeSans 256 0 0 0 VDD
port 0 nsew
<< end >>
