magic
tech sky130A
magscale 1 2
timestamp 1757772008
<< metal1 >>
rect 29370 22324 29376 22524
rect 29576 22324 29894 22524
rect 15026 22158 15226 22164
rect 15026 21704 15226 21958
rect 29694 21710 29894 22324
rect 14746 11428 14946 11766
rect 26664 11566 29614 11766
rect 14746 11228 18440 11428
rect 18240 10978 18440 11228
rect 26664 10996 26866 11566
rect 18594 6590 19194 6596
rect 18594 5984 19194 5990
rect 27022 6590 27622 6596
rect 27022 5984 27622 5990
rect 18588 5842 19188 5848
rect 18588 5236 19188 5242
rect 27008 5842 27608 5848
rect 27008 5236 27608 5242
rect 23026 4864 23226 4870
rect 14612 4728 14812 4734
rect 14612 2998 14812 4528
rect 18594 4252 19194 4258
rect 18594 3646 19194 3652
rect 18584 3502 19180 3508
rect 23026 2996 23226 4664
rect 27032 4252 27632 4258
rect 27032 3646 27632 3652
rect 27034 3502 27630 3508
rect 18584 2900 19180 2906
rect 27034 2900 27630 2906
rect 13696 2598 13702 2798
rect 13902 2598 14802 2798
rect 22334 2796 22534 2802
rect 22534 2596 23228 2796
rect 22334 2590 22534 2596
rect 20490 738 20690 1132
rect 28916 746 29116 1130
rect 28916 540 29116 546
rect 20490 532 20690 538
<< via1 >>
rect 29376 22324 29576 22524
rect 15026 21958 15226 22158
rect 18594 5990 19194 6590
rect 27022 5990 27622 6590
rect 18588 5242 19188 5842
rect 27008 5242 27608 5842
rect 14612 4528 14812 4728
rect 23026 4664 23226 4864
rect 18594 3652 19194 4252
rect 18584 2906 19180 3502
rect 27032 3652 27632 4252
rect 27034 2906 27630 3502
rect 13702 2598 13902 2798
rect 22334 2596 22534 2796
rect 20490 538 20690 738
rect 28916 546 29116 746
<< metal2 >>
rect 15026 22526 15226 22535
rect 29376 22524 29576 22530
rect 15026 22158 15226 22326
rect 29077 22324 29086 22524
rect 29286 22324 29376 22524
rect 29376 22318 29576 22324
rect 15020 21958 15026 22158
rect 15226 21958 15232 22158
rect 15442 13508 16876 13708
rect 2555 5990 2564 6590
rect 3164 5990 18594 6590
rect 19194 5990 27022 6590
rect 27622 5990 27628 6590
rect 2553 5242 2562 5842
rect 3162 5242 18588 5842
rect 19188 5242 27008 5842
rect 27608 5242 27614 5842
rect 14612 4728 14812 5242
rect 23026 4864 23226 5242
rect 14606 4528 14612 4728
rect 14812 4528 14818 4728
rect 23020 4664 23026 4864
rect 23226 4664 23232 4864
rect 4167 3652 4176 4252
rect 4776 3652 18594 4252
rect 19194 3652 27032 4252
rect 27632 3652 27638 4252
rect 4169 2906 4178 3502
rect 4774 2906 18584 3502
rect 19180 2906 27034 3502
rect 27630 2906 27636 3502
rect 13702 2798 13902 2906
rect 22334 2796 22534 2906
rect 13702 2592 13902 2598
rect 22328 2596 22334 2796
rect 22534 2596 22540 2796
rect 20484 538 20490 738
rect 20690 538 22502 738
rect 22702 538 22711 738
rect 28910 546 28916 746
rect 29116 546 29270 746
rect 29470 546 29479 746
<< via2 >>
rect 15026 22326 15226 22526
rect 29086 22324 29286 22524
rect 2564 5990 3164 6590
rect 2562 5242 3162 5842
rect 4176 3652 4776 4252
rect 4178 2906 4774 3502
rect 22502 538 22702 738
rect 29270 546 29470 746
<< metal3 >>
rect 5441 23964 5759 23965
rect 5436 23648 5442 23964
rect 5758 23648 5764 23964
rect 18872 23863 19192 23864
rect 12156 23773 12476 23774
rect 5441 22604 5759 23648
rect 12151 23455 12157 23773
rect 12475 23455 12481 23773
rect 18867 23545 18873 23863
rect 19191 23545 19197 23863
rect 25588 23739 25908 23740
rect 12156 22604 12476 23455
rect 18872 22606 19192 23545
rect 25583 23421 25589 23739
rect 25907 23421 25913 23739
rect 25588 22606 25908 23421
rect 18872 22604 25908 22606
rect 5441 22591 25908 22604
rect 205 22273 211 22591
rect 529 22526 25908 22591
rect 529 22326 15026 22526
rect 15226 22524 25908 22526
rect 29081 22524 29291 22529
rect 15226 22326 29086 22524
rect 529 22324 29086 22326
rect 29286 22324 29291 22524
rect 529 22286 25908 22324
rect 29081 22319 29291 22324
rect 529 22284 19192 22286
rect 529 22273 5759 22284
rect 2559 6590 3169 6595
rect 216 6584 2564 6590
rect 216 5996 222 6584
rect 594 5996 2564 6584
rect 216 5990 2564 5996
rect 3164 5990 3169 6590
rect 2559 5985 3169 5990
rect 2557 5842 3167 5847
rect 210 5836 2562 5842
rect 210 5248 216 5836
rect 594 5248 2562 5836
rect 210 5242 2562 5248
rect 3162 5242 3167 5842
rect 2557 5237 3167 5242
rect 4171 4252 4781 4257
rect 3206 3652 3212 4252
rect 3812 3652 4176 4252
rect 4776 3652 4781 4252
rect 4171 3647 4781 3652
rect 4173 3502 4779 3507
rect 3186 2906 3192 3502
rect 3788 2906 4178 3502
rect 4774 2906 4779 3502
rect 4173 2901 4779 2906
rect 29265 746 29475 751
rect 22497 738 22707 743
rect 22497 538 22502 738
rect 22702 538 24722 738
rect 24922 538 24928 738
rect 29265 546 29270 746
rect 29470 546 29682 746
rect 29882 546 29888 746
rect 29265 541 29475 546
rect 22497 533 22707 538
<< via3 >>
rect 5442 23648 5758 23964
rect 12157 23455 12475 23773
rect 18873 23545 19191 23863
rect 25589 23421 25907 23739
rect 211 22273 529 22591
rect 222 5996 594 6584
rect 216 5248 594 5836
rect 3212 3652 3812 4252
rect 3192 2906 3788 3502
rect 24722 538 24922 738
rect 29682 546 29882 746
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 22591 600 44152
rect 200 22273 211 22591
rect 529 22273 600 22591
rect 200 6584 600 22273
rect 200 5996 222 6584
rect 594 5996 600 6584
rect 200 5836 600 5996
rect 200 5248 216 5836
rect 594 5248 600 5836
rect 200 1000 600 5248
rect 800 23122 1200 44152
rect 5441 23964 5759 24526
rect 5441 23648 5442 23964
rect 5758 23648 5759 23964
rect 5441 23647 5759 23648
rect 8798 23122 9118 24496
rect 12156 23773 12476 24524
rect 12156 23455 12157 23773
rect 12475 23455 12476 23773
rect 12156 23454 12476 23455
rect 15514 23122 15834 24492
rect 18872 23863 19192 24582
rect 18872 23545 18873 23863
rect 19191 23545 19192 23863
rect 18872 23544 19192 23545
rect 22230 23122 22550 24490
rect 25588 23739 25908 24484
rect 25588 23421 25589 23739
rect 25907 23421 25908 23739
rect 25588 23420 25908 23421
rect 28946 23122 29266 24490
rect 800 22802 29266 23122
rect 800 4252 1200 22802
rect 3211 4252 3813 4253
rect 800 3652 3212 4252
rect 3812 3652 3813 4252
rect 800 3502 1200 3652
rect 3211 3651 3813 3652
rect 3191 3502 3789 3503
rect 800 2906 3192 3502
rect 3788 2906 3789 3502
rect 800 1000 1200 2906
rect 3191 2905 3789 2906
rect 29681 746 29883 747
rect 24721 738 24923 739
rect 24721 538 24722 738
rect 24922 538 26682 738
rect 29681 546 29682 746
rect 29882 730 29883 746
rect 29882 550 30542 730
rect 29882 546 29883 550
rect 29681 545 29883 546
rect 24721 537 24923 538
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 538
rect 30362 0 30542 550
use buffer  buffer_0
timestamp 1740347555
transform 1 0 23012 0 1 2996
box 14 -2066 6984 8200
use buffer  buffer_2
timestamp 1740347555
transform 1 0 14586 0 1 2998
box 14 -2066 6984 8200
use dac  dac_1
timestamp 1740347555
transform 1 0 23086 0 1 13038
box -6918 -1472 7384 8872
use dac  dac_2
timestamp 1740347555
transform 1 0 8418 0 1 13038
box -6918 -1472 7384 8872
use digital_top  digital_top_0
timestamp 1757770450
transform 1 0 1690 0 1 23594
box 514 0 27576 18000
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
