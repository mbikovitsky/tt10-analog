magic
tech sky130A
magscale 1 2
timestamp 1740250525
<< viali >>
rect 4640 2302 4688 2484
rect 4640 442 4690 622
rect 890 -390 948 -220
rect 2460 -392 2534 -226
<< metal1 >>
rect 1818 7850 2742 8050
rect 438 3908 1164 4108
rect 438 200 638 3908
rect 964 3212 1164 3908
rect 1818 1210 2018 7850
rect 2542 7112 2742 7850
rect 3654 4320 3854 8200
rect 3654 4120 4918 4320
rect 3654 3938 3854 4120
rect 3654 3732 3854 3738
rect 4718 3652 4918 4120
rect 2980 3118 4802 3608
rect 2974 3086 4802 3118
rect 2974 2862 3174 3086
rect 4280 2862 4802 3086
rect 4836 3016 5402 3608
rect 4836 2992 5416 3016
rect 2974 2685 4802 2862
rect 4840 2698 5416 2992
rect 5590 2698 6166 3016
rect 2974 2662 4800 2685
rect 1812 1010 1818 1210
rect 2018 1010 2024 1210
rect 2974 200 3174 2662
rect 4840 2596 6166 2698
rect 3322 2484 4704 2496
rect 3322 2302 4640 2484
rect 4688 2302 4704 2484
rect 3322 2296 4704 2302
rect 0 0 3178 200
rect 1818 -200 2018 -194
rect 3322 -200 3522 2296
rect 4842 2226 6166 2596
rect 4722 1888 4922 2190
rect 4716 1688 4722 1888
rect 4922 1688 4928 1888
rect 3691 1433 4905 1595
rect 5104 1472 6166 2226
rect 3691 411 3853 1433
rect 4743 1311 4905 1433
rect 4420 632 4816 1274
rect 4254 622 4816 632
rect 4254 442 4640 622
rect 4690 442 4816 622
rect 3685 249 3691 411
rect 3853 249 3859 411
rect 4254 -112 4816 442
rect 4844 812 5420 1278
rect 5590 812 6166 1472
rect 4844 236 6166 812
rect 4844 -108 5420 236
rect 4254 -200 4454 -112
rect 0 -220 1818 -200
rect 0 -390 890 -220
rect 948 -390 1818 -220
rect 0 -400 1818 -390
rect 2018 -226 4454 -200
rect 2018 -392 2460 -226
rect 2534 -392 4454 -226
rect 2018 -400 4454 -392
rect 1818 -406 2018 -400
rect 3691 -825 3853 -819
rect 992 -1517 1154 -894
rect 2563 -1517 2725 -983
rect 3691 -1517 3853 -987
rect 4739 -1517 4901 -149
rect 5928 -876 6128 236
rect 992 -1679 4901 -1517
<< via1 >>
rect 3654 3738 3854 3938
rect 1818 1010 2018 1210
rect 4722 1688 4922 1888
rect 3691 249 3853 411
rect 1818 -400 2018 -200
rect 3691 -987 3853 -825
<< metal2 >>
rect 3648 3738 3654 3938
rect 3854 3738 3860 3938
rect 3654 1888 3854 3738
rect 4722 1888 4922 1894
rect 3654 1688 4722 1888
rect 4722 1682 4922 1688
rect 1818 1210 2018 1216
rect 1818 -200 2018 1010
rect 3691 411 3853 417
rect 1812 -400 1818 -200
rect 2018 -400 2024 -200
rect 3691 -825 3853 249
rect 3685 -987 3691 -825
rect 3853 -987 3859 -825
use sky130_fd_pr__nfet_01v8_lvt_KBNS5F  XM1
timestamp 1740246064
transform 1 0 4825 0 1 582
box -211 -910 211 910
use sky130_fd_pr__nfet_01v8_lvt_KBNS5F  XM3
timestamp 1740246064
transform 1 0 4823 0 1 2920
box -211 -910 211 910
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR5
timestamp 1740246064
transform 1 0 2641 0 1 3090
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR6
timestamp 1740246064
transform 1 0 1065 0 1 1158
box -201 -2582 201 2582
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 3654 8000 3854 8200 0 FreeSans 256 0 0 0 in
port 3 nsew
flabel metal1 5928 -876 6128 -676 0 FreeSans 256 0 0 0 out
port 2 nsew
<< end >>
