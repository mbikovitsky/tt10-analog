magic
tech sky130A
magscale 1 2
timestamp 1757774869
<< metal1 >>
rect 29370 22324 29376 22524
rect 29576 22324 29894 22524
rect 15026 22158 15226 22164
rect 12360 21724 12416 21730
rect 6454 21716 6510 21722
rect 6454 21654 6510 21660
rect 8054 21712 8110 21718
rect 11056 21716 11112 21722
rect 9600 21656 9606 21712
rect 9662 21656 9668 21712
rect 12360 21662 12416 21668
rect 8054 21650 8110 21656
rect 11056 21654 11112 21660
rect 13710 21656 13716 21712
rect 13772 21656 13778 21712
rect 15026 21704 15226 21958
rect 21112 21710 21168 21716
rect 24270 21714 24326 21720
rect 21112 21648 21168 21654
rect 22720 21698 22776 21704
rect 24270 21652 24326 21658
rect 25718 21710 25774 21716
rect 27002 21654 27008 21710
rect 27064 21654 27070 21710
rect 28376 21706 28432 21712
rect 29694 21710 29894 22324
rect 25718 21648 25774 21654
rect 28376 21644 28432 21650
rect 22720 21636 22776 21642
rect 19560 21596 19616 21602
rect 4886 21582 4942 21588
rect 3066 21506 3072 21562
rect 3128 21506 3134 21562
rect 4886 21520 4942 21526
rect 17738 21518 17744 21574
rect 17800 21518 17806 21574
rect 19560 21534 19616 21540
rect 14746 11428 14946 11766
rect 26664 11566 29614 11766
rect 14746 11228 18440 11428
rect 18240 10978 18440 11228
rect 26664 10996 26866 11566
rect 18594 6590 19194 6596
rect 18594 5984 19194 5990
rect 27022 6590 27622 6596
rect 27022 5984 27622 5990
rect 18588 5842 19188 5848
rect 18588 5236 19188 5242
rect 27008 5842 27608 5848
rect 27008 5236 27608 5242
rect 23026 4864 23226 4870
rect 14612 4728 14812 4734
rect 14612 2998 14812 4528
rect 18594 4252 19194 4258
rect 18594 3646 19194 3652
rect 18584 3502 19180 3508
rect 23026 2996 23226 4664
rect 27032 4252 27632 4258
rect 27032 3646 27632 3652
rect 27034 3502 27630 3508
rect 18584 2900 19180 2906
rect 27034 2900 27630 2906
rect 13696 2598 13702 2798
rect 13902 2598 14802 2798
rect 22334 2796 22534 2802
rect 22534 2596 23228 2796
rect 22334 2590 22534 2596
rect 20490 738 20690 1132
rect 28916 746 29116 1130
rect 28916 540 29116 546
rect 20490 532 20690 538
<< via1 >>
rect 29376 22324 29576 22524
rect 15026 21958 15226 22158
rect 6454 21660 6510 21716
rect 8054 21656 8110 21712
rect 9606 21656 9662 21712
rect 11056 21660 11112 21716
rect 12360 21668 12416 21724
rect 13716 21656 13772 21712
rect 21112 21654 21168 21710
rect 22720 21642 22776 21698
rect 24270 21658 24326 21714
rect 25718 21654 25774 21710
rect 27008 21654 27064 21710
rect 28376 21650 28432 21706
rect 3072 21506 3128 21562
rect 4886 21526 4942 21582
rect 17744 21518 17800 21574
rect 19560 21540 19616 21596
rect 18594 5990 19194 6590
rect 27022 5990 27622 6590
rect 18588 5242 19188 5842
rect 27008 5242 27608 5842
rect 14612 4528 14812 4728
rect 23026 4664 23226 4864
rect 18594 3652 19194 4252
rect 18584 2906 19180 3502
rect 27032 3652 27632 4252
rect 27034 2906 27630 3502
rect 13702 2598 13902 2798
rect 22334 2596 22534 2796
rect 20490 538 20690 738
rect 28916 546 29116 746
<< metal2 >>
rect 2442 44862 2502 44871
rect 2442 44793 2502 44802
rect 2444 41522 2500 44793
rect 3086 44710 3146 44719
rect 3086 44641 3146 44650
rect 3088 41534 3144 44641
rect 3730 44578 3790 44587
rect 3730 44509 3790 44518
rect 28846 44518 28906 44527
rect 3732 41538 3788 44509
rect 23246 44504 23306 44506
rect 20486 44500 20546 44502
rect 22694 44500 22754 44502
rect 19934 44498 19994 44500
rect 19382 44486 19442 44488
rect 17726 44478 17786 44480
rect 18278 44478 18338 44480
rect 18830 44478 18890 44480
rect 4374 44434 4434 44443
rect 17719 44422 17728 44478
rect 17784 44422 17793 44478
rect 18271 44422 18280 44478
rect 18336 44422 18345 44478
rect 18823 44422 18832 44478
rect 18888 44422 18897 44478
rect 19375 44430 19384 44486
rect 19440 44430 19449 44486
rect 19927 44442 19936 44498
rect 19992 44442 20001 44498
rect 20479 44444 20488 44500
rect 20544 44444 20553 44500
rect 21038 44498 21098 44500
rect 21590 44498 21650 44500
rect 22142 44498 22202 44500
rect 4374 44365 4434 44374
rect 4376 41538 4432 44365
rect 5020 44308 5076 44315
rect 5018 44306 5078 44308
rect 5018 44250 5020 44306
rect 5076 44250 5078 44306
rect 5018 41490 5078 44250
rect 5668 44168 5724 44175
rect 5666 44166 5726 44168
rect 5666 44110 5668 44166
rect 5724 44110 5726 44166
rect 5666 41512 5726 44110
rect 6308 44036 6364 44043
rect 6306 44034 6366 44036
rect 6306 43978 6308 44034
rect 6364 43978 6366 44034
rect 17726 44014 17786 44422
rect 6306 41504 6366 43978
rect 15962 43954 17786 44014
rect 6950 43908 7006 43915
rect 6948 43906 7008 43908
rect 6948 43850 6950 43906
rect 7006 43850 7008 43906
rect 6948 41482 7008 43850
rect 7598 43780 7654 43787
rect 7596 43778 7656 43780
rect 7596 43722 7598 43778
rect 7654 43722 7656 43778
rect 7596 41476 7656 43722
rect 8238 43656 8294 43663
rect 8236 43654 8296 43656
rect 8236 43598 8238 43654
rect 8294 43598 8296 43654
rect 8236 41476 8296 43598
rect 8886 43510 8942 43517
rect 8884 43508 8944 43510
rect 8884 43452 8886 43508
rect 8942 43452 8944 43508
rect 8884 41460 8944 43452
rect 9528 43356 9584 43363
rect 9526 43354 9586 43356
rect 9526 43298 9528 43354
rect 9584 43298 9586 43354
rect 9526 41504 9586 43298
rect 10164 43204 10224 43206
rect 10157 43148 10166 43204
rect 10222 43148 10231 43204
rect 10164 41472 10224 43148
rect 10814 43062 10870 43069
rect 10812 43060 10872 43062
rect 10812 43004 10814 43060
rect 10870 43004 10872 43060
rect 10812 41516 10872 43004
rect 11458 42908 11514 42915
rect 11456 42906 11516 42908
rect 11456 42850 11458 42906
rect 11514 42850 11516 42906
rect 11456 41482 11516 42850
rect 12100 42766 12156 42773
rect 12098 42764 12158 42766
rect 12098 42708 12100 42764
rect 12156 42708 12158 42764
rect 12098 41504 12158 42708
rect 12750 42620 12806 42627
rect 12748 42618 12808 42620
rect 12748 42562 12750 42618
rect 12806 42562 12808 42618
rect 12748 41490 12808 42562
rect 13388 42480 13444 42487
rect 13386 42478 13446 42480
rect 13386 42422 13388 42478
rect 13444 42422 13446 42478
rect 13386 41490 13446 42422
rect 14036 42344 14092 42351
rect 14034 42342 14094 42344
rect 14034 42286 14036 42342
rect 14092 42286 14094 42342
rect 14034 41482 14094 42286
rect 14669 41540 14678 41596
rect 14734 41540 14743 41596
rect 15313 41524 15322 41580
rect 15378 41524 15387 41580
rect 15962 41530 16022 43954
rect 18278 43868 18338 44422
rect 16614 43808 18338 43868
rect 16614 41534 16674 43808
rect 18830 43740 18890 44422
rect 17250 43680 18890 43740
rect 17250 41522 17310 43680
rect 19382 43572 19442 44430
rect 17898 43512 19442 43572
rect 17898 41512 17958 43512
rect 19934 43436 19994 44442
rect 18540 43376 19994 43436
rect 18540 41492 18600 43376
rect 20486 43290 20546 44444
rect 21031 44442 21040 44498
rect 21096 44442 21105 44498
rect 21583 44442 21592 44498
rect 21648 44442 21657 44498
rect 22135 44442 22144 44498
rect 22200 44442 22209 44498
rect 22687 44444 22696 44500
rect 22752 44444 22761 44500
rect 23239 44448 23248 44504
rect 23304 44448 23313 44504
rect 23798 44500 23858 44502
rect 25454 44500 25514 44502
rect 26006 44500 26066 44502
rect 19186 43230 20546 43290
rect 19186 41492 19246 43230
rect 21038 43156 21098 44442
rect 19826 43096 21098 43156
rect 19826 41548 19886 43096
rect 21590 42976 21650 44442
rect 20476 42916 21650 42976
rect 20476 41518 20536 42916
rect 22142 42834 22202 44442
rect 21118 42774 22202 42834
rect 21118 41514 21178 42774
rect 22694 42622 22754 44444
rect 21760 42562 22754 42622
rect 21760 41548 21820 42562
rect 23246 42440 23306 44448
rect 23791 44444 23800 44500
rect 23856 44444 23865 44500
rect 24350 44498 24410 44500
rect 24902 44498 24962 44500
rect 22404 42380 23306 42440
rect 22404 41536 22464 42380
rect 23798 42254 23858 44444
rect 24343 44442 24352 44498
rect 24408 44442 24417 44498
rect 24895 44442 24904 44498
rect 24960 44442 24969 44498
rect 25447 44444 25456 44500
rect 25512 44444 25521 44500
rect 25999 44444 26008 44500
rect 26064 44444 26073 44500
rect 27110 44498 27170 44500
rect 26558 44494 26618 44496
rect 23054 42194 23858 42254
rect 23054 41536 23114 42194
rect 24350 42078 24410 44442
rect 23692 42018 24410 42078
rect 23692 41526 23752 42018
rect 24902 41830 24962 44442
rect 24338 41770 24962 41830
rect 24338 41508 24398 41770
rect 25454 41596 25514 44444
rect 24978 41536 25514 41596
rect 26006 41594 26066 44444
rect 26551 44438 26560 44494
rect 26616 44438 26625 44494
rect 27103 44442 27112 44498
rect 27168 44442 27177 44498
rect 27662 44494 27722 44496
rect 25630 41534 26066 41594
rect 26558 41574 26618 44438
rect 27110 41596 27170 44442
rect 27655 44438 27664 44494
rect 27720 44438 27729 44494
rect 28214 44490 28274 44492
rect 26274 41514 26618 41574
rect 26912 41536 27170 41596
rect 27662 41590 27722 44438
rect 28207 44434 28216 44490
rect 28272 44434 28281 44490
rect 28846 44449 28906 44458
rect 28214 41612 28274 44434
rect 27566 41530 27722 41590
rect 28180 41552 28274 41612
rect 28848 41508 28904 44449
rect 2536 23384 2592 23810
rect 2536 23328 3128 23384
rect 3072 21562 3128 23328
rect 4284 21582 4340 23748
rect 6032 21716 6088 23720
rect 6032 21660 6454 21716
rect 6510 21660 6516 21716
rect 7780 21712 7836 23732
rect 9528 22048 9584 23696
rect 9528 21992 9662 22048
rect 9606 21712 9662 21992
rect 11276 21716 11332 23732
rect 13024 21724 13080 23688
rect 14772 23392 14828 23680
rect 7780 21656 8054 21712
rect 8110 21656 8116 21712
rect 11050 21660 11056 21716
rect 11112 21660 11332 21716
rect 12354 21668 12360 21724
rect 12416 21668 13080 21724
rect 13716 23336 14828 23392
rect 13716 21712 13772 23336
rect 15026 22526 15226 22535
rect 15026 22158 15226 22326
rect 15020 21958 15026 22158
rect 15226 21958 15232 22158
rect 16520 21820 16576 23738
rect 16520 21764 17800 21820
rect 9606 21650 9662 21656
rect 13716 21650 13772 21656
rect 4284 21526 4886 21582
rect 4942 21526 4948 21582
rect 17744 21574 17800 21764
rect 18268 21596 18324 23778
rect 20016 21710 20072 23734
rect 20016 21654 21112 21710
rect 21168 21654 21174 21710
rect 21764 21698 21820 23762
rect 23512 21714 23568 23824
rect 21764 21642 22720 21698
rect 22776 21642 22782 21698
rect 23512 21658 24270 21714
rect 24326 21658 24332 21714
rect 25260 21710 25316 23766
rect 27008 21710 27064 23684
rect 25260 21654 25718 21710
rect 25774 21654 25780 21710
rect 28756 21706 28812 23652
rect 29376 22524 29576 22530
rect 29077 22324 29086 22524
rect 29286 22324 29376 22524
rect 29376 22318 29576 22324
rect 27008 21648 27064 21654
rect 28370 21650 28376 21706
rect 28432 21650 28812 21706
rect 18268 21540 19560 21596
rect 19616 21540 19622 21596
rect 17744 21512 17800 21518
rect 3072 21500 3128 21506
rect 15442 13508 16876 13708
rect 2555 5990 2564 6590
rect 3164 5990 18594 6590
rect 19194 5990 27022 6590
rect 27622 5990 27628 6590
rect 2553 5242 2562 5842
rect 3162 5242 18588 5842
rect 19188 5242 27008 5842
rect 27608 5242 27614 5842
rect 14612 4728 14812 5242
rect 23026 4864 23226 5242
rect 14606 4528 14612 4728
rect 14812 4528 14818 4728
rect 23020 4664 23026 4864
rect 23226 4664 23232 4864
rect 4167 3652 4176 4252
rect 4776 3652 18594 4252
rect 19194 3652 27032 4252
rect 27632 3652 27638 4252
rect 4169 2906 4178 3502
rect 4774 2906 18584 3502
rect 19180 2906 27034 3502
rect 27630 2906 27636 3502
rect 13702 2798 13902 2906
rect 22334 2796 22534 2906
rect 13702 2592 13902 2598
rect 22328 2596 22334 2796
rect 22534 2596 22540 2796
rect 20484 538 20490 738
rect 20690 538 22502 738
rect 22702 538 22711 738
rect 28910 546 28916 746
rect 29116 546 29270 746
rect 29470 546 29479 746
<< via2 >>
rect 2442 44802 2502 44862
rect 3086 44650 3146 44710
rect 3730 44518 3790 44578
rect 4374 44374 4434 44434
rect 17728 44422 17784 44478
rect 18280 44422 18336 44478
rect 18832 44422 18888 44478
rect 19384 44430 19440 44486
rect 19936 44442 19992 44498
rect 20488 44444 20544 44500
rect 5020 44250 5076 44306
rect 5668 44110 5724 44166
rect 6308 43978 6364 44034
rect 6950 43850 7006 43906
rect 7598 43722 7654 43778
rect 8238 43598 8294 43654
rect 8886 43452 8942 43508
rect 9528 43298 9584 43354
rect 10166 43148 10222 43204
rect 10814 43004 10870 43060
rect 11458 42850 11514 42906
rect 12100 42708 12156 42764
rect 12750 42562 12806 42618
rect 13388 42422 13444 42478
rect 14036 42286 14092 42342
rect 14678 41540 14734 41596
rect 15322 41524 15378 41580
rect 21040 44442 21096 44498
rect 21592 44442 21648 44498
rect 22144 44442 22200 44498
rect 22696 44444 22752 44500
rect 23248 44448 23304 44504
rect 23800 44444 23856 44500
rect 24352 44442 24408 44498
rect 24904 44442 24960 44498
rect 25456 44444 25512 44500
rect 26008 44444 26064 44500
rect 26560 44438 26616 44494
rect 27112 44442 27168 44498
rect 27664 44438 27720 44494
rect 28216 44434 28272 44490
rect 28846 44458 28906 44518
rect 15026 22326 15226 22526
rect 29086 22324 29286 22524
rect 2564 5990 3164 6590
rect 2562 5242 3162 5842
rect 4176 3652 4776 4252
rect 4178 2906 4774 3502
rect 22502 538 22702 738
rect 29270 546 29470 746
<< metal3 >>
rect 2437 44862 2507 44867
rect 6128 44862 6134 44864
rect 2437 44802 2442 44862
rect 2502 44802 6134 44862
rect 2437 44797 2507 44802
rect 6128 44800 6134 44802
rect 6198 44800 6204 44864
rect 3081 44710 3151 44715
rect 6674 44710 6680 44712
rect 3081 44650 3086 44710
rect 3146 44650 6680 44710
rect 3081 44645 3151 44650
rect 6674 44648 6680 44650
rect 6744 44648 6750 44712
rect 17718 44622 17724 44686
rect 17788 44622 17794 44686
rect 3725 44578 3795 44583
rect 7220 44578 7226 44580
rect 3725 44518 3730 44578
rect 3790 44518 7226 44578
rect 3725 44513 3795 44518
rect 7220 44516 7226 44518
rect 7290 44516 7296 44580
rect 17726 44483 17786 44622
rect 18270 44620 18276 44684
rect 18340 44620 18346 44684
rect 18822 44620 18828 44684
rect 18892 44620 18898 44684
rect 19374 44630 19380 44694
rect 19444 44630 19450 44694
rect 19926 44638 19932 44702
rect 19996 44638 20002 44702
rect 18278 44483 18338 44620
rect 18830 44483 18890 44620
rect 19382 44491 19442 44630
rect 19934 44503 19994 44638
rect 20478 44634 20484 44698
rect 20548 44634 20554 44698
rect 20486 44505 20546 44634
rect 21030 44630 21036 44694
rect 21100 44630 21106 44694
rect 21582 44634 21588 44698
rect 21652 44634 21658 44698
rect 19931 44498 19997 44503
rect 19379 44486 19445 44491
rect 17723 44478 17789 44483
rect 4369 44434 4439 44439
rect 7778 44434 7784 44436
rect 4369 44374 4374 44434
rect 4434 44374 7784 44434
rect 4369 44369 4439 44374
rect 7778 44372 7784 44374
rect 7848 44372 7854 44436
rect 17723 44422 17728 44478
rect 17784 44422 17789 44478
rect 17723 44417 17789 44422
rect 18275 44478 18341 44483
rect 18275 44422 18280 44478
rect 18336 44422 18341 44478
rect 18275 44417 18341 44422
rect 18827 44478 18893 44483
rect 18827 44422 18832 44478
rect 18888 44422 18893 44478
rect 19379 44430 19384 44486
rect 19440 44430 19445 44486
rect 19931 44442 19936 44498
rect 19992 44442 19997 44498
rect 19931 44437 19997 44442
rect 20483 44500 20549 44505
rect 21038 44503 21098 44630
rect 21590 44503 21650 44634
rect 22134 44630 22140 44694
rect 22204 44630 22210 44694
rect 22142 44503 22202 44630
rect 22686 44620 22692 44684
rect 22756 44620 22762 44684
rect 22694 44505 22754 44620
rect 23238 44616 23244 44680
rect 23308 44616 23314 44680
rect 23790 44616 23796 44680
rect 23860 44616 23866 44680
rect 23246 44509 23306 44616
rect 20483 44444 20488 44500
rect 20544 44444 20549 44500
rect 20483 44439 20549 44444
rect 21035 44498 21101 44503
rect 21035 44442 21040 44498
rect 21096 44442 21101 44498
rect 21035 44437 21101 44442
rect 21587 44498 21653 44503
rect 21587 44442 21592 44498
rect 21648 44442 21653 44498
rect 21587 44437 21653 44442
rect 22139 44498 22205 44503
rect 22139 44442 22144 44498
rect 22200 44442 22205 44498
rect 22139 44437 22205 44442
rect 22691 44500 22757 44505
rect 22691 44444 22696 44500
rect 22752 44444 22757 44500
rect 22691 44439 22757 44444
rect 23243 44504 23309 44509
rect 23798 44505 23858 44616
rect 24342 44608 24348 44672
rect 24412 44608 24418 44672
rect 23243 44448 23248 44504
rect 23304 44448 23309 44504
rect 23243 44443 23309 44448
rect 23795 44500 23861 44505
rect 24350 44503 24410 44608
rect 24894 44602 24900 44666
rect 24964 44602 24970 44666
rect 25446 44608 25452 44672
rect 25516 44608 25522 44672
rect 25998 44608 26004 44672
rect 26068 44608 26074 44672
rect 24902 44503 24962 44602
rect 25454 44505 25514 44608
rect 26006 44505 26066 44608
rect 26550 44602 26556 44666
rect 26620 44602 26626 44666
rect 23795 44444 23800 44500
rect 23856 44444 23861 44500
rect 23795 44439 23861 44444
rect 24347 44498 24413 44503
rect 24347 44442 24352 44498
rect 24408 44442 24413 44498
rect 24347 44437 24413 44442
rect 24899 44498 24965 44503
rect 24899 44442 24904 44498
rect 24960 44442 24965 44498
rect 24899 44437 24965 44442
rect 25451 44500 25517 44505
rect 25451 44444 25456 44500
rect 25512 44444 25517 44500
rect 25451 44439 25517 44444
rect 26003 44500 26069 44505
rect 26003 44444 26008 44500
rect 26064 44444 26069 44500
rect 26558 44499 26618 44602
rect 27102 44598 27108 44662
rect 27172 44598 27178 44662
rect 27110 44503 27170 44598
rect 27654 44594 27660 44658
rect 27724 44594 27730 44658
rect 28206 44598 28212 44662
rect 28276 44598 28282 44662
rect 28844 44656 28908 44662
rect 26003 44439 26069 44444
rect 26555 44494 26621 44499
rect 26555 44438 26560 44494
rect 26616 44438 26621 44494
rect 26555 44433 26621 44438
rect 27107 44498 27173 44503
rect 27662 44499 27722 44594
rect 27107 44442 27112 44498
rect 27168 44442 27173 44498
rect 27107 44437 27173 44442
rect 27659 44494 27725 44499
rect 28214 44495 28274 44598
rect 28844 44586 28908 44592
rect 28846 44523 28906 44586
rect 28841 44518 28911 44523
rect 27659 44438 27664 44494
rect 27720 44438 27725 44494
rect 27659 44433 27725 44438
rect 28211 44490 28277 44495
rect 28211 44434 28216 44490
rect 28272 44434 28277 44490
rect 28841 44458 28846 44518
rect 28906 44458 28911 44518
rect 28841 44453 28911 44458
rect 19379 44425 19445 44430
rect 28211 44429 28277 44434
rect 18827 44417 18893 44422
rect 5015 44308 5081 44311
rect 8334 44308 8340 44310
rect 5015 44306 8340 44308
rect 5015 44250 5020 44306
rect 5076 44250 8340 44306
rect 5015 44248 8340 44250
rect 5015 44245 5081 44248
rect 8334 44246 8340 44248
rect 8404 44246 8410 44310
rect 5663 44168 5729 44171
rect 8886 44168 8892 44170
rect 5663 44166 8892 44168
rect 5663 44110 5668 44166
rect 5724 44110 8892 44166
rect 5663 44108 8892 44110
rect 5663 44105 5729 44108
rect 8886 44106 8892 44108
rect 8956 44106 8962 44170
rect 6303 44036 6369 44039
rect 9438 44036 9444 44038
rect 6303 44034 9444 44036
rect 6303 43978 6308 44034
rect 6364 43978 9444 44034
rect 6303 43976 9444 43978
rect 6303 43973 6369 43976
rect 9438 43974 9444 43976
rect 9508 43974 9514 44038
rect 6945 43908 7011 43911
rect 9990 43908 9996 43910
rect 6945 43906 9996 43908
rect 6945 43850 6950 43906
rect 7006 43850 9996 43906
rect 6945 43848 9996 43850
rect 6945 43845 7011 43848
rect 9990 43846 9996 43848
rect 10060 43846 10066 43910
rect 7593 43780 7659 43783
rect 10542 43780 10548 43782
rect 7593 43778 10548 43780
rect 7593 43722 7598 43778
rect 7654 43722 10548 43778
rect 7593 43720 10548 43722
rect 7593 43717 7659 43720
rect 10542 43718 10548 43720
rect 10612 43718 10618 43782
rect 8233 43656 8299 43659
rect 11094 43656 11100 43658
rect 8233 43654 11100 43656
rect 8233 43598 8238 43654
rect 8294 43598 11100 43654
rect 8233 43596 11100 43598
rect 8233 43593 8299 43596
rect 11094 43594 11100 43596
rect 11164 43594 11170 43658
rect 8881 43510 8947 43513
rect 11646 43510 11652 43512
rect 8881 43508 11652 43510
rect 8881 43452 8886 43508
rect 8942 43452 11652 43508
rect 8881 43450 11652 43452
rect 8881 43447 8947 43450
rect 11646 43448 11652 43450
rect 11716 43448 11722 43512
rect 9523 43356 9589 43359
rect 12198 43356 12204 43358
rect 9523 43354 12204 43356
rect 9523 43298 9528 43354
rect 9584 43298 12204 43354
rect 9523 43296 12204 43298
rect 9523 43293 9589 43296
rect 12198 43294 12204 43296
rect 12268 43294 12274 43358
rect 10161 43206 10227 43209
rect 12750 43206 12756 43208
rect 10161 43204 12756 43206
rect 10161 43148 10166 43204
rect 10222 43148 12756 43204
rect 10161 43146 12756 43148
rect 10161 43143 10227 43146
rect 12750 43144 12756 43146
rect 12820 43144 12826 43208
rect 10809 43062 10875 43065
rect 13302 43062 13308 43064
rect 10809 43060 13308 43062
rect 10809 43004 10814 43060
rect 10870 43004 13308 43060
rect 10809 43002 13308 43004
rect 10809 42999 10875 43002
rect 13302 43000 13308 43002
rect 13372 43000 13378 43064
rect 11453 42908 11519 42911
rect 13854 42908 13860 42910
rect 11453 42906 13860 42908
rect 11453 42850 11458 42906
rect 11514 42850 13860 42906
rect 11453 42848 13860 42850
rect 11453 42845 11519 42848
rect 13854 42846 13860 42848
rect 13924 42846 13930 42910
rect 12095 42766 12161 42769
rect 14406 42766 14412 42768
rect 12095 42764 14412 42766
rect 12095 42708 12100 42764
rect 12156 42708 14412 42764
rect 12095 42706 14412 42708
rect 12095 42703 12161 42706
rect 14406 42704 14412 42706
rect 14476 42704 14482 42768
rect 12745 42620 12811 42623
rect 14958 42620 14964 42622
rect 12745 42618 14964 42620
rect 12745 42562 12750 42618
rect 12806 42562 14964 42618
rect 12745 42560 14964 42562
rect 12745 42557 12811 42560
rect 14958 42558 14964 42560
rect 15028 42558 15034 42622
rect 13383 42480 13449 42483
rect 15510 42480 15516 42482
rect 13383 42478 15516 42480
rect 13383 42422 13388 42478
rect 13444 42422 15516 42478
rect 13383 42420 15516 42422
rect 13383 42417 13449 42420
rect 15510 42418 15516 42420
rect 15580 42418 15586 42482
rect 14031 42344 14097 42347
rect 15740 42344 15746 42346
rect 14031 42342 15746 42344
rect 14031 42286 14036 42342
rect 14092 42286 15746 42342
rect 14031 42284 15746 42286
rect 14031 42281 14097 42284
rect 15740 42282 15746 42284
rect 15810 42282 15816 42346
rect 14674 42164 14738 42170
rect 14674 42094 14738 42100
rect 14676 41601 14736 42094
rect 15318 41882 15382 41888
rect 15318 41812 15382 41818
rect 14673 41596 14739 41601
rect 14673 41540 14678 41596
rect 14734 41540 14739 41596
rect 15320 41585 15380 41812
rect 14673 41535 14739 41540
rect 15317 41580 15383 41585
rect 15317 41524 15322 41580
rect 15378 41524 15383 41580
rect 15317 41519 15383 41524
rect 5441 23964 5759 23965
rect 5436 23648 5442 23964
rect 5758 23648 5764 23964
rect 18872 23863 19192 23864
rect 12156 23773 12476 23774
rect 5441 22604 5759 23648
rect 12151 23455 12157 23773
rect 12475 23455 12481 23773
rect 18867 23545 18873 23863
rect 19191 23545 19197 23863
rect 25588 23739 25908 23740
rect 12156 22604 12476 23455
rect 18872 22606 19192 23545
rect 25583 23421 25589 23739
rect 25907 23421 25913 23739
rect 25588 22606 25908 23421
rect 18872 22604 25908 22606
rect 5441 22591 25908 22604
rect 205 22273 211 22591
rect 529 22526 25908 22591
rect 529 22326 15026 22526
rect 15226 22524 25908 22526
rect 29081 22524 29291 22529
rect 15226 22326 29086 22524
rect 529 22324 29086 22326
rect 29286 22324 29291 22524
rect 529 22286 25908 22324
rect 29081 22319 29291 22324
rect 529 22284 19192 22286
rect 529 22273 5759 22284
rect 2559 6590 3169 6595
rect 216 6584 2564 6590
rect 216 5996 222 6584
rect 594 5996 2564 6584
rect 216 5990 2564 5996
rect 3164 5990 3169 6590
rect 2559 5985 3169 5990
rect 2557 5842 3167 5847
rect 210 5836 2562 5842
rect 210 5248 216 5836
rect 594 5248 2562 5836
rect 210 5242 2562 5248
rect 3162 5242 3167 5842
rect 2557 5237 3167 5242
rect 4171 4252 4781 4257
rect 3206 3652 3212 4252
rect 3812 3652 4176 4252
rect 4776 3652 4781 4252
rect 4171 3647 4781 3652
rect 4173 3502 4779 3507
rect 3186 2906 3192 3502
rect 3788 2906 4178 3502
rect 4774 2906 4779 3502
rect 4173 2901 4779 2906
rect 29265 746 29475 751
rect 22497 738 22707 743
rect 22497 538 22502 738
rect 22702 538 24722 738
rect 24922 538 24928 738
rect 29265 546 29270 746
rect 29470 546 29682 746
rect 29882 546 29888 746
rect 29265 541 29475 546
rect 22497 533 22707 538
<< via3 >>
rect 6134 44800 6198 44864
rect 6680 44648 6744 44712
rect 17724 44622 17788 44686
rect 7226 44516 7290 44580
rect 18276 44620 18340 44684
rect 18828 44620 18892 44684
rect 19380 44630 19444 44694
rect 19932 44638 19996 44702
rect 20484 44634 20548 44698
rect 21036 44630 21100 44694
rect 21588 44634 21652 44698
rect 7784 44372 7848 44436
rect 22140 44630 22204 44694
rect 22692 44620 22756 44684
rect 23244 44616 23308 44680
rect 23796 44616 23860 44680
rect 24348 44608 24412 44672
rect 24900 44602 24964 44666
rect 25452 44608 25516 44672
rect 26004 44608 26068 44672
rect 26556 44602 26620 44666
rect 27108 44598 27172 44662
rect 27660 44594 27724 44658
rect 28212 44598 28276 44662
rect 28844 44592 28908 44656
rect 8340 44246 8404 44310
rect 8892 44106 8956 44170
rect 9444 43974 9508 44038
rect 9996 43846 10060 43910
rect 10548 43718 10612 43782
rect 11100 43594 11164 43658
rect 11652 43448 11716 43512
rect 12204 43294 12268 43358
rect 12756 43144 12820 43208
rect 13308 43000 13372 43064
rect 13860 42846 13924 42910
rect 14412 42704 14476 42768
rect 14964 42558 15028 42622
rect 15516 42418 15580 42482
rect 15746 42282 15810 42346
rect 14674 42100 14738 42164
rect 15318 41818 15382 41882
rect 5442 23648 5758 23964
rect 12157 23455 12475 23773
rect 18873 23545 19191 23863
rect 25589 23421 25907 23739
rect 211 22273 529 22591
rect 222 5996 594 6584
rect 216 5248 594 5836
rect 3212 3652 3812 4252
rect 3192 2906 3788 3502
rect 24722 538 24922 738
rect 29682 546 29882 746
<< metal4 >>
rect 6134 45030 6194 45152
rect 6134 44952 6196 45030
rect 6686 45024 6746 45152
rect 7238 45042 7298 45152
rect 6136 44865 6196 44952
rect 6682 44952 6746 45024
rect 7228 44952 7298 45042
rect 7790 45012 7850 45152
rect 7786 44952 7850 45012
rect 6133 44864 6199 44865
rect 6133 44800 6134 44864
rect 6198 44800 6199 44864
rect 6133 44799 6199 44800
rect 6682 44713 6742 44952
rect 6679 44712 6745 44713
rect 6679 44648 6680 44712
rect 6744 44648 6745 44712
rect 6679 44647 6745 44648
rect 7228 44581 7288 44952
rect 7225 44580 7291 44581
rect 7225 44516 7226 44580
rect 7290 44516 7291 44580
rect 7225 44515 7291 44516
rect 7786 44437 7846 44952
rect 7783 44436 7849 44437
rect 7783 44372 7784 44436
rect 7848 44372 7849 44436
rect 7783 44371 7849 44372
rect 8342 44311 8402 45152
rect 8339 44310 8405 44311
rect 8339 44246 8340 44310
rect 8404 44246 8405 44310
rect 8339 44245 8405 44246
rect 8894 44171 8954 45152
rect 8891 44170 8957 44171
rect 200 22591 600 44152
rect 200 22273 211 22591
rect 529 22273 600 22591
rect 200 6584 600 22273
rect 200 5996 222 6584
rect 594 5996 600 6584
rect 200 5836 600 5996
rect 200 5248 216 5836
rect 594 5248 600 5836
rect 200 1000 600 5248
rect 800 23122 1200 44152
rect 8891 44106 8892 44170
rect 8956 44106 8957 44170
rect 8891 44105 8957 44106
rect 9446 44039 9506 45152
rect 9443 44038 9509 44039
rect 9443 43974 9444 44038
rect 9508 43974 9509 44038
rect 9443 43973 9509 43974
rect 9998 43911 10058 45152
rect 9995 43910 10061 43911
rect 9995 43846 9996 43910
rect 10060 43846 10061 43910
rect 9995 43845 10061 43846
rect 10550 43783 10610 45152
rect 10547 43782 10613 43783
rect 10547 43718 10548 43782
rect 10612 43718 10613 43782
rect 10547 43717 10613 43718
rect 11102 43659 11162 45152
rect 11099 43658 11165 43659
rect 11099 43594 11100 43658
rect 11164 43594 11165 43658
rect 11099 43593 11165 43594
rect 11654 43513 11714 45152
rect 11651 43512 11717 43513
rect 11651 43448 11652 43512
rect 11716 43448 11717 43512
rect 11651 43447 11717 43448
rect 12206 43359 12266 45152
rect 12203 43358 12269 43359
rect 12203 43294 12204 43358
rect 12268 43294 12269 43358
rect 12203 43293 12269 43294
rect 12758 43209 12818 45152
rect 12755 43208 12821 43209
rect 12755 43144 12756 43208
rect 12820 43144 12821 43208
rect 12755 43143 12821 43144
rect 13310 43065 13370 45152
rect 13307 43064 13373 43065
rect 13307 43000 13308 43064
rect 13372 43000 13373 43064
rect 13307 42999 13373 43000
rect 13862 42911 13922 45152
rect 13859 42910 13925 42911
rect 13859 42846 13860 42910
rect 13924 42846 13925 42910
rect 13859 42845 13925 42846
rect 14414 42769 14474 45152
rect 14411 42768 14477 42769
rect 14411 42704 14412 42768
rect 14476 42704 14477 42768
rect 14411 42703 14477 42704
rect 14966 42623 15026 45152
rect 14963 42622 15029 42623
rect 14963 42558 14964 42622
rect 15028 42558 15029 42622
rect 14963 42557 15029 42558
rect 15518 42483 15578 45152
rect 16070 44662 16130 45152
rect 15748 44602 16130 44662
rect 15515 42482 15581 42483
rect 15515 42418 15516 42482
rect 15580 42418 15581 42482
rect 15515 42417 15581 42418
rect 15748 42347 15808 44602
rect 16622 44476 16682 45152
rect 17174 44648 17234 45152
rect 17726 44687 17786 45152
rect 16266 44416 16682 44476
rect 16958 44588 17234 44648
rect 17723 44686 17789 44687
rect 17723 44622 17724 44686
rect 17788 44622 17789 44686
rect 18278 44685 18338 45152
rect 18830 44685 18890 45152
rect 19382 44695 19442 45152
rect 19934 44703 19994 45152
rect 19931 44702 19997 44703
rect 19379 44694 19445 44695
rect 17723 44621 17789 44622
rect 18275 44684 18341 44685
rect 18275 44620 18276 44684
rect 18340 44620 18341 44684
rect 18275 44619 18341 44620
rect 18827 44684 18893 44685
rect 18827 44620 18828 44684
rect 18892 44620 18893 44684
rect 19379 44630 19380 44694
rect 19444 44630 19445 44694
rect 19931 44638 19932 44702
rect 19996 44638 19997 44702
rect 20486 44699 20546 45152
rect 19931 44637 19997 44638
rect 20483 44698 20549 44699
rect 20483 44634 20484 44698
rect 20548 44634 20549 44698
rect 21038 44695 21098 45152
rect 21590 44699 21650 45152
rect 21587 44698 21653 44699
rect 20483 44633 20549 44634
rect 21035 44694 21101 44695
rect 19379 44629 19445 44630
rect 21035 44630 21036 44694
rect 21100 44630 21101 44694
rect 21587 44634 21588 44698
rect 21652 44634 21653 44698
rect 22142 44695 22202 45152
rect 21587 44633 21653 44634
rect 22139 44694 22205 44695
rect 21035 44629 21101 44630
rect 22139 44630 22140 44694
rect 22204 44630 22205 44694
rect 22694 44685 22754 45152
rect 22139 44629 22205 44630
rect 22691 44684 22757 44685
rect 18827 44619 18893 44620
rect 22691 44620 22692 44684
rect 22756 44620 22757 44684
rect 23246 44681 23306 45152
rect 23798 44681 23858 45152
rect 22691 44619 22757 44620
rect 23243 44680 23309 44681
rect 23243 44616 23244 44680
rect 23308 44616 23309 44680
rect 23243 44615 23309 44616
rect 23795 44680 23861 44681
rect 23795 44616 23796 44680
rect 23860 44616 23861 44680
rect 24350 44673 24410 45152
rect 23795 44615 23861 44616
rect 24347 44672 24413 44673
rect 24347 44608 24348 44672
rect 24412 44608 24413 44672
rect 24902 44667 24962 45152
rect 25454 44673 25514 45152
rect 26006 44673 26066 45152
rect 25451 44672 25517 44673
rect 24347 44607 24413 44608
rect 24899 44666 24965 44667
rect 24899 44602 24900 44666
rect 24964 44602 24965 44666
rect 25451 44608 25452 44672
rect 25516 44608 25517 44672
rect 25451 44607 25517 44608
rect 26003 44672 26069 44673
rect 26003 44608 26004 44672
rect 26068 44608 26069 44672
rect 26558 44667 26618 45152
rect 26003 44607 26069 44608
rect 26555 44666 26621 44667
rect 24899 44601 24965 44602
rect 26555 44602 26556 44666
rect 26620 44602 26621 44666
rect 27110 44663 27170 45152
rect 26555 44601 26621 44602
rect 27107 44662 27173 44663
rect 27107 44598 27108 44662
rect 27172 44598 27173 44662
rect 27662 44659 27722 45152
rect 28214 44663 28274 45152
rect 28766 45012 28826 45152
rect 28766 44952 28830 45012
rect 29318 44952 29378 45152
rect 28770 44858 28830 44952
rect 28770 44798 28906 44858
rect 28211 44662 28277 44663
rect 27107 44597 27173 44598
rect 27659 44658 27725 44659
rect 27659 44594 27660 44658
rect 27724 44594 27725 44658
rect 28211 44598 28212 44662
rect 28276 44598 28277 44662
rect 28846 44657 28906 44798
rect 28211 44597 28277 44598
rect 28843 44656 28909 44657
rect 27659 44593 27725 44594
rect 28843 44592 28844 44656
rect 28908 44592 28909 44656
rect 28843 44591 28909 44592
rect 15745 42346 15811 42347
rect 15745 42282 15746 42346
rect 15810 42282 15811 42346
rect 15745 42281 15811 42282
rect 14673 42164 14739 42165
rect 14673 42100 14674 42164
rect 14738 42162 14739 42164
rect 16266 42162 16326 44416
rect 14738 42102 16326 42162
rect 14738 42100 14739 42102
rect 14673 42099 14739 42100
rect 15317 41882 15383 41883
rect 15317 41818 15318 41882
rect 15382 41880 15383 41882
rect 16958 41880 17018 44588
rect 15382 41820 17018 41880
rect 15382 41818 15383 41820
rect 15317 41817 15383 41818
rect 5441 23964 5759 24526
rect 5441 23648 5442 23964
rect 5758 23648 5759 23964
rect 5441 23647 5759 23648
rect 8798 23122 9118 24496
rect 12156 23773 12476 24524
rect 12156 23455 12157 23773
rect 12475 23455 12476 23773
rect 12156 23454 12476 23455
rect 15514 23122 15834 24492
rect 18872 23863 19192 24582
rect 18872 23545 18873 23863
rect 19191 23545 19192 23863
rect 18872 23544 19192 23545
rect 22230 23122 22550 24490
rect 25588 23739 25908 24484
rect 25588 23421 25589 23739
rect 25907 23421 25908 23739
rect 25588 23420 25908 23421
rect 28946 23122 29266 24490
rect 800 22802 29266 23122
rect 800 4252 1200 22802
rect 3211 4252 3813 4253
rect 800 3652 3212 4252
rect 3812 3652 3813 4252
rect 800 3502 1200 3652
rect 3211 3651 3813 3652
rect 3191 3502 3789 3503
rect 800 2906 3192 3502
rect 3788 2906 3789 3502
rect 800 1000 1200 2906
rect 3191 2905 3789 2906
rect 29681 746 29883 747
rect 24721 738 24923 739
rect 24721 538 24722 738
rect 24922 538 26682 738
rect 29681 546 29682 746
rect 29882 730 29883 746
rect 29882 550 30542 730
rect 29882 546 29883 550
rect 29681 545 29883 546
rect 24721 537 24923 538
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 538
rect 30362 0 30542 550
use buffer  buffer_0
timestamp 1740347555
transform 1 0 23012 0 1 2996
box 14 -2066 6984 8200
use buffer  buffer_2
timestamp 1740347555
transform 1 0 14586 0 1 2998
box 14 -2066 6984 8200
use dac  dac_1
timestamp 1740347555
transform 1 0 23086 0 1 13038
box -6918 -1472 7384 8872
use dac  dac_2
timestamp 1740347555
transform 1 0 8418 0 1 13038
box -6918 -1472 7384 8872
use digital_top  digital_top_0
timestamp 1757770450
transform 1 0 1690 0 1 23594
box 514 0 27576 18000
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
