magic
tech sky130A
magscale 1 2
timestamp 1757869722
<< viali >>
rect 857 17289 891 17323
rect 1501 17289 1535 17323
rect 4077 17289 4111 17323
rect 6009 17289 6043 17323
rect 6653 17289 6687 17323
rect 8125 17289 8159 17323
rect 9229 17289 9263 17323
rect 10609 17289 10643 17323
rect 12081 17289 12115 17323
rect 14197 17289 14231 17323
rect 22753 17289 22787 17323
rect 24685 17289 24719 17323
rect 25145 17289 25179 17323
rect 18337 17221 18371 17255
rect 23397 17221 23431 17255
rect 24041 17221 24075 17255
rect 2789 17153 2823 17187
rect 3433 17153 3467 17187
rect 4721 17153 4755 17187
rect 5365 17153 5399 17187
rect 19717 17153 19751 17187
rect 20269 17153 20303 17187
rect 21741 17153 21775 17187
rect 21833 17153 21867 17187
rect 25421 17153 25455 17187
rect 7941 17085 7975 17119
rect 10149 17085 10183 17119
rect 10793 17085 10827 17119
rect 11897 17085 11931 17119
rect 14381 17085 14415 17119
rect 16497 17085 16531 17119
rect 16957 17085 16991 17119
rect 17785 17085 17819 17119
rect 18521 17085 18555 17119
rect 18981 17085 19015 17119
rect 19073 17085 19107 17119
rect 19533 17085 19567 17119
rect 20085 17085 20119 17119
rect 20637 17085 20671 17119
rect 20729 17085 20763 17119
rect 21097 17085 21131 17119
rect 21557 17085 21591 17119
rect 22017 17085 22051 17119
rect 22569 17085 22603 17119
rect 22937 17085 22971 17119
rect 23581 17085 23615 17119
rect 24225 17085 24259 17119
rect 24869 17085 24903 17119
rect 25329 17085 25363 17119
rect 25697 17085 25731 17119
rect 26433 17085 26467 17119
rect 22201 17017 22235 17051
rect 9597 16949 9631 16983
rect 16313 16949 16347 16983
rect 17141 16949 17175 16983
rect 17601 16949 17635 16983
rect 18797 16949 18831 16983
rect 19349 16949 19383 16983
rect 19901 16949 19935 16983
rect 20453 16949 20487 16983
rect 20913 16949 20947 16983
rect 21373 16949 21407 16983
rect 22385 16949 22419 16983
rect 27077 16949 27111 16983
rect 7941 16745 7975 16779
rect 9781 16745 9815 16779
rect 10977 16745 11011 16779
rect 12817 16745 12851 16779
rect 13645 16745 13679 16779
rect 15485 16745 15519 16779
rect 15853 16745 15887 16779
rect 6736 16677 6770 16711
rect 13093 16677 13127 16711
rect 13461 16677 13495 16711
rect 14841 16677 14875 16711
rect 15025 16677 15059 16711
rect 19257 16677 19291 16711
rect 24777 16677 24811 16711
rect 26433 16677 26467 16711
rect 8125 16609 8159 16643
rect 8217 16609 8251 16643
rect 8484 16609 8518 16643
rect 9965 16609 9999 16643
rect 10793 16609 10827 16643
rect 12090 16609 12124 16643
rect 12357 16609 12391 16643
rect 13001 16609 13035 16643
rect 14013 16609 14047 16643
rect 14105 16609 14139 16643
rect 15301 16609 15335 16643
rect 15669 16609 15703 16643
rect 16589 16609 16623 16643
rect 16773 16609 16807 16643
rect 19533 16609 19567 16643
rect 19625 16609 19659 16643
rect 19717 16609 19751 16643
rect 19901 16609 19935 16643
rect 22109 16609 22143 16643
rect 22477 16609 22511 16643
rect 22569 16609 22603 16643
rect 22661 16609 22695 16643
rect 22845 16609 22879 16643
rect 24133 16609 24167 16643
rect 24317 16609 24351 16643
rect 24409 16609 24443 16643
rect 24501 16609 24535 16643
rect 25513 16609 25547 16643
rect 26249 16609 26283 16643
rect 26709 16609 26743 16643
rect 26801 16609 26835 16643
rect 26893 16609 26927 16643
rect 27077 16609 27111 16643
rect 6469 16541 6503 16575
rect 14197 16541 14231 16575
rect 15117 16541 15151 16575
rect 16957 16541 16991 16575
rect 18521 16541 18555 16575
rect 20637 16541 20671 16575
rect 22201 16541 22235 16575
rect 23489 16541 23523 16575
rect 9597 16473 9631 16507
rect 19993 16473 20027 16507
rect 22937 16473 22971 16507
rect 7849 16405 7883 16439
rect 10149 16405 10183 16439
rect 14565 16405 14599 16439
rect 19073 16405 19107 16439
rect 21465 16405 21499 16439
rect 24961 16405 24995 16439
rect 26065 16405 26099 16439
rect 7113 16201 7147 16235
rect 8493 16201 8527 16235
rect 10149 16201 10183 16235
rect 10333 16201 10367 16235
rect 11529 16201 11563 16235
rect 12081 16201 12115 16235
rect 14473 16201 14507 16235
rect 22569 16201 22603 16235
rect 25329 16201 25363 16235
rect 6469 16133 6503 16167
rect 10057 16133 10091 16167
rect 10977 16133 11011 16167
rect 13369 16133 13403 16167
rect 22477 16133 22511 16167
rect 9229 16065 9263 16099
rect 10517 16065 10551 16099
rect 11161 16065 11195 16099
rect 20729 16065 20763 16099
rect 6929 15997 6963 16031
rect 8769 15997 8803 16031
rect 8861 15997 8895 16031
rect 8953 15997 8987 16031
rect 9137 15997 9171 16031
rect 9413 15997 9447 16031
rect 9689 15997 9723 16031
rect 9781 15997 9815 16031
rect 10057 15997 10091 16031
rect 10333 15997 10367 16031
rect 10885 15997 10919 16031
rect 11713 15997 11747 16031
rect 12265 15997 12299 16031
rect 12449 15997 12483 16031
rect 13185 15997 13219 16031
rect 13369 15997 13403 16031
rect 14197 15997 14231 16031
rect 14657 15997 14691 16031
rect 15117 15997 15151 16031
rect 17233 15997 17267 16031
rect 18705 15997 18739 16031
rect 21097 15997 21131 16031
rect 21364 15997 21398 16031
rect 22707 15997 22741 16031
rect 22845 15997 22879 16031
rect 23120 15997 23154 16031
rect 23213 15997 23247 16031
rect 23397 15997 23431 16031
rect 23489 15997 23523 16031
rect 25237 15997 25271 16031
rect 25881 15997 25915 16031
rect 26249 15997 26283 16031
rect 6837 15929 6871 15963
rect 7665 15929 7699 15963
rect 7849 15929 7883 15963
rect 10793 15929 10827 15963
rect 11161 15929 11195 15963
rect 13553 15929 13587 15963
rect 18972 15929 19006 15963
rect 20177 15929 20211 15963
rect 22937 15929 22971 15963
rect 24970 15929 25004 15963
rect 6377 15861 6411 15895
rect 9597 15861 9631 15895
rect 9873 15861 9907 15895
rect 13093 15861 13127 15895
rect 15301 15861 15335 15895
rect 17877 15861 17911 15895
rect 20085 15861 20119 15895
rect 23857 15861 23891 15895
rect 26801 15861 26835 15895
rect 8769 15657 8803 15691
rect 12081 15657 12115 15691
rect 18613 15657 18647 15691
rect 22109 15657 22143 15691
rect 27077 15657 27111 15691
rect 10701 15589 10735 15623
rect 11069 15589 11103 15623
rect 12808 15589 12842 15623
rect 19441 15589 19475 15623
rect 22477 15589 22511 15623
rect 25136 15589 25170 15623
rect 5365 15521 5399 15555
rect 5549 15521 5583 15555
rect 5825 15521 5859 15555
rect 6092 15521 6126 15555
rect 8585 15521 8619 15555
rect 8769 15521 8803 15555
rect 10609 15521 10643 15555
rect 10977 15521 11011 15555
rect 11253 15521 11287 15555
rect 11713 15521 11747 15555
rect 11805 15521 11839 15555
rect 12541 15521 12575 15555
rect 17233 15521 17267 15555
rect 17500 15521 17534 15555
rect 18705 15521 18739 15555
rect 18889 15521 18923 15555
rect 18981 15521 19015 15555
rect 19073 15521 19107 15555
rect 22247 15521 22281 15555
rect 22385 15521 22419 15555
rect 22660 15521 22694 15555
rect 22753 15521 22787 15555
rect 22845 15521 22879 15555
rect 23029 15521 23063 15555
rect 23121 15521 23155 15555
rect 23213 15521 23247 15555
rect 23581 15521 23615 15555
rect 26433 15521 26467 15555
rect 26581 15521 26615 15555
rect 26709 15521 26743 15555
rect 26801 15521 26835 15555
rect 26898 15521 26932 15555
rect 5641 15453 5675 15487
rect 11621 15453 11655 15487
rect 11897 15453 11931 15487
rect 14749 15453 14783 15487
rect 19349 15453 19383 15487
rect 19993 15453 20027 15487
rect 20177 15453 20211 15487
rect 21373 15453 21407 15487
rect 24225 15453 24259 15487
rect 24869 15453 24903 15487
rect 7205 15385 7239 15419
rect 13921 15385 13955 15419
rect 5181 15317 5215 15351
rect 11437 15317 11471 15351
rect 14105 15317 14139 15351
rect 20821 15317 20855 15351
rect 22017 15317 22051 15351
rect 23489 15317 23523 15351
rect 26249 15317 26283 15351
rect 6469 15113 6503 15147
rect 7481 15113 7515 15147
rect 10425 15113 10459 15147
rect 10885 15113 10919 15147
rect 11253 15113 11287 15147
rect 15485 15113 15519 15147
rect 17049 15113 17083 15147
rect 20177 15113 20211 15147
rect 25237 15113 25271 15147
rect 9689 15045 9723 15079
rect 9873 15045 9907 15079
rect 10609 15045 10643 15079
rect 18245 15045 18279 15079
rect 2973 14977 3007 15011
rect 7113 14977 7147 15011
rect 7665 14977 7699 15011
rect 8125 14977 8159 15011
rect 21189 14977 21223 15011
rect 23857 14977 23891 15011
rect 26341 14977 26375 15011
rect 26985 14977 27019 15011
rect 2789 14909 2823 14943
rect 3065 14909 3099 14943
rect 3893 14909 3927 14943
rect 5089 14909 5123 14943
rect 7481 14909 7515 14943
rect 8033 14909 8067 14943
rect 8217 14909 8251 14943
rect 9505 14909 9539 14943
rect 9781 14909 9815 14943
rect 10057 14909 10091 14943
rect 10149 14909 10183 14943
rect 11345 14909 11379 14943
rect 11621 14909 11655 14943
rect 11805 14909 11839 14943
rect 11989 14909 12023 14943
rect 14105 14909 14139 14943
rect 15669 14909 15703 14943
rect 17601 14909 17635 14943
rect 17749 14909 17783 14943
rect 18107 14909 18141 14943
rect 18981 14909 19015 14943
rect 19073 14909 19107 14943
rect 19165 14909 19199 14943
rect 19349 14909 19383 14943
rect 20085 14909 20119 14943
rect 20356 14909 20390 14943
rect 20453 14909 20487 14943
rect 20728 14909 20762 14943
rect 20821 14909 20855 14943
rect 23213 14909 23247 14943
rect 25697 14909 25731 14943
rect 25881 14909 25915 14943
rect 25973 14909 26007 14943
rect 26065 14909 26099 14943
rect 3249 14841 3283 14875
rect 5334 14841 5368 14875
rect 7941 14841 7975 14875
rect 9873 14841 9907 14875
rect 10241 14841 10275 14875
rect 11069 14841 11103 14875
rect 11713 14841 11747 14875
rect 12234 14841 12268 14875
rect 14372 14841 14406 14875
rect 15936 14841 15970 14875
rect 17877 14841 17911 14875
rect 17969 14841 18003 14875
rect 20545 14841 20579 14875
rect 21456 14841 21490 14875
rect 22661 14841 22695 14875
rect 24102 14841 24136 14875
rect 2605 14773 2639 14807
rect 6561 14773 6595 14807
rect 7297 14773 7331 14807
rect 9321 14773 9355 14807
rect 10451 14773 10485 14807
rect 10701 14773 10735 14807
rect 10869 14773 10903 14807
rect 13369 14773 13403 14807
rect 18705 14773 18739 14807
rect 19441 14773 19475 14807
rect 22569 14773 22603 14807
rect 26433 14773 26467 14807
rect 3801 14569 3835 14603
rect 6377 14569 6411 14603
rect 10701 14569 10735 14603
rect 11529 14569 11563 14603
rect 13829 14569 13863 14603
rect 17049 14569 17083 14603
rect 19717 14569 19751 14603
rect 21281 14569 21315 14603
rect 22753 14569 22787 14603
rect 26249 14569 26283 14603
rect 27077 14569 27111 14603
rect 6009 14501 6043 14535
rect 7465 14501 7499 14535
rect 7665 14501 7699 14535
rect 11989 14501 12023 14535
rect 18604 14501 18638 14535
rect 25136 14501 25170 14535
rect 2053 14433 2087 14467
rect 2329 14433 2363 14467
rect 2688 14433 2722 14467
rect 4445 14433 4479 14467
rect 5181 14433 5215 14467
rect 6561 14433 6595 14467
rect 6745 14433 6779 14467
rect 6837 14433 6871 14467
rect 8401 14433 8435 14467
rect 8493 14433 8527 14467
rect 8769 14433 8803 14467
rect 9045 14433 9079 14467
rect 9505 14433 9539 14467
rect 10149 14431 10183 14465
rect 10333 14423 10367 14457
rect 10609 14433 10643 14467
rect 10793 14433 10827 14467
rect 11161 14433 11195 14467
rect 11345 14433 11379 14467
rect 11897 14433 11931 14467
rect 13369 14433 13403 14467
rect 13553 14433 13587 14467
rect 14105 14433 14139 14467
rect 14197 14433 14231 14467
rect 14289 14433 14323 14467
rect 14473 14433 14507 14467
rect 14565 14433 14599 14467
rect 14749 14433 14783 14467
rect 14841 14433 14875 14467
rect 14933 14433 14967 14467
rect 16129 14433 16163 14467
rect 16865 14433 16899 14467
rect 18337 14433 18371 14467
rect 20545 14433 20579 14467
rect 22394 14433 22428 14467
rect 23029 14433 23063 14467
rect 23121 14433 23155 14467
rect 23213 14433 23247 14467
rect 23397 14433 23431 14467
rect 24041 14433 24075 14467
rect 2421 14365 2455 14399
rect 4905 14365 4939 14399
rect 6653 14365 6687 14399
rect 8677 14365 8711 14399
rect 9229 14365 9263 14399
rect 12081 14365 12115 14399
rect 15209 14365 15243 14399
rect 15853 14365 15887 14399
rect 16681 14365 16715 14399
rect 18061 14365 18095 14399
rect 20361 14365 20395 14399
rect 22661 14365 22695 14399
rect 24869 14365 24903 14399
rect 26433 14365 26467 14399
rect 3893 14297 3927 14331
rect 5825 14297 5859 14331
rect 7297 14297 7331 14331
rect 10241 14297 10275 14331
rect 1869 14229 1903 14263
rect 2237 14229 2271 14263
rect 4629 14229 4663 14263
rect 4813 14229 4847 14263
rect 7481 14229 7515 14263
rect 8861 14229 8895 14263
rect 10977 14229 11011 14263
rect 13461 14229 13495 14263
rect 15301 14229 15335 14263
rect 17509 14229 17543 14263
rect 19809 14229 19843 14263
rect 20729 14229 20763 14263
rect 23489 14229 23523 14263
rect 3249 14025 3283 14059
rect 6193 14025 6227 14059
rect 10333 14025 10367 14059
rect 11989 14025 12023 14059
rect 15485 14025 15519 14059
rect 16405 14025 16439 14059
rect 20177 14025 20211 14059
rect 24041 14025 24075 14059
rect 26985 14025 27019 14059
rect 2881 13957 2915 13991
rect 4813 13957 4847 13991
rect 7573 13957 7607 13991
rect 8217 13957 8251 13991
rect 15393 13957 15427 13991
rect 18521 13957 18555 13991
rect 5733 13889 5767 13923
rect 7297 13889 7331 13923
rect 9965 13889 9999 13923
rect 18705 13889 18739 13923
rect 19257 13889 19291 13923
rect 1501 13821 1535 13855
rect 3525 13821 3559 13855
rect 3617 13821 3651 13855
rect 3709 13821 3743 13855
rect 3893 13821 3927 13855
rect 3985 13821 4019 13855
rect 4169 13821 4203 13855
rect 4905 13821 4939 13855
rect 5089 13821 5123 13855
rect 5365 13821 5399 13855
rect 6101 13821 6135 13855
rect 6193 13821 6227 13855
rect 6377 13821 6411 13855
rect 7849 13821 7883 13855
rect 8677 13821 8711 13855
rect 8861 13821 8895 13855
rect 9045 13821 9079 13855
rect 9873 13821 9907 13855
rect 10057 13821 10091 13855
rect 10609 13821 10643 13855
rect 14013 13821 14047 13855
rect 14280 13821 14314 13855
rect 15623 13821 15657 13855
rect 16036 13821 16070 13855
rect 16129 13821 16163 13855
rect 16543 13821 16577 13855
rect 16681 13821 16715 13855
rect 16773 13821 16807 13855
rect 16956 13821 16990 13855
rect 17049 13821 17083 13855
rect 17141 13821 17175 13855
rect 19717 13821 19751 13855
rect 19809 13821 19843 13855
rect 19901 13821 19935 13855
rect 20085 13821 20119 13855
rect 20453 13821 20487 13855
rect 20545 13821 20579 13855
rect 20637 13821 20671 13855
rect 20821 13821 20855 13855
rect 20913 13821 20947 13855
rect 21061 13821 21095 13855
rect 21189 13821 21223 13855
rect 21281 13821 21315 13855
rect 21378 13821 21412 13855
rect 21649 13821 21683 13855
rect 21833 13821 21867 13855
rect 21925 13821 21959 13855
rect 22017 13821 22051 13855
rect 22937 13821 22971 13855
rect 24179 13821 24213 13855
rect 24317 13821 24351 13855
rect 24409 13821 24443 13855
rect 24592 13821 24626 13855
rect 24685 13821 24719 13855
rect 24961 13821 24995 13855
rect 25605 13821 25639 13855
rect 25698 13821 25732 13855
rect 25881 13821 25915 13855
rect 25973 13821 26007 13855
rect 26070 13821 26104 13855
rect 26341 13821 26375 13855
rect 26489 13821 26523 13855
rect 26617 13821 26651 13855
rect 26709 13821 26743 13855
rect 26806 13821 26840 13855
rect 1768 13753 1802 13787
rect 5917 13753 5951 13787
rect 8033 13753 8067 13787
rect 10149 13753 10183 13787
rect 10349 13753 10383 13787
rect 10876 13753 10910 13787
rect 15761 13753 15795 13787
rect 15853 13753 15887 13787
rect 17408 13753 17442 13787
rect 22293 13753 22327 13787
rect 4353 13685 4387 13719
rect 5181 13685 5215 13719
rect 5549 13685 5583 13719
rect 7757 13685 7791 13719
rect 10517 13685 10551 13719
rect 19441 13685 19475 13719
rect 21557 13685 21591 13719
rect 22385 13685 22419 13719
rect 25513 13685 25547 13719
rect 26249 13685 26283 13719
rect 1777 13481 1811 13515
rect 5917 13481 5951 13515
rect 8309 13481 8343 13515
rect 10793 13481 10827 13515
rect 16129 13481 16163 13515
rect 17693 13481 17727 13515
rect 18613 13481 18647 13515
rect 21097 13481 21131 13515
rect 24869 13481 24903 13515
rect 1961 13413 1995 13447
rect 2789 13413 2823 13447
rect 3985 13413 4019 13447
rect 5273 13413 5307 13447
rect 5365 13413 5399 13447
rect 5503 13413 5537 13447
rect 12725 13413 12759 13447
rect 21916 13413 21950 13447
rect 1685 13345 1719 13379
rect 2329 13345 2363 13379
rect 2421 13345 2455 13379
rect 2513 13345 2547 13379
rect 2697 13345 2731 13379
rect 3709 13345 3743 13379
rect 5181 13345 5215 13379
rect 5825 13345 5859 13379
rect 6009 13345 6043 13379
rect 6561 13345 6595 13379
rect 6929 13345 6963 13379
rect 7196 13345 7230 13379
rect 8401 13345 8435 13379
rect 8493 13345 8527 13379
rect 9965 13345 9999 13379
rect 10333 13345 10367 13379
rect 10425 13345 10459 13379
rect 11069 13345 11103 13379
rect 11217 13345 11251 13379
rect 11345 13345 11379 13379
rect 11437 13345 11471 13379
rect 11575 13345 11609 13379
rect 14841 13345 14875 13379
rect 14933 13345 14967 13379
rect 15025 13345 15059 13379
rect 15209 13345 15243 13379
rect 17969 13345 18003 13379
rect 18061 13345 18095 13379
rect 18153 13345 18187 13379
rect 18337 13345 18371 13379
rect 18429 13345 18463 13379
rect 19533 13345 19567 13379
rect 19717 13345 19751 13379
rect 19984 13345 20018 13379
rect 21649 13345 21683 13379
rect 23756 13345 23790 13379
rect 24961 13345 24995 13379
rect 26985 13345 27019 13379
rect 1888 13277 1922 13311
rect 3433 13277 3467 13311
rect 3893 13277 3927 13311
rect 5641 13277 5675 13311
rect 6285 13277 6319 13311
rect 10517 13277 10551 13311
rect 10609 13277 10643 13311
rect 13369 13277 13403 13311
rect 14289 13277 14323 13311
rect 15853 13277 15887 13311
rect 16681 13277 16715 13311
rect 16957 13277 16991 13311
rect 23489 13277 23523 13311
rect 25513 13277 25547 13311
rect 3525 13209 3559 13243
rect 6377 13209 6411 13243
rect 8769 13209 8803 13243
rect 2053 13141 2087 13175
rect 3985 13141 4019 13175
rect 4997 13141 5031 13175
rect 6745 13141 6779 13175
rect 8401 13141 8435 13175
rect 9781 13141 9815 13175
rect 11713 13141 11747 13175
rect 13645 13141 13679 13175
rect 14565 13141 14599 13175
rect 15301 13141 15335 13175
rect 17601 13141 17635 13175
rect 18981 13141 19015 13175
rect 23029 13141 23063 13175
rect 26433 13141 26467 13175
rect 2973 12937 3007 12971
rect 4169 12937 4203 12971
rect 4353 12937 4387 12971
rect 7389 12937 7423 12971
rect 11069 12937 11103 12971
rect 15485 12937 15519 12971
rect 16589 12937 16623 12971
rect 22937 12937 22971 12971
rect 25237 12937 25271 12971
rect 26709 12937 26743 12971
rect 2789 12869 2823 12903
rect 4721 12869 4755 12903
rect 7665 12869 7699 12903
rect 4077 12801 4111 12835
rect 4445 12801 4479 12835
rect 17969 12801 18003 12835
rect 18705 12801 18739 12835
rect 21097 12801 21131 12835
rect 25329 12801 25363 12835
rect 1409 12733 1443 12767
rect 2881 12733 2915 12767
rect 3430 12733 3464 12767
rect 3801 12733 3835 12767
rect 3893 12733 3927 12767
rect 3985 12733 4019 12767
rect 4629 12733 4663 12767
rect 4721 12733 4755 12767
rect 4905 12733 4939 12767
rect 7573 12733 7607 12767
rect 7757 12733 7791 12767
rect 7849 12733 7883 12767
rect 8401 12733 8435 12767
rect 9597 12733 9631 12767
rect 9965 12733 9999 12767
rect 10885 12733 10919 12767
rect 14105 12733 14139 12767
rect 14372 12733 14406 12767
rect 15669 12733 15703 12767
rect 18245 12733 18279 12767
rect 23857 12733 23891 12767
rect 23950 12733 23984 12767
rect 24133 12733 24167 12767
rect 24322 12733 24356 12767
rect 24593 12733 24627 12767
rect 24777 12733 24811 12767
rect 24869 12733 24903 12767
rect 24961 12733 24995 12767
rect 1676 12665 1710 12699
rect 5172 12665 5206 12699
rect 17702 12665 17736 12699
rect 20453 12665 20487 12699
rect 21649 12665 21683 12699
rect 24225 12665 24259 12699
rect 25596 12665 25630 12699
rect 3249 12597 3283 12631
rect 3433 12597 3467 12631
rect 6285 12597 6319 12631
rect 8585 12597 8619 12631
rect 9413 12597 9447 12631
rect 9781 12597 9815 12631
rect 15761 12597 15795 12631
rect 18429 12597 18463 12631
rect 20545 12597 20579 12631
rect 24501 12597 24535 12631
rect 3801 12393 3835 12427
rect 5273 12393 5307 12427
rect 14749 12393 14783 12427
rect 16221 12393 16255 12427
rect 16957 12393 16991 12427
rect 20085 12393 20119 12427
rect 22753 12393 22787 12427
rect 25513 12393 25547 12427
rect 26433 12393 26467 12427
rect 7021 12325 7055 12359
rect 8677 12325 8711 12359
rect 9781 12325 9815 12359
rect 18880 12325 18914 12359
rect 2605 12257 2639 12291
rect 2697 12257 2731 12291
rect 2789 12257 2823 12291
rect 2973 12257 3007 12291
rect 4261 12257 4295 12291
rect 4997 12257 5031 12291
rect 5181 12257 5215 12291
rect 5457 12257 5491 12291
rect 7205 12257 7239 12291
rect 7481 12257 7515 12291
rect 7757 12257 7791 12291
rect 7941 12257 7975 12291
rect 8953 12257 8987 12291
rect 9137 12257 9171 12291
rect 9505 12257 9539 12291
rect 9965 12257 9999 12291
rect 10241 12257 10275 12291
rect 10977 12257 11011 12291
rect 11161 12257 11195 12291
rect 11437 12257 11471 12291
rect 11704 12257 11738 12291
rect 13369 12257 13403 12291
rect 13636 12257 13670 12291
rect 14841 12257 14875 12291
rect 15485 12257 15519 12291
rect 15669 12257 15703 12291
rect 15945 12257 15979 12291
rect 16129 12257 16163 12291
rect 16313 12257 16347 12291
rect 17233 12257 17267 12291
rect 17325 12257 17359 12291
rect 17417 12257 17451 12291
rect 17601 12257 17635 12291
rect 18613 12257 18647 12291
rect 20361 12257 20395 12291
rect 20453 12257 20487 12291
rect 20545 12257 20579 12291
rect 20729 12257 20763 12291
rect 22109 12257 22143 12291
rect 22293 12257 22327 12291
rect 22385 12257 22419 12291
rect 22477 12257 22511 12291
rect 22845 12257 22879 12291
rect 23489 12257 23523 12291
rect 23581 12257 23615 12291
rect 24777 12257 24811 12291
rect 24961 12257 24995 12291
rect 25053 12257 25087 12291
rect 25145 12257 25179 12291
rect 25789 12257 25823 12291
rect 25881 12257 25915 12291
rect 25973 12257 26007 12291
rect 26157 12257 26191 12291
rect 3065 12189 3099 12223
rect 3617 12189 3651 12223
rect 4813 12189 4847 12223
rect 6837 12189 6871 12223
rect 8033 12189 8067 12223
rect 9229 12189 9263 12223
rect 9321 12189 9355 12223
rect 10149 12189 10183 12223
rect 21925 12189 21959 12223
rect 26985 12189 27019 12223
rect 7573 12121 7607 12155
rect 7665 12121 7699 12155
rect 10425 12121 10459 12155
rect 19993 12121 20027 12155
rect 23765 12121 23799 12155
rect 2329 12053 2363 12087
rect 3985 12053 4019 12087
rect 7297 12053 7331 12087
rect 9689 12053 9723 12087
rect 11345 12053 11379 12087
rect 12817 12053 12851 12087
rect 15853 12053 15887 12087
rect 21373 12053 21407 12087
rect 25421 12053 25455 12087
rect 3065 11849 3099 11883
rect 8953 11849 8987 11883
rect 12081 11849 12115 11883
rect 13369 11849 13403 11883
rect 15117 11849 15151 11883
rect 17417 11849 17451 11883
rect 18245 11849 18279 11883
rect 19349 11849 19383 11883
rect 20085 11849 20119 11883
rect 22569 11849 22603 11883
rect 23489 11849 23523 11883
rect 26249 11849 26283 11883
rect 15209 11781 15243 11815
rect 22477 11781 22511 11815
rect 11345 11713 11379 11747
rect 14105 11713 14139 11747
rect 14473 11713 14507 11747
rect 15761 11713 15795 11747
rect 23121 11713 23155 11747
rect 24409 11713 24443 11747
rect 24869 11713 24903 11747
rect 1685 11645 1719 11679
rect 8401 11645 8435 11679
rect 8493 11645 8527 11679
rect 8677 11645 8711 11679
rect 8769 11645 8803 11679
rect 11437 11645 11471 11679
rect 11621 11645 11655 11679
rect 11713 11645 11747 11679
rect 11805 11645 11839 11679
rect 12725 11645 12759 11679
rect 12909 11645 12943 11679
rect 13001 11645 13035 11679
rect 13093 11645 13127 11679
rect 16221 11645 16255 11679
rect 16497 11645 16531 11679
rect 16957 11645 16991 11679
rect 17233 11645 17267 11679
rect 17775 11623 17809 11657
rect 18061 11645 18095 11679
rect 18705 11645 18739 11679
rect 18798 11645 18832 11679
rect 18981 11645 19015 11679
rect 19211 11645 19245 11679
rect 19441 11645 19475 11679
rect 19534 11645 19568 11679
rect 19906 11645 19940 11679
rect 21097 11645 21131 11679
rect 23305 11645 23339 11679
rect 25136 11645 25170 11679
rect 26893 11645 26927 11679
rect 1952 11577 1986 11611
rect 6285 11577 6319 11611
rect 8033 11577 8067 11611
rect 9597 11577 9631 11611
rect 12265 11577 12299 11611
rect 12449 11577 12483 11611
rect 16037 11577 16071 11611
rect 19073 11577 19107 11611
rect 19717 11577 19751 11611
rect 19809 11577 19843 11611
rect 21364 11577 21398 11611
rect 13553 11509 13587 11543
rect 14657 11509 14691 11543
rect 14749 11509 14783 11543
rect 15577 11509 15611 11543
rect 15669 11509 15703 11543
rect 16405 11509 16439 11543
rect 17049 11509 17083 11543
rect 17877 11509 17911 11543
rect 23857 11509 23891 11543
rect 26341 11509 26375 11543
rect 3525 11305 3559 11339
rect 7205 11305 7239 11339
rect 10609 11305 10643 11339
rect 12265 11305 12299 11339
rect 13737 11305 13771 11339
rect 18521 11305 18555 11339
rect 20085 11305 20119 11339
rect 21281 11305 21315 11339
rect 24133 11305 24167 11339
rect 26249 11305 26283 11339
rect 6092 11237 6126 11271
rect 8401 11237 8435 11271
rect 9496 11237 9530 11271
rect 12602 11237 12636 11271
rect 13921 11237 13955 11271
rect 3341 11169 3375 11203
rect 4629 11169 4663 11203
rect 8217 11169 8251 11203
rect 8493 11169 8527 11203
rect 8677 11169 8711 11203
rect 8769 11169 8803 11203
rect 8861 11169 8895 11203
rect 12357 11169 12391 11203
rect 14013 11169 14047 11203
rect 14105 11169 14139 11203
rect 15117 11169 15151 11203
rect 15301 11169 15335 11203
rect 18061 11169 18095 11203
rect 18153 11169 18187 11203
rect 18337 11169 18371 11203
rect 18613 11169 18647 11203
rect 18797 11169 18831 11203
rect 18889 11169 18923 11203
rect 18981 11169 19015 11203
rect 21557 11169 21591 11203
rect 21649 11169 21683 11203
rect 21741 11169 21775 11203
rect 21925 11169 21959 11203
rect 22109 11169 22143 11203
rect 23020 11169 23054 11203
rect 24869 11169 24903 11203
rect 25136 11169 25170 11203
rect 26433 11169 26467 11203
rect 5825 11101 5859 11135
rect 7297 11101 7331 11135
rect 9229 11101 9263 11135
rect 11713 11101 11747 11135
rect 14749 11101 14783 11135
rect 17969 11101 18003 11135
rect 19257 11101 19291 11135
rect 19901 11101 19935 11135
rect 20729 11101 20763 11135
rect 22753 11101 22787 11135
rect 26985 11101 27019 11135
rect 4813 11033 4847 11067
rect 8033 11033 8067 11067
rect 15485 11033 15519 11067
rect 7941 10965 7975 10999
rect 9137 10965 9171 10999
rect 14289 10965 14323 10999
rect 17325 10965 17359 10999
rect 19349 10965 19383 10999
rect 22293 10965 22327 10999
rect 7205 10761 7239 10795
rect 8217 10761 8251 10795
rect 10977 10761 11011 10795
rect 12449 10761 12483 10795
rect 14841 10761 14875 10795
rect 17233 10761 17267 10795
rect 20085 10761 20119 10795
rect 22017 10761 22051 10795
rect 23857 10761 23891 10795
rect 26617 10761 26651 10795
rect 14289 10625 14323 10659
rect 18705 10625 18739 10659
rect 23581 10625 23615 10659
rect 24409 10625 24443 10659
rect 25237 10625 25271 10659
rect 4353 10557 4387 10591
rect 5825 10557 5859 10591
rect 7573 10557 7607 10591
rect 7721 10557 7755 10591
rect 7941 10557 7975 10591
rect 8038 10557 8072 10591
rect 8861 10557 8895 10591
rect 9045 10557 9079 10591
rect 9137 10557 9171 10591
rect 9229 10557 9263 10591
rect 9597 10557 9631 10591
rect 12725 10557 12759 10591
rect 12817 10557 12851 10591
rect 12909 10557 12943 10591
rect 13093 10557 13127 10591
rect 15025 10557 15059 10591
rect 15209 10557 15243 10591
rect 15301 10557 15335 10591
rect 15393 10557 15427 10591
rect 15853 10557 15887 10591
rect 17877 10557 17911 10591
rect 18972 10557 19006 10591
rect 20177 10557 20211 10591
rect 22201 10557 22235 10591
rect 22385 10557 22419 10591
rect 22477 10557 22511 10591
rect 22937 10557 22971 10591
rect 23121 10557 23155 10591
rect 23213 10557 23247 10591
rect 23305 10557 23339 10591
rect 24777 10557 24811 10591
rect 25053 10557 25087 10591
rect 4620 10489 4654 10523
rect 6092 10489 6126 10523
rect 7849 10489 7883 10523
rect 9505 10489 9539 10523
rect 9842 10489 9876 10523
rect 16098 10489 16132 10523
rect 24593 10489 24627 10523
rect 25482 10489 25516 10523
rect 5733 10421 5767 10455
rect 14381 10421 14415 10455
rect 14473 10421 14507 10455
rect 15669 10421 15703 10455
rect 17325 10421 17359 10455
rect 20361 10421 20395 10455
rect 24961 10421 24995 10455
rect 2145 10217 2179 10251
rect 6009 10217 6043 10251
rect 7941 10217 7975 10251
rect 8953 10217 8987 10251
rect 12817 10217 12851 10251
rect 13369 10217 13403 10251
rect 14197 10217 14231 10251
rect 15669 10217 15703 10251
rect 15853 10217 15887 10251
rect 20269 10217 20303 10251
rect 21925 10217 21959 10251
rect 22109 10217 22143 10251
rect 22937 10217 22971 10251
rect 25421 10217 25455 10251
rect 2688 10149 2722 10183
rect 8677 10149 8711 10183
rect 12541 10149 12575 10183
rect 18797 10149 18831 10183
rect 19134 10149 19168 10183
rect 21557 10149 21591 10183
rect 22477 10149 22511 10183
rect 2421 10081 2455 10115
rect 4997 10081 5031 10115
rect 5457 10081 5491 10115
rect 6193 10081 6227 10115
rect 6469 10081 6503 10115
rect 6653 10081 6687 10115
rect 7021 10081 7055 10115
rect 7205 10081 7239 10115
rect 7297 10081 7331 10115
rect 8309 10081 8343 10115
rect 8457 10081 8491 10115
rect 8585 10081 8619 10115
rect 8815 10081 8849 10115
rect 9045 10081 9079 10115
rect 9301 10081 9335 10115
rect 12173 10081 12207 10115
rect 12266 10081 12300 10115
rect 12449 10081 12483 10115
rect 12638 10081 12672 10115
rect 13737 10081 13771 10115
rect 14565 10081 14599 10115
rect 15025 10081 15059 10115
rect 15761 10081 15795 10115
rect 15945 10081 15979 10115
rect 16681 10081 16715 10115
rect 17049 10081 17083 10115
rect 17141 10081 17175 10115
rect 17325 10081 17359 10115
rect 18889 10081 18923 10115
rect 20913 10081 20947 10115
rect 21465 10081 21499 10115
rect 21741 10081 21775 10115
rect 22017 10081 22051 10115
rect 22293 10081 22327 10115
rect 23121 10081 23155 10115
rect 23305 10081 23339 10115
rect 23397 10081 23431 10115
rect 24065 10081 24099 10115
rect 24225 10081 24259 10115
rect 24317 10081 24351 10115
rect 24409 10081 24443 10115
rect 24777 10081 24811 10115
rect 24961 10081 24995 10115
rect 25053 10081 25087 10115
rect 25145 10081 25179 10115
rect 25697 10081 25731 10115
rect 25881 10081 25915 10115
rect 25973 10081 26007 10115
rect 26985 10081 27019 10115
rect 4813 10013 4847 10047
rect 5273 10013 5307 10047
rect 5641 10013 5675 10047
rect 6837 10013 6871 10047
rect 13829 10013 13863 10047
rect 14013 10013 14047 10047
rect 14657 10013 14691 10047
rect 14749 10013 14783 10047
rect 17969 10013 18003 10047
rect 18245 10013 18279 10047
rect 25513 10013 25547 10047
rect 1777 9945 1811 9979
rect 6285 9945 6319 9979
rect 6377 9945 6411 9979
rect 17325 9945 17359 9979
rect 20361 9945 20395 9979
rect 24685 9945 24719 9979
rect 26433 9945 26467 9979
rect 2145 9877 2179 9911
rect 2329 9877 2363 9911
rect 3801 9877 3835 9911
rect 5181 9877 5215 9911
rect 10425 9877 10459 9911
rect 16129 9877 16163 9911
rect 17417 9877 17451 9911
rect 5641 9673 5675 9707
rect 18981 9673 19015 9707
rect 2789 9605 2823 9639
rect 2881 9605 2915 9639
rect 3985 9605 4019 9639
rect 6101 9605 6135 9639
rect 14473 9605 14507 9639
rect 16681 9605 16715 9639
rect 20545 9605 20579 9639
rect 21373 9605 21407 9639
rect 24685 9605 24719 9639
rect 24869 9605 24903 9639
rect 3801 9537 3835 9571
rect 4905 9537 4939 9571
rect 5273 9537 5307 9571
rect 5733 9537 5767 9571
rect 11621 9537 11655 9571
rect 16957 9537 16991 9571
rect 17049 9537 17083 9571
rect 17325 9537 17359 9571
rect 17509 9537 17543 9571
rect 22753 9537 22787 9571
rect 23213 9537 23247 9571
rect 23305 9537 23339 9571
rect 1409 9469 1443 9503
rect 3065 9469 3099 9503
rect 4169 9469 4203 9503
rect 4445 9469 4479 9503
rect 4721 9469 4755 9503
rect 5457 9469 5491 9503
rect 5917 9469 5951 9503
rect 6009 9469 6043 9503
rect 6193 9469 6227 9503
rect 6377 9469 6411 9503
rect 7665 9469 7699 9503
rect 8953 9469 8987 9503
rect 9137 9469 9171 9503
rect 9229 9469 9263 9503
rect 9321 9469 9355 9503
rect 9689 9469 9723 9503
rect 16129 9469 16163 9503
rect 16221 9469 16255 9503
rect 16313 9469 16347 9503
rect 16497 9469 16531 9503
rect 16865 9469 16899 9503
rect 17141 9469 17175 9503
rect 17601 9469 17635 9503
rect 19257 9469 19291 9503
rect 19349 9469 19383 9503
rect 19441 9469 19475 9503
rect 19625 9469 19659 9503
rect 19901 9469 19935 9503
rect 20177 9469 20211 9503
rect 20361 9469 20395 9503
rect 23029 9469 23063 9503
rect 23121 9469 23155 9503
rect 24225 9469 24259 9503
rect 24501 9469 24535 9503
rect 25053 9469 25087 9503
rect 25329 9469 25363 9503
rect 1676 9401 1710 9435
rect 4353 9401 4387 9435
rect 9934 9401 9968 9435
rect 11888 9401 11922 9435
rect 15761 9401 15795 9435
rect 19717 9401 19751 9435
rect 22486 9401 22520 9435
rect 3249 9333 3283 9367
rect 4537 9333 4571 9367
rect 8217 9333 8251 9367
rect 9597 9333 9631 9367
rect 11069 9333 11103 9367
rect 13001 9333 13035 9367
rect 15853 9333 15887 9367
rect 17325 9333 17359 9367
rect 20085 9333 20119 9367
rect 22845 9333 22879 9367
rect 24317 9333 24351 9367
rect 25237 9333 25271 9367
rect 1691 9129 1725 9163
rect 4445 9129 4479 9163
rect 4997 9129 5031 9163
rect 8125 9129 8159 9163
rect 9321 9129 9355 9163
rect 11897 9129 11931 9163
rect 12633 9129 12667 9163
rect 14381 9129 14415 9163
rect 17877 9129 17911 9163
rect 19165 9129 19199 9163
rect 22661 9129 22695 9163
rect 23949 9129 23983 9163
rect 1777 9061 1811 9095
rect 5181 9061 5215 9095
rect 8401 9061 8435 9095
rect 9045 9061 9079 9095
rect 15494 9061 15528 9095
rect 23029 9061 23063 9095
rect 23673 9061 23707 9095
rect 25154 9061 25188 9095
rect 25697 9061 25731 9095
rect 1593 8993 1627 9027
rect 1869 8993 1903 9027
rect 1961 8993 1995 9027
rect 2973 8993 3007 9027
rect 3893 8993 3927 9027
rect 4077 8993 4111 9027
rect 4629 8993 4663 9027
rect 4905 8993 4939 9027
rect 6745 8993 6779 9027
rect 7012 8993 7046 9027
rect 8585 8993 8619 9027
rect 8677 8993 8711 9027
rect 8770 8993 8804 9027
rect 8953 8993 8987 9027
rect 9142 8993 9176 9027
rect 13185 8993 13219 9027
rect 13548 8993 13582 9027
rect 13645 8993 13679 9027
rect 13737 8993 13771 9027
rect 13920 8993 13954 9027
rect 14013 8993 14047 9027
rect 16764 8993 16798 9027
rect 18521 8993 18555 9027
rect 18705 8993 18739 9027
rect 18797 8993 18831 9027
rect 18981 8993 19015 9027
rect 19809 8993 19843 9027
rect 21281 8993 21315 9027
rect 21465 8993 21499 9027
rect 22753 8993 22787 9027
rect 22845 8993 22879 9027
rect 23305 8993 23339 9027
rect 23397 8993 23431 9027
rect 23489 8993 23523 9027
rect 23765 8993 23799 9027
rect 25513 8993 25547 9027
rect 25789 8993 25823 9027
rect 26157 8993 26191 9027
rect 2237 8925 2271 8959
rect 3157 8925 3191 8959
rect 3801 8925 3835 8959
rect 4353 8925 4387 8959
rect 4813 8925 4847 8959
rect 12449 8925 12483 8959
rect 15761 8925 15795 8959
rect 16497 8925 16531 8959
rect 22385 8925 22419 8959
rect 22477 8925 22511 8959
rect 25421 8925 25455 8959
rect 2053 8857 2087 8891
rect 2145 8857 2179 8891
rect 5181 8857 5215 8891
rect 13369 8857 13403 8891
rect 24041 8857 24075 8891
rect 25973 8857 26007 8891
rect 2329 8789 2363 8823
rect 4261 8789 4295 8823
rect 8217 8789 8251 8823
rect 17969 8789 18003 8823
rect 19625 8789 19659 8823
rect 21373 8789 21407 8823
rect 21741 8789 21775 8823
rect 23121 8789 23155 8823
rect 25513 8789 25547 8823
rect 2973 8585 3007 8619
rect 7021 8585 7055 8619
rect 14933 8585 14967 8619
rect 16405 8585 16439 8619
rect 17141 8585 17175 8619
rect 20637 8585 20671 8619
rect 22201 8585 22235 8619
rect 22753 8585 22787 8619
rect 22937 8585 22971 8619
rect 24133 8585 24167 8619
rect 11805 8517 11839 8551
rect 17785 8517 17819 8551
rect 22385 8517 22419 8551
rect 24041 8517 24075 8551
rect 3801 8449 3835 8483
rect 11897 8449 11931 8483
rect 16313 8449 16347 8483
rect 19257 8449 19291 8483
rect 20913 8449 20947 8483
rect 21189 8449 21223 8483
rect 24225 8449 24259 8483
rect 24961 8449 24995 8483
rect 25145 8449 25179 8483
rect 1593 8381 1627 8415
rect 3617 8381 3651 8415
rect 3709 8381 3743 8415
rect 3893 8381 3927 8415
rect 4629 8381 4663 8415
rect 5549 8381 5583 8415
rect 5733 8381 5767 8415
rect 7573 8381 7607 8415
rect 7941 8381 7975 8415
rect 9321 8381 9355 8415
rect 9414 8381 9448 8415
rect 9597 8381 9631 8415
rect 9786 8381 9820 8415
rect 11161 8381 11195 8415
rect 11254 8381 11288 8415
rect 11626 8381 11660 8415
rect 12173 8381 12207 8415
rect 12265 8381 12299 8415
rect 12357 8381 12391 8415
rect 12541 8381 12575 8415
rect 12633 8381 12667 8415
rect 12817 8381 12851 8415
rect 12909 8381 12943 8415
rect 13001 8381 13035 8415
rect 16046 8381 16080 8415
rect 16957 8381 16991 8415
rect 17141 8381 17175 8415
rect 17417 8381 17451 8415
rect 17601 8381 17635 8415
rect 19524 8381 19558 8415
rect 21005 8381 21039 8415
rect 21097 8381 21131 8415
rect 21557 8381 21591 8415
rect 21741 8381 21775 8415
rect 21833 8381 21867 8415
rect 21925 8381 21959 8415
rect 23949 8381 23983 8415
rect 24317 8381 24351 8415
rect 1860 8313 1894 8347
rect 4261 8313 4295 8347
rect 5917 8313 5951 8347
rect 8125 8313 8159 8347
rect 8401 8313 8435 8347
rect 8585 8313 8619 8347
rect 9689 8313 9723 8347
rect 11437 8313 11471 8347
rect 11529 8313 11563 8347
rect 17325 8313 17359 8347
rect 22753 8313 22787 8347
rect 25412 8313 25446 8347
rect 3433 8245 3467 8279
rect 4077 8245 4111 8279
rect 4353 8245 4387 8279
rect 4445 8245 4479 8279
rect 7757 8245 7791 8279
rect 8769 8245 8803 8279
rect 9965 8245 9999 8279
rect 13277 8245 13311 8279
rect 20729 8245 20763 8279
rect 26525 8245 26559 8279
rect 2605 8041 2639 8075
rect 4077 8041 4111 8075
rect 6929 8041 6963 8075
rect 8493 8041 8527 8075
rect 9321 8041 9355 8075
rect 19901 8041 19935 8075
rect 21649 8041 21683 8075
rect 21741 8041 21775 8075
rect 24685 8041 24719 8075
rect 26433 8041 26467 8075
rect 2942 7973 2976 8007
rect 9781 7973 9815 8007
rect 13084 7973 13118 8007
rect 2421 7905 2455 7939
rect 2697 7905 2731 7939
rect 6193 7905 6227 7939
rect 6377 7905 6411 7939
rect 6653 7905 6687 7939
rect 7113 7905 7147 7939
rect 7297 7905 7331 7939
rect 7389 7905 7423 7939
rect 7573 7905 7607 7939
rect 9413 7905 9447 7939
rect 9506 7905 9540 7939
rect 9689 7905 9723 7939
rect 9878 7905 9912 7939
rect 10149 7905 10183 7939
rect 10333 7905 10367 7939
rect 10425 7905 10459 7939
rect 10517 7905 10551 7939
rect 11345 7905 11379 7939
rect 12081 7905 12115 7939
rect 12265 7905 12299 7939
rect 12360 7905 12394 7939
rect 12495 7905 12529 7939
rect 20729 7905 20763 7939
rect 21373 7905 21407 7939
rect 21557 7905 21591 7939
rect 22569 7905 22603 7939
rect 23029 7905 23063 7939
rect 23213 7905 23247 7939
rect 23305 7905 23339 7939
rect 23489 7905 23523 7939
rect 24041 7905 24075 7939
rect 24133 7905 24167 7939
rect 24409 7905 24443 7939
rect 25798 7905 25832 7939
rect 26065 7905 26099 7939
rect 26985 7905 27019 7939
rect 7941 7837 7975 7871
rect 8769 7837 8803 7871
rect 11989 7837 12023 7871
rect 12817 7837 12851 7871
rect 21005 7837 21039 7871
rect 22385 7837 22419 7871
rect 22477 7837 22511 7871
rect 22661 7837 22695 7871
rect 23857 7837 23891 7871
rect 24225 7837 24259 7871
rect 6469 7769 6503 7803
rect 6561 7769 6595 7803
rect 7205 7769 7239 7803
rect 10057 7769 10091 7803
rect 19533 7769 19567 7803
rect 20085 7769 20119 7803
rect 23213 7769 23247 7803
rect 23949 7769 23983 7803
rect 6837 7701 6871 7735
rect 10793 7701 10827 7735
rect 12725 7701 12759 7735
rect 14197 7701 14231 7735
rect 19901 7701 19935 7735
rect 21925 7701 21959 7735
rect 22201 7701 22235 7735
rect 22937 7701 22971 7735
rect 24593 7701 24627 7735
rect 3249 7497 3283 7531
rect 3433 7497 3467 7531
rect 5917 7497 5951 7531
rect 7941 7497 7975 7531
rect 15393 7497 15427 7531
rect 15945 7497 15979 7531
rect 18521 7497 18555 7531
rect 25145 7497 25179 7531
rect 25329 7497 25363 7531
rect 4077 7429 4111 7463
rect 19073 7429 19107 7463
rect 3801 7361 3835 7395
rect 3893 7361 3927 7395
rect 6009 7361 6043 7395
rect 8677 7361 8711 7395
rect 17141 7361 17175 7395
rect 4169 7293 4203 7327
rect 4261 7293 4295 7327
rect 4445 7293 4479 7327
rect 4537 7293 4571 7327
rect 5549 7293 5583 7327
rect 5733 7293 5767 7327
rect 6193 7293 6227 7327
rect 6561 7293 6595 7327
rect 6828 7293 6862 7327
rect 8585 7293 8619 7327
rect 8769 7293 8803 7327
rect 8861 7293 8895 7327
rect 9045 7293 9079 7327
rect 9597 7293 9631 7327
rect 11069 7293 11103 7327
rect 13553 7293 13587 7327
rect 13820 7293 13854 7327
rect 15577 7293 15611 7327
rect 15853 7293 15887 7327
rect 16129 7293 16163 7327
rect 16405 7293 16439 7327
rect 18889 7293 18923 7327
rect 19441 7293 19475 7327
rect 21465 7293 21499 7327
rect 21741 7293 21775 7327
rect 25053 7293 25087 7327
rect 25329 7293 25363 7327
rect 25513 7293 25547 7327
rect 25605 7293 25639 7327
rect 25789 7293 25823 7327
rect 3433 7225 3467 7259
rect 3893 7225 3927 7259
rect 6377 7225 6411 7259
rect 9864 7225 9898 7259
rect 11336 7225 11370 7259
rect 17408 7225 17442 7259
rect 19257 7225 19291 7259
rect 23397 7225 23431 7259
rect 4353 7157 4387 7191
rect 4721 7157 4755 7191
rect 8401 7157 8435 7191
rect 10977 7157 11011 7191
rect 12449 7157 12483 7191
rect 14933 7157 14967 7191
rect 15761 7157 15795 7191
rect 16313 7157 16347 7191
rect 18705 7157 18739 7191
rect 19349 7157 19383 7191
rect 19625 7157 19659 7191
rect 21649 7157 21683 7191
rect 25697 7157 25731 7191
rect 4093 6953 4127 6987
rect 4353 6953 4387 6987
rect 5273 6953 5307 6987
rect 5365 6953 5399 6987
rect 5457 6953 5491 6987
rect 8861 6953 8895 6987
rect 13921 6953 13955 6987
rect 18337 6953 18371 6987
rect 23213 6953 23247 6987
rect 23949 6953 23983 6987
rect 24317 6953 24351 6987
rect 25789 6953 25823 6987
rect 3893 6885 3927 6919
rect 18153 6885 18187 6919
rect 22100 6885 22134 6919
rect 24133 6885 24167 6919
rect 1501 6817 1535 6851
rect 1768 6817 1802 6851
rect 4997 6817 5031 6851
rect 7748 6817 7782 6851
rect 9137 6817 9171 6851
rect 11437 6817 11471 6851
rect 12081 6817 12115 6851
rect 12173 6817 12207 6851
rect 12357 6817 12391 6851
rect 13461 6817 13495 6851
rect 13645 6817 13679 6851
rect 13829 6817 13863 6851
rect 14381 6817 14415 6851
rect 14749 6817 14783 6851
rect 14841 6817 14875 6851
rect 15577 6817 15611 6851
rect 18705 6817 18739 6851
rect 18889 6817 18923 6851
rect 20361 6817 20395 6851
rect 20453 6817 20487 6851
rect 20637 6817 20671 6851
rect 20821 6817 20855 6851
rect 24225 6817 24259 6851
rect 24593 6817 24627 6851
rect 25329 6817 25363 6851
rect 25513 6817 25547 6851
rect 26065 6817 26099 6851
rect 26433 6817 26467 6851
rect 3617 6749 3651 6783
rect 7481 6749 7515 6783
rect 8953 6749 8987 6783
rect 14264 6749 14298 6783
rect 14473 6749 14507 6783
rect 15117 6749 15151 6783
rect 18429 6749 18463 6783
rect 18613 6749 18647 6783
rect 18797 6749 18831 6783
rect 19441 6749 19475 6783
rect 21833 6749 21867 6783
rect 25145 6749 25179 6783
rect 25697 6749 25731 6783
rect 25789 6749 25823 6783
rect 26985 6749 27019 6783
rect 2973 6681 3007 6715
rect 5641 6681 5675 6715
rect 13553 6681 13587 6715
rect 14933 6681 14967 6715
rect 17785 6681 17819 6715
rect 20177 6681 20211 6715
rect 24501 6681 24535 6715
rect 2881 6613 2915 6647
rect 4077 6613 4111 6647
rect 4261 6613 4295 6647
rect 5089 6613 5123 6647
rect 9321 6613 9355 6647
rect 12541 6613 12575 6647
rect 14105 6613 14139 6647
rect 15301 6613 15335 6647
rect 15853 6613 15887 6647
rect 18153 6613 18187 6647
rect 20085 6613 20119 6647
rect 20729 6613 20763 6647
rect 25973 6613 26007 6647
rect 2053 6409 2087 6443
rect 2513 6409 2547 6443
rect 4813 6409 4847 6443
rect 6285 6409 6319 6443
rect 11805 6409 11839 6443
rect 14381 6409 14415 6443
rect 18521 6409 18555 6443
rect 22017 6409 22051 6443
rect 22201 6409 22235 6443
rect 24777 6409 24811 6443
rect 24961 6409 24995 6443
rect 26525 6409 26559 6443
rect 9781 6341 9815 6375
rect 11345 6341 11379 6375
rect 13645 6341 13679 6375
rect 15853 6341 15887 6375
rect 23029 6341 23063 6375
rect 2329 6273 2363 6307
rect 10977 6273 11011 6307
rect 12449 6273 12483 6307
rect 15761 6273 15795 6307
rect 17141 6273 17175 6307
rect 21833 6273 21867 6307
rect 22845 6273 22879 6307
rect 24409 6273 24443 6307
rect 25145 6273 25179 6307
rect 2053 6205 2087 6239
rect 2237 6205 2271 6239
rect 2605 6205 2639 6239
rect 2881 6205 2915 6239
rect 3065 6205 3099 6239
rect 3433 6205 3467 6239
rect 4905 6205 4939 6239
rect 8125 6205 8159 6239
rect 8401 6205 8435 6239
rect 10241 6205 10275 6239
rect 10333 6205 10367 6239
rect 10425 6205 10459 6239
rect 10609 6205 10643 6239
rect 10701 6205 10735 6239
rect 11161 6205 11195 6239
rect 11253 6205 11287 6239
rect 11436 6205 11470 6239
rect 11633 6215 11667 6249
rect 12173 6205 12207 6239
rect 13829 6205 13863 6239
rect 16129 6205 16163 6239
rect 16865 6205 16899 6239
rect 17049 6205 17083 6239
rect 18705 6205 18739 6239
rect 20453 6205 20487 6239
rect 20729 6205 20763 6239
rect 21005 6205 21039 6239
rect 21649 6205 21683 6239
rect 21741 6205 21775 6239
rect 23121 6205 23155 6239
rect 23857 6205 23891 6239
rect 25412 6205 25446 6239
rect 2329 6137 2363 6171
rect 2697 6137 2731 6171
rect 3700 6137 3734 6171
rect 5172 6137 5206 6171
rect 6377 6137 6411 6171
rect 8668 6137 8702 6171
rect 10885 6137 10919 6171
rect 15494 6137 15528 6171
rect 15853 6137 15887 6171
rect 16957 6137 16991 6171
rect 17386 6137 17420 6171
rect 20545 6137 20579 6171
rect 22185 6137 22219 6171
rect 22385 6137 22419 6171
rect 24593 6137 24627 6171
rect 24793 6137 24827 6171
rect 10057 6069 10091 6103
rect 12265 6069 12299 6103
rect 16037 6069 16071 6103
rect 20913 6069 20947 6103
rect 22845 6069 22879 6103
rect 6469 5865 6503 5899
rect 8677 5865 8711 5899
rect 14933 5865 14967 5899
rect 17325 5865 17359 5899
rect 17693 5865 17727 5899
rect 20821 5865 20855 5899
rect 24041 5865 24075 5899
rect 24593 5865 24627 5899
rect 4997 5797 5031 5831
rect 13185 5797 13219 5831
rect 18153 5797 18187 5831
rect 19708 5797 19742 5831
rect 21433 5797 21467 5831
rect 21649 5797 21683 5831
rect 5181 5729 5215 5763
rect 5273 5729 5307 5763
rect 5365 5729 5399 5763
rect 5549 5729 5583 5763
rect 5917 5729 5951 5763
rect 8493 5729 8527 5763
rect 8953 5729 8987 5763
rect 9137 5729 9171 5763
rect 10977 5729 11011 5763
rect 11244 5729 11278 5763
rect 13645 5729 13679 5763
rect 14013 5729 14047 5763
rect 14197 5729 14231 5763
rect 14749 5729 14783 5763
rect 14841 5729 14875 5763
rect 15025 5729 15059 5763
rect 17601 5729 17635 5763
rect 17877 5729 17911 5763
rect 18061 5729 18095 5763
rect 18705 5729 18739 5763
rect 19441 5729 19475 5763
rect 21097 5729 21131 5763
rect 22385 5729 22419 5763
rect 22569 5729 22603 5763
rect 22661 5729 22695 5763
rect 22917 5729 22951 5763
rect 24501 5729 24535 5763
rect 25706 5729 25740 5763
rect 25973 5729 26007 5763
rect 4997 5661 5031 5695
rect 8217 5661 8251 5695
rect 13001 5661 13035 5695
rect 17325 5661 17359 5695
rect 22477 5661 22511 5695
rect 12357 5593 12391 5627
rect 12449 5593 12483 5627
rect 17509 5593 17543 5627
rect 21281 5593 21315 5627
rect 5365 5525 5399 5559
rect 8309 5525 8343 5559
rect 8769 5525 8803 5559
rect 14565 5525 14599 5559
rect 20913 5525 20947 5559
rect 21465 5525 21499 5559
rect 24409 5525 24443 5559
rect 10149 5321 10183 5355
rect 11713 5321 11747 5355
rect 13553 5321 13587 5355
rect 14381 5321 14415 5355
rect 19901 5321 19935 5355
rect 22753 5321 22787 5355
rect 23489 5321 23523 5355
rect 24409 5321 24443 5355
rect 25789 5321 25823 5355
rect 12541 5253 12575 5287
rect 16681 5253 16715 5287
rect 9045 5185 9079 5219
rect 12357 5185 12391 5219
rect 13093 5185 13127 5219
rect 14197 5185 14231 5219
rect 14933 5185 14967 5219
rect 17233 5185 17267 5219
rect 19349 5185 19383 5219
rect 21281 5185 21315 5219
rect 4261 5117 4295 5151
rect 5917 5117 5951 5151
rect 6469 5117 6503 5151
rect 6837 5117 6871 5151
rect 6929 5117 6963 5151
rect 7021 5117 7055 5151
rect 7205 5117 7239 5151
rect 7941 5117 7975 5151
rect 8125 5117 8159 5151
rect 8585 5117 8619 5151
rect 8677 5117 8711 5151
rect 8861 5117 8895 5151
rect 8953 5117 8987 5151
rect 9229 5117 9263 5151
rect 9321 5117 9355 5151
rect 9505 5117 9539 5151
rect 9597 5117 9631 5151
rect 11437 5117 11471 5151
rect 12081 5117 12115 5151
rect 12909 5117 12943 5151
rect 15485 5117 15519 5151
rect 15669 5117 15703 5151
rect 15853 5117 15887 5151
rect 16129 5117 16163 5151
rect 16313 5117 16347 5151
rect 16401 5117 16435 5151
rect 16497 5117 16531 5151
rect 16865 5117 16899 5151
rect 16957 5117 16991 5151
rect 17417 5117 17451 5151
rect 17601 5117 17635 5151
rect 18061 5117 18095 5151
rect 18797 5117 18831 5151
rect 18889 5117 18923 5151
rect 19257 5117 19291 5151
rect 21014 5117 21048 5151
rect 22385 5117 22419 5151
rect 23029 5117 23063 5151
rect 23213 5117 23247 5151
rect 23857 5117 23891 5151
rect 24041 5117 24075 5151
rect 24317 5117 24351 5151
rect 24501 5117 24535 5151
rect 24593 5117 24627 5151
rect 25145 5117 25179 5151
rect 4528 5049 4562 5083
rect 6561 5049 6595 5083
rect 8401 5049 8435 5083
rect 14749 5049 14783 5083
rect 14841 5049 14875 5083
rect 15761 5049 15795 5083
rect 19073 5049 19107 5083
rect 19165 5049 19199 5083
rect 22569 5049 22603 5083
rect 23305 5049 23339 5083
rect 23521 5049 23555 5083
rect 23949 5049 23983 5083
rect 24133 5049 24167 5083
rect 5641 4981 5675 5015
rect 7941 4981 7975 5015
rect 12173 4981 12207 5015
rect 13001 4981 13035 5015
rect 13921 4981 13955 5015
rect 14013 4981 14047 5015
rect 16037 4981 16071 5015
rect 17141 4981 17175 5015
rect 18245 4981 18279 5015
rect 22845 4981 22879 5015
rect 23673 4981 23707 5015
rect 11621 4777 11655 4811
rect 15301 4777 15335 4811
rect 23949 4777 23983 4811
rect 5825 4709 5859 4743
rect 6837 4709 6871 4743
rect 19134 4709 19168 4743
rect 3709 4641 3743 4675
rect 3801 4641 3835 4675
rect 3893 4641 3927 4675
rect 4077 4641 4111 4675
rect 5181 4641 5215 4675
rect 5273 4641 5307 4675
rect 5365 4641 5399 4675
rect 5549 4641 5583 4675
rect 6745 4641 6779 4675
rect 6929 4641 6963 4675
rect 7113 4641 7147 4675
rect 7481 4641 7515 4675
rect 7573 4641 7607 4675
rect 7757 4641 7791 4675
rect 7849 4641 7883 4675
rect 8125 4641 8159 4675
rect 8217 4641 8251 4675
rect 8401 4641 8435 4675
rect 8493 4641 8527 4675
rect 8585 4641 8619 4675
rect 8677 4641 8711 4675
rect 8861 4641 8895 4675
rect 8953 4641 8987 4675
rect 9229 4641 9263 4675
rect 9321 4641 9355 4675
rect 9459 4641 9493 4675
rect 9597 4641 9631 4675
rect 10241 4641 10275 4675
rect 10333 4641 10367 4675
rect 10517 4641 10551 4675
rect 10609 4641 10643 4675
rect 10977 4641 11011 4675
rect 11161 4641 11195 4675
rect 11253 4641 11287 4675
rect 11345 4641 11379 4675
rect 12173 4641 12207 4675
rect 12357 4641 12391 4675
rect 12449 4641 12483 4675
rect 12541 4641 12575 4675
rect 15117 4641 15151 4675
rect 17141 4641 17175 4675
rect 17417 4641 17451 4675
rect 17673 4641 17707 4675
rect 18889 4641 18923 4675
rect 22569 4641 22603 4675
rect 22836 4641 22870 4675
rect 4813 4573 4847 4607
rect 6377 4573 6411 4607
rect 7297 4505 7331 4539
rect 17325 4505 17359 4539
rect 3433 4437 3467 4471
rect 4169 4437 4203 4471
rect 4905 4437 4939 4471
rect 6561 4437 6595 4471
rect 7941 4437 7975 4471
rect 9137 4437 9171 4471
rect 9781 4437 9815 4471
rect 10793 4437 10827 4471
rect 12725 4437 12759 4471
rect 18797 4437 18831 4471
rect 20269 4437 20303 4471
rect 5457 4233 5491 4267
rect 12633 4233 12667 4267
rect 13553 4233 13587 4267
rect 22845 4233 22879 4267
rect 15853 4165 15887 4199
rect 13277 4097 13311 4131
rect 14197 4097 14231 4131
rect 19073 4097 19107 4131
rect 19441 4097 19475 4131
rect 3801 4029 3835 4063
rect 3985 4029 4019 4063
rect 4077 4029 4111 4063
rect 7113 4029 7147 4063
rect 7205 4029 7239 4063
rect 7297 4029 7331 4063
rect 7481 4029 7515 4063
rect 8125 4029 8159 4063
rect 8861 4029 8895 4063
rect 8953 4029 8987 4063
rect 9045 4029 9079 4063
rect 9229 4029 9263 4063
rect 9873 4029 9907 4063
rect 10333 4029 10367 4063
rect 10425 4029 10459 4063
rect 10517 4029 10551 4063
rect 10701 4029 10735 4063
rect 10977 4029 11011 4063
rect 11161 4029 11195 4063
rect 11253 4029 11287 4063
rect 11345 4029 11379 4063
rect 11897 4029 11931 4063
rect 12449 4029 12483 4063
rect 13093 4029 13127 4063
rect 14657 4029 14691 4063
rect 14841 4029 14875 4063
rect 15025 4029 15059 4063
rect 15301 4029 15335 4063
rect 15485 4029 15519 4063
rect 15669 4029 15703 4063
rect 15945 4029 15979 4063
rect 16313 4029 16347 4063
rect 17969 4029 18003 4063
rect 18153 4029 18187 4063
rect 18889 4029 18923 4063
rect 23029 4029 23063 4063
rect 4344 3961 4378 3995
rect 7573 3961 7607 3995
rect 9321 3961 9355 3995
rect 13001 3961 13035 3995
rect 13921 3961 13955 3995
rect 14933 3961 14967 3995
rect 15577 3961 15611 3995
rect 16129 3961 16163 3995
rect 16221 3961 16255 3995
rect 19686 3961 19720 3995
rect 3617 3893 3651 3927
rect 6837 3893 6871 3927
rect 8585 3893 8619 3927
rect 10057 3893 10091 3927
rect 11621 3893 11655 3927
rect 14013 3893 14047 3927
rect 15209 3893 15243 3927
rect 16497 3893 16531 3927
rect 18337 3893 18371 3927
rect 18705 3893 18739 3927
rect 20821 3893 20855 3927
rect 5181 3689 5215 3723
rect 7849 3689 7883 3723
rect 10793 3689 10827 3723
rect 12449 3689 12483 3723
rect 13921 3689 13955 3723
rect 14749 3689 14783 3723
rect 18705 3689 18739 3723
rect 18981 3689 19015 3723
rect 4046 3621 4080 3655
rect 6736 3621 6770 3655
rect 11336 3621 11370 3655
rect 14289 3621 14323 3655
rect 19318 3621 19352 3655
rect 3709 3553 3743 3587
rect 3801 3553 3835 3587
rect 6469 3553 6503 3587
rect 8309 3553 8343 3587
rect 8576 3553 8610 3587
rect 11069 3553 11103 3587
rect 12725 3553 12759 3587
rect 14381 3553 14415 3587
rect 15117 3553 15151 3587
rect 16129 3553 16163 3587
rect 16313 3553 16347 3587
rect 16405 3553 16439 3587
rect 16497 3553 16531 3587
rect 17785 3553 17819 3587
rect 17969 3553 18003 3587
rect 18521 3553 18555 3587
rect 18797 3553 18831 3587
rect 19073 3553 19107 3587
rect 10149 3485 10183 3519
rect 12541 3485 12575 3519
rect 14565 3485 14599 3519
rect 15209 3485 15243 3519
rect 15301 3485 15335 3519
rect 3525 3349 3559 3383
rect 9689 3349 9723 3383
rect 12909 3349 12943 3383
rect 16681 3349 16715 3383
rect 18153 3349 18187 3383
rect 20453 3349 20487 3383
rect 4721 3145 4755 3179
rect 10149 3145 10183 3179
rect 15945 3145 15979 3179
rect 20085 3077 20119 3111
rect 3341 3009 3375 3043
rect 15301 3009 15335 3043
rect 17509 3009 17543 3043
rect 18705 3009 18739 3043
rect 3608 2941 3642 2975
rect 5273 2941 5307 2975
rect 5365 2941 5399 2975
rect 5641 2941 5675 2975
rect 5733 2941 5767 2975
rect 5917 2941 5951 2975
rect 6009 2941 6043 2975
rect 6101 2941 6135 2975
rect 7481 2941 7515 2975
rect 7573 2941 7607 2975
rect 7849 2941 7883 2975
rect 8769 2941 8803 2975
rect 12081 2941 12115 2975
rect 12357 2941 12391 2975
rect 12449 2941 12483 2975
rect 12909 2941 12943 2975
rect 15485 2941 15519 2975
rect 16037 2941 16071 2975
rect 16221 2941 16255 2975
rect 16405 2941 16439 2975
rect 16773 2941 16807 2975
rect 16865 2941 16899 2975
rect 17325 2941 17359 2975
rect 18337 2941 18371 2975
rect 5457 2873 5491 2907
rect 7665 2873 7699 2907
rect 9036 2873 9070 2907
rect 12265 2873 12299 2907
rect 15577 2873 15611 2907
rect 16313 2873 16347 2907
rect 18950 2873 18984 2907
rect 5089 2805 5123 2839
rect 6285 2805 6319 2839
rect 7297 2805 7331 2839
rect 12633 2805 12667 2839
rect 12725 2805 12759 2839
rect 16589 2805 16623 2839
rect 17049 2805 17083 2839
rect 17141 2805 17175 2839
rect 18521 2805 18555 2839
rect 5181 2601 5215 2635
rect 9137 2601 9171 2635
rect 13277 2601 13311 2635
rect 14657 2601 14691 2635
rect 5641 2533 5675 2567
rect 9413 2533 9447 2567
rect 10057 2533 10091 2567
rect 12164 2533 12198 2567
rect 14381 2533 14415 2567
rect 16589 2533 16623 2567
rect 3801 2465 3835 2499
rect 4068 2465 4102 2499
rect 5457 2465 5491 2499
rect 6009 2465 6043 2499
rect 6469 2465 6503 2499
rect 7573 2465 7607 2499
rect 8861 2465 8895 2499
rect 9321 2465 9355 2499
rect 9505 2465 9539 2499
rect 9689 2465 9723 2499
rect 9965 2465 9999 2499
rect 10149 2465 10183 2499
rect 10333 2465 10367 2499
rect 14197 2465 14231 2499
rect 14289 2465 14323 2499
rect 14565 2465 14599 2499
rect 15025 2465 15059 2499
rect 16773 2465 16807 2499
rect 17233 2465 17267 2499
rect 5273 2397 5307 2431
rect 6193 2397 6227 2431
rect 7389 2397 7423 2431
rect 8677 2397 8711 2431
rect 11897 2397 11931 2431
rect 15117 2397 15151 2431
rect 15301 2397 15335 2431
rect 16313 2397 16347 2431
rect 5825 2261 5859 2295
rect 6285 2261 6319 2295
rect 7757 2261 7791 2295
rect 9045 2261 9079 2295
rect 9781 2261 9815 2295
rect 14013 2261 14047 2295
rect 16957 2261 16991 2295
rect 17049 2261 17083 2295
rect 4353 2057 4387 2091
rect 11345 2057 11379 2091
rect 15301 1989 15335 2023
rect 6377 1921 6411 1955
rect 9954 1921 9988 1955
rect 14197 1921 14231 1955
rect 20269 1921 20303 1955
rect 4537 1853 4571 1887
rect 6121 1853 6155 1887
rect 7665 1853 7699 1887
rect 8953 1853 8987 1887
rect 9229 1853 9263 1887
rect 9505 1853 9539 1887
rect 9689 1853 9723 1887
rect 9873 1853 9907 1887
rect 12357 1853 12391 1887
rect 12449 1853 12483 1887
rect 12633 1853 12667 1887
rect 12725 1853 12759 1887
rect 13737 1853 13771 1887
rect 13921 1853 13955 1887
rect 14381 1853 14415 1887
rect 14933 1853 14967 1887
rect 15117 1853 15151 1887
rect 15853 1853 15887 1887
rect 17417 1853 17451 1887
rect 19809 1853 19843 1887
rect 19993 1853 20027 1887
rect 20361 1853 20395 1887
rect 10210 1785 10244 1819
rect 14105 1785 14139 1819
rect 17150 1785 17184 1819
rect 21005 1785 21039 1819
rect 4997 1717 5031 1751
rect 7481 1717 7515 1751
rect 9137 1717 9171 1751
rect 9413 1717 9447 1751
rect 12909 1717 12943 1751
rect 15669 1717 15703 1751
rect 16037 1717 16071 1751
rect 5917 1513 5951 1547
rect 8677 1513 8711 1547
rect 10701 1513 10735 1547
rect 12081 1513 12115 1547
rect 18153 1513 18187 1547
rect 22201 1513 22235 1547
rect 9566 1445 9600 1479
rect 11529 1445 11563 1479
rect 13194 1445 13228 1479
rect 17040 1445 17074 1479
rect 18613 1445 18647 1479
rect 18705 1445 18739 1479
rect 19550 1445 19584 1479
rect 20913 1445 20947 1479
rect 4445 1377 4479 1411
rect 4905 1377 4939 1411
rect 5089 1377 5123 1411
rect 5457 1377 5491 1411
rect 6285 1377 6319 1411
rect 6469 1377 6503 1411
rect 6837 1377 6871 1411
rect 7564 1377 7598 1411
rect 11432 1377 11466 1411
rect 11621 1377 11655 1411
rect 11805 1377 11839 1411
rect 14197 1377 14231 1411
rect 14289 1377 14323 1411
rect 14565 1377 14599 1411
rect 15025 1377 15059 1411
rect 15117 1377 15151 1411
rect 18469 1377 18503 1411
rect 18889 1377 18923 1411
rect 18981 1377 19015 1411
rect 19165 1377 19199 1411
rect 19257 1377 19291 1411
rect 19354 1377 19388 1411
rect 19809 1377 19843 1411
rect 19901 1377 19935 1411
rect 20269 1377 20303 1411
rect 21465 1377 21499 1411
rect 21833 1377 21867 1411
rect 22017 1377 22051 1411
rect 5365 1309 5399 1343
rect 6745 1309 6779 1343
rect 7297 1309 7331 1343
rect 9321 1309 9355 1343
rect 13461 1309 13495 1343
rect 14381 1309 14415 1343
rect 16773 1309 16807 1343
rect 20453 1309 20487 1343
rect 21557 1309 21591 1343
rect 11253 1173 11287 1207
rect 15577 1173 15611 1207
rect 18337 1173 18371 1207
rect 14105 969 14139 1003
rect 5917 901 5951 935
rect 8033 901 8067 935
rect 9597 901 9631 935
rect 13093 901 13127 935
rect 16681 901 16715 935
rect 15485 833 15519 867
rect 20177 833 20211 867
rect 6096 765 6130 799
rect 6193 765 6227 799
rect 6285 765 6319 799
rect 6469 765 6503 799
rect 7481 765 7515 799
rect 7901 765 7935 799
rect 9045 765 9079 799
rect 9465 765 9499 799
rect 12541 765 12575 799
rect 12817 765 12851 799
rect 12961 765 12995 799
rect 15229 765 15263 799
rect 16129 765 16163 799
rect 16313 765 16347 799
rect 16405 765 16439 799
rect 16502 765 16536 799
rect 19809 765 19843 799
rect 19901 765 19935 799
rect 20269 765 20303 799
rect 7665 697 7699 731
rect 7757 697 7791 731
rect 9229 697 9263 731
rect 9321 697 9355 731
rect 12725 697 12759 731
rect 20913 697 20947 731
<< metal1 >>
rect 10226 17552 10232 17604
rect 10284 17592 10290 17604
rect 10410 17592 10416 17604
rect 10284 17564 10416 17592
rect 10284 17552 10290 17564
rect 10410 17552 10416 17564
rect 10468 17552 10474 17604
rect 16758 17552 16764 17604
rect 16816 17592 16822 17604
rect 25130 17592 25136 17604
rect 16816 17564 25136 17592
rect 16816 17552 16822 17564
rect 25130 17552 25136 17564
rect 25188 17552 25194 17604
rect 3602 17484 3608 17536
rect 3660 17524 3666 17536
rect 3970 17524 3976 17536
rect 3660 17496 3976 17524
rect 3660 17484 3666 17496
rect 3970 17484 3976 17496
rect 4028 17484 4034 17536
rect 18966 17484 18972 17536
rect 19024 17524 19030 17536
rect 24670 17524 24676 17536
rect 19024 17496 24676 17524
rect 19024 17484 19030 17496
rect 24670 17484 24676 17496
rect 24728 17484 24734 17536
rect 552 17434 27416 17456
rect 552 17382 3756 17434
rect 3808 17382 3820 17434
rect 3872 17382 3884 17434
rect 3936 17382 3948 17434
rect 4000 17382 4012 17434
rect 4064 17382 10472 17434
rect 10524 17382 10536 17434
rect 10588 17382 10600 17434
rect 10652 17382 10664 17434
rect 10716 17382 10728 17434
rect 10780 17382 17188 17434
rect 17240 17382 17252 17434
rect 17304 17382 17316 17434
rect 17368 17382 17380 17434
rect 17432 17382 17444 17434
rect 17496 17382 23904 17434
rect 23956 17382 23968 17434
rect 24020 17382 24032 17434
rect 24084 17382 24096 17434
rect 24148 17382 24160 17434
rect 24212 17382 27416 17434
rect 552 17360 27416 17382
rect 842 17280 848 17332
rect 900 17280 906 17332
rect 1486 17280 1492 17332
rect 1544 17280 1550 17332
rect 3602 17280 3608 17332
rect 3660 17320 3666 17332
rect 4065 17323 4123 17329
rect 4065 17320 4077 17323
rect 3660 17292 4077 17320
rect 3660 17280 3666 17292
rect 4065 17289 4077 17292
rect 4111 17289 4123 17323
rect 4065 17283 4123 17289
rect 5902 17280 5908 17332
rect 5960 17320 5966 17332
rect 5997 17323 6055 17329
rect 5997 17320 6009 17323
rect 5960 17292 6009 17320
rect 5960 17280 5966 17292
rect 5997 17289 6009 17292
rect 6043 17289 6055 17323
rect 5997 17283 6055 17289
rect 6546 17280 6552 17332
rect 6604 17320 6610 17332
rect 6641 17323 6699 17329
rect 6641 17320 6653 17323
rect 6604 17292 6653 17320
rect 6604 17280 6610 17292
rect 6641 17289 6653 17292
rect 6687 17289 6699 17323
rect 6641 17283 6699 17289
rect 8113 17323 8171 17329
rect 8113 17289 8125 17323
rect 8159 17320 8171 17323
rect 8478 17320 8484 17332
rect 8159 17292 8484 17320
rect 8159 17289 8171 17292
rect 8113 17283 8171 17289
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 9122 17280 9128 17332
rect 9180 17320 9186 17332
rect 9217 17323 9275 17329
rect 9217 17320 9229 17323
rect 9180 17292 9229 17320
rect 9180 17280 9186 17292
rect 9217 17289 9229 17292
rect 9263 17289 9275 17323
rect 9217 17283 9275 17289
rect 10226 17280 10232 17332
rect 10284 17320 10290 17332
rect 10597 17323 10655 17329
rect 10597 17320 10609 17323
rect 10284 17292 10609 17320
rect 10284 17280 10290 17292
rect 10597 17289 10609 17292
rect 10643 17289 10655 17323
rect 10597 17283 10655 17289
rect 11698 17280 11704 17332
rect 11756 17320 11762 17332
rect 12069 17323 12127 17329
rect 12069 17320 12081 17323
rect 11756 17292 12081 17320
rect 11756 17280 11762 17292
rect 12069 17289 12081 17292
rect 12115 17289 12127 17323
rect 12069 17283 12127 17289
rect 13630 17280 13636 17332
rect 13688 17320 13694 17332
rect 14185 17323 14243 17329
rect 14185 17320 14197 17323
rect 13688 17292 14197 17320
rect 13688 17280 13694 17292
rect 14185 17289 14197 17292
rect 14231 17289 14243 17323
rect 14185 17283 14243 17289
rect 20346 17280 20352 17332
rect 20404 17320 20410 17332
rect 22741 17323 22799 17329
rect 22741 17320 22753 17323
rect 20404 17292 22753 17320
rect 20404 17280 20410 17292
rect 22741 17289 22753 17292
rect 22787 17289 22799 17323
rect 22741 17283 22799 17289
rect 24670 17280 24676 17332
rect 24728 17280 24734 17332
rect 25130 17280 25136 17332
rect 25188 17280 25194 17332
rect 12158 17212 12164 17264
rect 12216 17252 12222 17264
rect 18325 17255 18383 17261
rect 18325 17252 18337 17255
rect 12216 17224 18337 17252
rect 12216 17212 12222 17224
rect 18325 17221 18337 17224
rect 18371 17221 18383 17255
rect 18325 17215 18383 17221
rect 19058 17212 19064 17264
rect 19116 17252 19122 17264
rect 20714 17252 20720 17264
rect 19116 17224 19748 17252
rect 19116 17212 19122 17224
rect 2682 17144 2688 17196
rect 2740 17184 2746 17196
rect 2777 17187 2835 17193
rect 2777 17184 2789 17187
rect 2740 17156 2789 17184
rect 2740 17144 2746 17156
rect 2777 17153 2789 17156
rect 2823 17153 2835 17187
rect 2777 17147 2835 17153
rect 3418 17144 3424 17196
rect 3476 17144 3482 17196
rect 4706 17144 4712 17196
rect 4764 17144 4770 17196
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 5353 17187 5411 17193
rect 5353 17184 5365 17187
rect 5316 17156 5365 17184
rect 5316 17144 5322 17156
rect 5353 17153 5365 17156
rect 5399 17153 5411 17187
rect 19426 17184 19432 17196
rect 5353 17147 5411 17153
rect 18524 17156 19432 17184
rect 7834 17076 7840 17128
rect 7892 17116 7898 17128
rect 7929 17119 7987 17125
rect 7929 17116 7941 17119
rect 7892 17088 7941 17116
rect 7892 17076 7898 17088
rect 7929 17085 7941 17088
rect 7975 17085 7987 17119
rect 7929 17079 7987 17085
rect 9950 17076 9956 17128
rect 10008 17116 10014 17128
rect 10137 17119 10195 17125
rect 10137 17116 10149 17119
rect 10008 17088 10149 17116
rect 10008 17076 10014 17088
rect 10137 17085 10149 17088
rect 10183 17085 10195 17119
rect 10137 17079 10195 17085
rect 10778 17076 10784 17128
rect 10836 17076 10842 17128
rect 11882 17076 11888 17128
rect 11940 17076 11946 17128
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17116 14427 17119
rect 14550 17116 14556 17128
rect 14415 17088 14556 17116
rect 14415 17085 14427 17088
rect 14369 17079 14427 17085
rect 14550 17076 14556 17088
rect 14608 17076 14614 17128
rect 16482 17076 16488 17128
rect 16540 17076 16546 17128
rect 16850 17076 16856 17128
rect 16908 17116 16914 17128
rect 16945 17119 17003 17125
rect 16945 17116 16957 17119
rect 16908 17088 16957 17116
rect 16908 17076 16914 17088
rect 16945 17085 16957 17088
rect 16991 17085 17003 17119
rect 16945 17079 17003 17085
rect 17770 17076 17776 17128
rect 17828 17076 17834 17128
rect 18524 17125 18552 17156
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 19720 17193 19748 17224
rect 20272 17224 20720 17252
rect 19705 17187 19763 17193
rect 19705 17153 19717 17187
rect 19751 17184 19763 17187
rect 19978 17184 19984 17196
rect 19751 17156 19984 17184
rect 19751 17153 19763 17156
rect 19705 17147 19763 17153
rect 19978 17144 19984 17156
rect 20036 17144 20042 17196
rect 20162 17144 20168 17196
rect 20220 17184 20226 17196
rect 20272 17193 20300 17224
rect 20714 17212 20720 17224
rect 20772 17212 20778 17264
rect 23385 17255 23443 17261
rect 21008 17224 21772 17252
rect 20257 17187 20315 17193
rect 20257 17184 20269 17187
rect 20220 17156 20269 17184
rect 20220 17144 20226 17156
rect 20257 17153 20269 17156
rect 20303 17153 20315 17187
rect 20257 17147 20315 17153
rect 18509 17119 18567 17125
rect 18509 17085 18521 17119
rect 18555 17085 18567 17119
rect 18509 17079 18567 17085
rect 18966 17076 18972 17128
rect 19024 17076 19030 17128
rect 19058 17076 19064 17128
rect 19116 17076 19122 17128
rect 19518 17076 19524 17128
rect 19576 17076 19582 17128
rect 20073 17119 20131 17125
rect 20073 17085 20085 17119
rect 20119 17116 20131 17119
rect 20346 17116 20352 17128
rect 20119 17088 20352 17116
rect 20119 17085 20131 17088
rect 20073 17079 20131 17085
rect 20346 17076 20352 17088
rect 20404 17076 20410 17128
rect 20625 17119 20683 17125
rect 20625 17085 20637 17119
rect 20671 17085 20683 17119
rect 20625 17079 20683 17085
rect 20640 17048 20668 17079
rect 20714 17076 20720 17128
rect 20772 17116 20778 17128
rect 21008 17116 21036 17224
rect 21744 17193 21772 17224
rect 23385 17221 23397 17255
rect 23431 17221 23443 17255
rect 23385 17215 23443 17221
rect 21729 17187 21787 17193
rect 21729 17153 21741 17187
rect 21775 17184 21787 17187
rect 21821 17187 21879 17193
rect 21821 17184 21833 17187
rect 21775 17156 21833 17184
rect 21775 17153 21787 17156
rect 21729 17147 21787 17153
rect 21821 17153 21833 17156
rect 21867 17153 21879 17187
rect 23400 17184 23428 17215
rect 24026 17212 24032 17264
rect 24084 17212 24090 17264
rect 21821 17147 21879 17153
rect 22020 17156 23428 17184
rect 25409 17187 25467 17193
rect 20772 17088 21036 17116
rect 21085 17119 21143 17125
rect 20772 17076 20778 17088
rect 21085 17085 21097 17119
rect 21131 17116 21143 17119
rect 21358 17116 21364 17128
rect 21131 17088 21364 17116
rect 21131 17085 21143 17088
rect 21085 17079 21143 17085
rect 21358 17076 21364 17088
rect 21416 17076 21422 17128
rect 22020 17125 22048 17156
rect 25409 17153 25421 17187
rect 25455 17184 25467 17187
rect 25866 17184 25872 17196
rect 25455 17156 25872 17184
rect 25455 17153 25467 17156
rect 25409 17147 25467 17153
rect 25866 17144 25872 17156
rect 25924 17144 25930 17196
rect 21545 17119 21603 17125
rect 21545 17085 21557 17119
rect 21591 17085 21603 17119
rect 21545 17079 21603 17085
rect 22005 17119 22063 17125
rect 22005 17085 22017 17119
rect 22051 17085 22063 17119
rect 22005 17079 22063 17085
rect 17144 17020 17816 17048
rect 20640 17020 20944 17048
rect 9398 16940 9404 16992
rect 9456 16980 9462 16992
rect 9585 16983 9643 16989
rect 9585 16980 9597 16983
rect 9456 16952 9597 16980
rect 9456 16940 9462 16952
rect 9585 16949 9597 16952
rect 9631 16949 9643 16983
rect 9585 16943 9643 16949
rect 15102 16940 15108 16992
rect 15160 16980 15166 16992
rect 17144 16989 17172 17020
rect 17788 16992 17816 17020
rect 16301 16983 16359 16989
rect 16301 16980 16313 16983
rect 15160 16952 16313 16980
rect 15160 16940 15166 16952
rect 16301 16949 16313 16952
rect 16347 16949 16359 16983
rect 16301 16943 16359 16949
rect 17129 16983 17187 16989
rect 17129 16949 17141 16983
rect 17175 16949 17187 16983
rect 17129 16943 17187 16949
rect 17586 16940 17592 16992
rect 17644 16940 17650 16992
rect 17770 16940 17776 16992
rect 17828 16940 17834 16992
rect 18414 16940 18420 16992
rect 18472 16980 18478 16992
rect 18785 16983 18843 16989
rect 18785 16980 18797 16983
rect 18472 16952 18797 16980
rect 18472 16940 18478 16952
rect 18785 16949 18797 16952
rect 18831 16949 18843 16983
rect 18785 16943 18843 16949
rect 19334 16940 19340 16992
rect 19392 16940 19398 16992
rect 19886 16940 19892 16992
rect 19944 16940 19950 16992
rect 19978 16940 19984 16992
rect 20036 16980 20042 16992
rect 20916 16989 20944 17020
rect 20441 16983 20499 16989
rect 20441 16980 20453 16983
rect 20036 16952 20453 16980
rect 20036 16940 20042 16952
rect 20441 16949 20453 16952
rect 20487 16949 20499 16983
rect 20441 16943 20499 16949
rect 20901 16983 20959 16989
rect 20901 16949 20913 16983
rect 20947 16949 20959 16983
rect 20901 16943 20959 16949
rect 21361 16983 21419 16989
rect 21361 16949 21373 16983
rect 21407 16980 21419 16983
rect 21450 16980 21456 16992
rect 21407 16952 21456 16980
rect 21407 16949 21419 16952
rect 21361 16943 21419 16949
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 21560 16980 21588 17079
rect 22278 17076 22284 17128
rect 22336 17116 22342 17128
rect 22557 17119 22615 17125
rect 22557 17116 22569 17119
rect 22336 17088 22569 17116
rect 22336 17076 22342 17088
rect 22557 17085 22569 17088
rect 22603 17085 22615 17119
rect 22557 17079 22615 17085
rect 22646 17076 22652 17128
rect 22704 17116 22710 17128
rect 22925 17119 22983 17125
rect 22925 17116 22937 17119
rect 22704 17088 22937 17116
rect 22704 17076 22710 17088
rect 22925 17085 22937 17088
rect 22971 17085 22983 17119
rect 22925 17079 22983 17085
rect 23290 17076 23296 17128
rect 23348 17116 23354 17128
rect 23569 17119 23627 17125
rect 23569 17116 23581 17119
rect 23348 17088 23581 17116
rect 23348 17076 23354 17088
rect 23569 17085 23581 17088
rect 23615 17085 23627 17119
rect 23569 17079 23627 17085
rect 23750 17076 23756 17128
rect 23808 17116 23814 17128
rect 24213 17119 24271 17125
rect 24213 17116 24225 17119
rect 23808 17088 24225 17116
rect 23808 17076 23814 17088
rect 24213 17085 24225 17088
rect 24259 17085 24271 17119
rect 24213 17079 24271 17085
rect 24578 17076 24584 17128
rect 24636 17116 24642 17128
rect 24857 17119 24915 17125
rect 24857 17116 24869 17119
rect 24636 17088 24869 17116
rect 24636 17076 24642 17088
rect 24857 17085 24869 17088
rect 24903 17085 24915 17119
rect 24857 17079 24915 17085
rect 25222 17076 25228 17128
rect 25280 17116 25286 17128
rect 25317 17119 25375 17125
rect 25317 17116 25329 17119
rect 25280 17088 25329 17116
rect 25280 17076 25286 17088
rect 25317 17085 25329 17088
rect 25363 17085 25375 17119
rect 25317 17079 25375 17085
rect 25498 17076 25504 17128
rect 25556 17116 25562 17128
rect 25685 17119 25743 17125
rect 25685 17116 25697 17119
rect 25556 17088 25697 17116
rect 25556 17076 25562 17088
rect 25685 17085 25697 17088
rect 25731 17085 25743 17119
rect 25685 17079 25743 17085
rect 26326 17076 26332 17128
rect 26384 17116 26390 17128
rect 26421 17119 26479 17125
rect 26421 17116 26433 17119
rect 26384 17088 26433 17116
rect 26384 17076 26390 17088
rect 26421 17085 26433 17088
rect 26467 17085 26479 17119
rect 26421 17079 26479 17085
rect 22189 17051 22247 17057
rect 22189 17017 22201 17051
rect 22235 17048 22247 17051
rect 22235 17020 22968 17048
rect 22235 17017 22247 17020
rect 22189 17011 22247 17017
rect 22373 16983 22431 16989
rect 22373 16980 22385 16983
rect 21560 16952 22385 16980
rect 22373 16949 22385 16952
rect 22419 16949 22431 16983
rect 22940 16980 22968 17020
rect 24118 17008 24124 17060
rect 24176 17048 24182 17060
rect 24670 17048 24676 17060
rect 24176 17020 24676 17048
rect 24176 17008 24182 17020
rect 24670 17008 24676 17020
rect 24728 17048 24734 17060
rect 26970 17048 26976 17060
rect 24728 17020 26976 17048
rect 24728 17008 24734 17020
rect 26970 17008 26976 17020
rect 27028 17008 27034 17060
rect 23106 16980 23112 16992
rect 22940 16952 23112 16980
rect 22373 16943 22431 16949
rect 23106 16940 23112 16952
rect 23164 16940 23170 16992
rect 26694 16940 26700 16992
rect 26752 16980 26758 16992
rect 27065 16983 27123 16989
rect 27065 16980 27077 16983
rect 26752 16952 27077 16980
rect 26752 16940 26758 16952
rect 27065 16949 27077 16952
rect 27111 16949 27123 16983
rect 27065 16943 27123 16949
rect 552 16890 27576 16912
rect 552 16838 7114 16890
rect 7166 16838 7178 16890
rect 7230 16838 7242 16890
rect 7294 16838 7306 16890
rect 7358 16838 7370 16890
rect 7422 16838 13830 16890
rect 13882 16838 13894 16890
rect 13946 16838 13958 16890
rect 14010 16838 14022 16890
rect 14074 16838 14086 16890
rect 14138 16838 20546 16890
rect 20598 16838 20610 16890
rect 20662 16838 20674 16890
rect 20726 16838 20738 16890
rect 20790 16838 20802 16890
rect 20854 16838 27262 16890
rect 27314 16838 27326 16890
rect 27378 16838 27390 16890
rect 27442 16838 27454 16890
rect 27506 16838 27518 16890
rect 27570 16838 27576 16890
rect 552 16816 27576 16838
rect 7929 16779 7987 16785
rect 7929 16745 7941 16779
rect 7975 16745 7987 16779
rect 9674 16776 9680 16788
rect 7929 16739 7987 16745
rect 8128 16748 9680 16776
rect 6724 16711 6782 16717
rect 6724 16677 6736 16711
rect 6770 16708 6782 16711
rect 7944 16708 7972 16739
rect 6770 16680 7972 16708
rect 6770 16677 6782 16680
rect 6724 16671 6782 16677
rect 8128 16649 8156 16748
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 9766 16736 9772 16788
rect 9824 16736 9830 16788
rect 10778 16736 10784 16788
rect 10836 16776 10842 16788
rect 10965 16779 11023 16785
rect 10965 16776 10977 16779
rect 10836 16748 10977 16776
rect 10836 16736 10842 16748
rect 10965 16745 10977 16748
rect 11011 16745 11023 16779
rect 10965 16739 11023 16745
rect 12805 16779 12863 16785
rect 12805 16745 12817 16779
rect 12851 16776 12863 16779
rect 12986 16776 12992 16788
rect 12851 16748 12992 16776
rect 12851 16745 12863 16748
rect 12805 16739 12863 16745
rect 12986 16736 12992 16748
rect 13044 16736 13050 16788
rect 13633 16779 13691 16785
rect 13633 16776 13645 16779
rect 13464 16748 13645 16776
rect 8220 16680 12388 16708
rect 8220 16649 8248 16680
rect 12360 16652 12388 16680
rect 12710 16668 12716 16720
rect 12768 16708 12774 16720
rect 13464 16717 13492 16748
rect 13633 16745 13645 16748
rect 13679 16745 13691 16779
rect 13633 16739 13691 16745
rect 14274 16736 14280 16788
rect 14332 16776 14338 16788
rect 15473 16779 15531 16785
rect 15473 16776 15485 16779
rect 14332 16748 15485 16776
rect 14332 16736 14338 16748
rect 15473 16745 15485 16748
rect 15519 16745 15531 16779
rect 15473 16739 15531 16745
rect 15838 16736 15844 16788
rect 15896 16736 15902 16788
rect 19794 16736 19800 16788
rect 19852 16776 19858 16788
rect 24118 16776 24124 16788
rect 19852 16748 24124 16776
rect 19852 16736 19858 16748
rect 13081 16711 13139 16717
rect 13081 16708 13093 16711
rect 12768 16680 13093 16708
rect 12768 16668 12774 16680
rect 13081 16677 13093 16680
rect 13127 16677 13139 16711
rect 13081 16671 13139 16677
rect 13449 16711 13507 16717
rect 13449 16677 13461 16711
rect 13495 16677 13507 16711
rect 14829 16711 14887 16717
rect 14829 16708 14841 16711
rect 13449 16671 13507 16677
rect 14016 16680 14841 16708
rect 14016 16652 14044 16680
rect 14829 16677 14841 16680
rect 14875 16677 14887 16711
rect 14829 16671 14887 16677
rect 15013 16711 15071 16717
rect 15013 16677 15025 16711
rect 15059 16708 15071 16711
rect 17586 16708 17592 16720
rect 15059 16680 17592 16708
rect 15059 16677 15071 16680
rect 15013 16671 15071 16677
rect 17586 16668 17592 16680
rect 17644 16668 17650 16720
rect 19245 16711 19303 16717
rect 19245 16677 19257 16711
rect 19291 16708 19303 16711
rect 20714 16708 20720 16720
rect 19291 16680 20720 16708
rect 19291 16677 19303 16680
rect 19245 16671 19303 16677
rect 20714 16668 20720 16680
rect 20772 16668 20778 16720
rect 23032 16708 23060 16748
rect 24118 16736 24124 16748
rect 24176 16736 24182 16788
rect 25958 16776 25964 16788
rect 24412 16748 25964 16776
rect 24412 16708 24440 16748
rect 25958 16736 25964 16748
rect 26016 16776 26022 16788
rect 26016 16748 26832 16776
rect 26016 16736 26022 16748
rect 22480 16680 22784 16708
rect 8478 16649 8484 16652
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16609 8171 16643
rect 8113 16603 8171 16609
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16609 8263 16643
rect 8205 16603 8263 16609
rect 8472 16603 8484 16649
rect 8478 16600 8484 16603
rect 8536 16600 8542 16652
rect 9950 16640 9956 16652
rect 9600 16612 9956 16640
rect 5810 16532 5816 16584
rect 5868 16572 5874 16584
rect 6457 16575 6515 16581
rect 6457 16572 6469 16575
rect 5868 16544 6469 16572
rect 5868 16532 5874 16544
rect 6457 16541 6469 16544
rect 6503 16541 6515 16575
rect 6457 16535 6515 16541
rect 9600 16513 9628 16612
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10778 16600 10784 16652
rect 10836 16600 10842 16652
rect 11146 16600 11152 16652
rect 11204 16640 11210 16652
rect 12078 16643 12136 16649
rect 12078 16640 12090 16643
rect 11204 16612 12090 16640
rect 11204 16600 11210 16612
rect 12078 16609 12090 16612
rect 12124 16609 12136 16643
rect 12078 16603 12136 16609
rect 12342 16600 12348 16652
rect 12400 16600 12406 16652
rect 12986 16600 12992 16652
rect 13044 16600 13050 16652
rect 13998 16600 14004 16652
rect 14056 16600 14062 16652
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16640 14151 16643
rect 14274 16640 14280 16652
rect 14139 16612 14280 16640
rect 14139 16609 14151 16612
rect 14093 16603 14151 16609
rect 14274 16600 14280 16612
rect 14332 16600 14338 16652
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15289 16643 15347 16649
rect 15289 16640 15301 16643
rect 15252 16612 15301 16640
rect 15252 16600 15258 16612
rect 15289 16609 15301 16612
rect 15335 16609 15347 16643
rect 15289 16603 15347 16609
rect 15562 16600 15568 16652
rect 15620 16640 15626 16652
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 15620 16612 15669 16640
rect 15620 16600 15626 16612
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 15657 16603 15715 16609
rect 16574 16600 16580 16652
rect 16632 16600 16638 16652
rect 16758 16600 16764 16652
rect 16816 16600 16822 16652
rect 19058 16640 19064 16652
rect 18432 16612 19064 16640
rect 14185 16575 14243 16581
rect 14185 16541 14197 16575
rect 14231 16572 14243 16575
rect 14826 16572 14832 16584
rect 14231 16544 14832 16572
rect 14231 16541 14243 16544
rect 14185 16535 14243 16541
rect 14826 16532 14832 16544
rect 14884 16532 14890 16584
rect 15102 16532 15108 16584
rect 15160 16532 15166 16584
rect 16945 16575 17003 16581
rect 16945 16541 16957 16575
rect 16991 16572 17003 16575
rect 18432 16572 18460 16612
rect 19058 16600 19064 16612
rect 19116 16600 19122 16652
rect 19521 16643 19579 16649
rect 19521 16609 19533 16643
rect 19567 16609 19579 16643
rect 19521 16603 19579 16609
rect 16991 16544 18460 16572
rect 16991 16541 17003 16544
rect 16945 16535 17003 16541
rect 9585 16507 9643 16513
rect 9585 16473 9597 16507
rect 9631 16473 9643 16507
rect 14844 16504 14872 16532
rect 16960 16504 16988 16535
rect 18506 16532 18512 16584
rect 18564 16532 18570 16584
rect 14844 16476 16988 16504
rect 19536 16504 19564 16603
rect 19610 16600 19616 16652
rect 19668 16600 19674 16652
rect 19705 16643 19763 16649
rect 19705 16609 19717 16643
rect 19751 16609 19763 16643
rect 19705 16603 19763 16609
rect 19720 16572 19748 16603
rect 19794 16600 19800 16652
rect 19852 16640 19858 16652
rect 22480 16649 22508 16680
rect 19889 16643 19947 16649
rect 19889 16640 19901 16643
rect 19852 16612 19901 16640
rect 19852 16600 19858 16612
rect 19889 16609 19901 16612
rect 19935 16609 19947 16643
rect 22097 16643 22155 16649
rect 22465 16643 22523 16649
rect 19889 16603 19947 16609
rect 19996 16612 22048 16640
rect 19996 16572 20024 16612
rect 19720 16544 20024 16572
rect 20625 16575 20683 16581
rect 20625 16541 20637 16575
rect 20671 16572 20683 16575
rect 20898 16572 20904 16584
rect 20671 16544 20904 16572
rect 20671 16541 20683 16544
rect 20625 16535 20683 16541
rect 20898 16532 20904 16544
rect 20956 16532 20962 16584
rect 22020 16572 22048 16612
rect 22097 16609 22109 16643
rect 22143 16615 22232 16643
rect 22143 16609 22155 16615
rect 22097 16603 22155 16609
rect 22204 16581 22232 16615
rect 22465 16609 22477 16643
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16609 22615 16643
rect 22557 16603 22615 16609
rect 22189 16575 22247 16581
rect 22020 16544 22094 16572
rect 22066 16516 22094 16544
rect 22189 16541 22201 16575
rect 22235 16541 22247 16575
rect 22572 16572 22600 16603
rect 22646 16600 22652 16652
rect 22704 16600 22710 16652
rect 22189 16535 22247 16541
rect 22388 16544 22600 16572
rect 22756 16572 22784 16680
rect 22940 16680 23060 16708
rect 24044 16680 24440 16708
rect 22833 16643 22891 16649
rect 22833 16609 22845 16643
rect 22879 16640 22891 16643
rect 22940 16640 22968 16680
rect 24044 16640 24072 16680
rect 22879 16612 22968 16640
rect 23032 16612 24072 16640
rect 22879 16609 22891 16612
rect 22833 16603 22891 16609
rect 22756 16544 22968 16572
rect 19981 16507 20039 16513
rect 19981 16504 19993 16507
rect 19536 16476 19993 16504
rect 9585 16467 9643 16473
rect 19981 16473 19993 16476
rect 20027 16473 20039 16507
rect 19981 16467 20039 16473
rect 20088 16476 21588 16504
rect 22066 16476 22100 16516
rect 7834 16396 7840 16448
rect 7892 16396 7898 16448
rect 10134 16396 10140 16448
rect 10192 16396 10198 16448
rect 13354 16396 13360 16448
rect 13412 16436 13418 16448
rect 14553 16439 14611 16445
rect 14553 16436 14565 16439
rect 13412 16408 14565 16436
rect 13412 16396 13418 16408
rect 14553 16405 14565 16408
rect 14599 16405 14611 16439
rect 14553 16399 14611 16405
rect 19058 16396 19064 16448
rect 19116 16396 19122 16448
rect 19610 16396 19616 16448
rect 19668 16436 19674 16448
rect 20088 16436 20116 16476
rect 19668 16408 20116 16436
rect 19668 16396 19674 16408
rect 21358 16396 21364 16448
rect 21416 16436 21422 16448
rect 21453 16439 21511 16445
rect 21453 16436 21465 16439
rect 21416 16408 21465 16436
rect 21416 16396 21422 16408
rect 21453 16405 21465 16408
rect 21499 16405 21511 16439
rect 21560 16436 21588 16476
rect 22094 16464 22100 16476
rect 22152 16464 22158 16516
rect 22388 16436 22416 16544
rect 22940 16513 22968 16544
rect 22925 16507 22983 16513
rect 22925 16473 22937 16507
rect 22971 16473 22983 16507
rect 22925 16467 22983 16473
rect 23032 16436 23060 16612
rect 24118 16600 24124 16652
rect 24176 16600 24182 16652
rect 24302 16600 24308 16652
rect 24360 16600 24366 16652
rect 24412 16649 24440 16680
rect 24765 16711 24823 16717
rect 24765 16677 24777 16711
rect 24811 16708 24823 16711
rect 24811 16680 25544 16708
rect 24811 16677 24823 16680
rect 24765 16671 24823 16677
rect 24397 16643 24455 16649
rect 24397 16609 24409 16643
rect 24443 16609 24455 16643
rect 24397 16603 24455 16609
rect 24489 16643 24547 16649
rect 24489 16609 24501 16643
rect 24535 16640 24547 16643
rect 25314 16640 25320 16652
rect 24535 16612 25320 16640
rect 24535 16609 24547 16612
rect 24489 16603 24547 16609
rect 25314 16600 25320 16612
rect 25372 16600 25378 16652
rect 25516 16649 25544 16680
rect 25590 16668 25596 16720
rect 25648 16708 25654 16720
rect 26421 16711 26479 16717
rect 26421 16708 26433 16711
rect 25648 16680 26433 16708
rect 25648 16668 25654 16680
rect 26421 16677 26433 16680
rect 26467 16677 26479 16711
rect 26421 16671 26479 16677
rect 25501 16643 25559 16649
rect 25501 16609 25513 16643
rect 25547 16609 25559 16643
rect 25501 16603 25559 16609
rect 26234 16600 26240 16652
rect 26292 16600 26298 16652
rect 26694 16600 26700 16652
rect 26752 16600 26758 16652
rect 26804 16649 26832 16748
rect 26789 16643 26847 16649
rect 26789 16609 26801 16643
rect 26835 16609 26847 16643
rect 26789 16603 26847 16609
rect 26878 16600 26884 16652
rect 26936 16600 26942 16652
rect 26970 16600 26976 16652
rect 27028 16640 27034 16652
rect 27065 16643 27123 16649
rect 27065 16640 27077 16643
rect 27028 16612 27077 16640
rect 27028 16600 27034 16612
rect 27065 16609 27077 16612
rect 27111 16609 27123 16643
rect 27065 16603 27123 16609
rect 23474 16532 23480 16584
rect 23532 16532 23538 16584
rect 21560 16408 23060 16436
rect 21453 16399 21511 16405
rect 24946 16396 24952 16448
rect 25004 16396 25010 16448
rect 25682 16396 25688 16448
rect 25740 16436 25746 16448
rect 26053 16439 26111 16445
rect 26053 16436 26065 16439
rect 25740 16408 26065 16436
rect 25740 16396 25746 16408
rect 26053 16405 26065 16408
rect 26099 16405 26111 16439
rect 26053 16399 26111 16405
rect 552 16346 27416 16368
rect 552 16294 3756 16346
rect 3808 16294 3820 16346
rect 3872 16294 3884 16346
rect 3936 16294 3948 16346
rect 4000 16294 4012 16346
rect 4064 16294 10472 16346
rect 10524 16294 10536 16346
rect 10588 16294 10600 16346
rect 10652 16294 10664 16346
rect 10716 16294 10728 16346
rect 10780 16294 17188 16346
rect 17240 16294 17252 16346
rect 17304 16294 17316 16346
rect 17368 16294 17380 16346
rect 17432 16294 17444 16346
rect 17496 16294 23904 16346
rect 23956 16294 23968 16346
rect 24020 16294 24032 16346
rect 24084 16294 24096 16346
rect 24148 16294 24160 16346
rect 24212 16294 27416 16346
rect 552 16272 27416 16294
rect 7101 16235 7159 16241
rect 7101 16201 7113 16235
rect 7147 16232 7159 16235
rect 7466 16232 7472 16244
rect 7147 16204 7472 16232
rect 7147 16201 7159 16204
rect 7101 16195 7159 16201
rect 7466 16192 7472 16204
rect 7524 16192 7530 16244
rect 8478 16192 8484 16244
rect 8536 16192 8542 16244
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 10137 16235 10195 16241
rect 10137 16232 10149 16235
rect 9732 16204 10149 16232
rect 9732 16192 9738 16204
rect 10137 16201 10149 16204
rect 10183 16201 10195 16235
rect 10137 16195 10195 16201
rect 10318 16192 10324 16244
rect 10376 16192 10382 16244
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11517 16235 11575 16241
rect 11517 16232 11529 16235
rect 11112 16204 11529 16232
rect 11112 16192 11118 16204
rect 11517 16201 11529 16204
rect 11563 16201 11575 16235
rect 11517 16195 11575 16201
rect 12069 16235 12127 16241
rect 12069 16201 12081 16235
rect 12115 16232 12127 16235
rect 12250 16232 12256 16244
rect 12115 16204 12256 16232
rect 12115 16201 12127 16204
rect 12069 16195 12127 16201
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 14461 16235 14519 16241
rect 14461 16201 14473 16235
rect 14507 16232 14519 16235
rect 14918 16232 14924 16244
rect 14507 16204 14924 16232
rect 14507 16201 14519 16204
rect 14461 16195 14519 16201
rect 14918 16192 14924 16204
rect 14976 16192 14982 16244
rect 22557 16235 22615 16241
rect 22557 16201 22569 16235
rect 22603 16232 22615 16235
rect 22646 16232 22652 16244
rect 22603 16204 22652 16232
rect 22603 16201 22615 16204
rect 22557 16195 22615 16201
rect 22646 16192 22652 16204
rect 22704 16192 22710 16244
rect 23584 16204 25268 16232
rect 6454 16124 6460 16176
rect 6512 16124 6518 16176
rect 10045 16167 10103 16173
rect 10045 16133 10057 16167
rect 10091 16164 10103 16167
rect 10965 16167 11023 16173
rect 10965 16164 10977 16167
rect 10091 16136 10977 16164
rect 10091 16133 10103 16136
rect 10045 16127 10103 16133
rect 10965 16133 10977 16136
rect 11011 16133 11023 16167
rect 13357 16167 13415 16173
rect 13357 16164 13369 16167
rect 10965 16127 11023 16133
rect 11072 16136 13369 16164
rect 9217 16099 9275 16105
rect 9217 16096 9229 16099
rect 8956 16068 9229 16096
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 16028 6975 16031
rect 7558 16028 7564 16040
rect 6963 16000 7564 16028
rect 6963 15997 6975 16000
rect 6917 15991 6975 15997
rect 7558 15988 7564 16000
rect 7616 15988 7622 16040
rect 8754 15988 8760 16040
rect 8812 15988 8818 16040
rect 8846 15988 8852 16040
rect 8904 15988 8910 16040
rect 8956 16037 8984 16068
rect 9217 16065 9229 16068
rect 9263 16065 9275 16099
rect 10505 16099 10563 16105
rect 10505 16096 10517 16099
rect 9217 16059 9275 16065
rect 9784 16068 10517 16096
rect 8941 16031 8999 16037
rect 8941 15997 8953 16031
rect 8987 15997 8999 16031
rect 8941 15991 8999 15997
rect 9125 16031 9183 16037
rect 9125 15997 9137 16031
rect 9171 15997 9183 16031
rect 9125 15991 9183 15997
rect 6730 15920 6736 15972
rect 6788 15960 6794 15972
rect 6825 15963 6883 15969
rect 6825 15960 6837 15963
rect 6788 15932 6837 15960
rect 6788 15920 6794 15932
rect 6825 15929 6837 15932
rect 6871 15960 6883 15963
rect 7650 15960 7656 15972
rect 6871 15932 7656 15960
rect 6871 15929 6883 15932
rect 6825 15923 6883 15929
rect 7650 15920 7656 15932
rect 7708 15920 7714 15972
rect 7834 15920 7840 15972
rect 7892 15920 7898 15972
rect 8662 15920 8668 15972
rect 8720 15960 8726 15972
rect 9140 15960 9168 15991
rect 9398 15988 9404 16040
rect 9456 15988 9462 16040
rect 9674 15988 9680 16040
rect 9732 15988 9738 16040
rect 9784 16037 9812 16068
rect 10505 16065 10517 16068
rect 10551 16096 10563 16099
rect 11072 16096 11100 16136
rect 13357 16133 13369 16136
rect 13403 16133 13415 16167
rect 13357 16127 13415 16133
rect 22465 16167 22523 16173
rect 22465 16133 22477 16167
rect 22511 16164 22523 16167
rect 23474 16164 23480 16176
rect 22511 16136 23480 16164
rect 22511 16133 22523 16136
rect 22465 16127 22523 16133
rect 23474 16124 23480 16136
rect 23532 16124 23538 16176
rect 10551 16068 11100 16096
rect 11149 16099 11207 16105
rect 10551 16065 10563 16068
rect 10505 16059 10563 16065
rect 11149 16065 11161 16099
rect 11195 16065 11207 16099
rect 11149 16059 11207 16065
rect 9769 16031 9827 16037
rect 9769 15997 9781 16031
rect 9815 15997 9827 16031
rect 9769 15991 9827 15997
rect 10045 16031 10103 16037
rect 10045 15997 10057 16031
rect 10091 16028 10103 16031
rect 10134 16028 10140 16040
rect 10091 16000 10140 16028
rect 10091 15997 10103 16000
rect 10045 15991 10103 15997
rect 10134 15988 10140 16000
rect 10192 16028 10198 16040
rect 10321 16031 10379 16037
rect 10321 16028 10333 16031
rect 10192 16000 10333 16028
rect 10192 15988 10198 16000
rect 10321 15997 10333 16000
rect 10367 15997 10379 16031
rect 10321 15991 10379 15997
rect 10870 15988 10876 16040
rect 10928 15988 10934 16040
rect 11054 15988 11060 16040
rect 11112 16028 11118 16040
rect 11164 16028 11192 16059
rect 11238 16056 11244 16108
rect 11296 16096 11302 16108
rect 11296 16068 12296 16096
rect 11296 16056 11302 16068
rect 11112 16000 11468 16028
rect 11112 15988 11118 16000
rect 10781 15963 10839 15969
rect 10781 15960 10793 15963
rect 8720 15932 9168 15960
rect 9692 15932 10793 15960
rect 8720 15920 8726 15932
rect 9692 15904 9720 15932
rect 10781 15929 10793 15932
rect 10827 15929 10839 15963
rect 10781 15923 10839 15929
rect 11146 15920 11152 15972
rect 11204 15920 11210 15972
rect 6365 15895 6423 15901
rect 6365 15861 6377 15895
rect 6411 15892 6423 15895
rect 7466 15892 7472 15904
rect 6411 15864 7472 15892
rect 6411 15861 6423 15864
rect 6365 15855 6423 15861
rect 7466 15852 7472 15864
rect 7524 15852 7530 15904
rect 9585 15895 9643 15901
rect 9585 15861 9597 15895
rect 9631 15892 9643 15895
rect 9674 15892 9680 15904
rect 9631 15864 9680 15892
rect 9631 15861 9643 15864
rect 9585 15855 9643 15861
rect 9674 15852 9680 15864
rect 9732 15852 9738 15904
rect 9861 15895 9919 15901
rect 9861 15861 9873 15895
rect 9907 15892 9919 15895
rect 10134 15892 10140 15904
rect 9907 15864 10140 15892
rect 9907 15861 9919 15864
rect 9861 15855 9919 15861
rect 10134 15852 10140 15864
rect 10192 15892 10198 15904
rect 10962 15892 10968 15904
rect 10192 15864 10968 15892
rect 10192 15852 10198 15864
rect 10962 15852 10968 15864
rect 11020 15852 11026 15904
rect 11440 15892 11468 16000
rect 11514 15988 11520 16040
rect 11572 16028 11578 16040
rect 12268 16037 12296 16068
rect 20714 16056 20720 16108
rect 20772 16056 20778 16108
rect 22922 16056 22928 16108
rect 22980 16096 22986 16108
rect 23584 16096 23612 16204
rect 25240 16164 25268 16204
rect 25314 16192 25320 16244
rect 25372 16192 25378 16244
rect 25682 16164 25688 16176
rect 25240 16136 25688 16164
rect 25682 16124 25688 16136
rect 25740 16124 25746 16176
rect 22980 16068 23244 16096
rect 22980 16056 22986 16068
rect 11701 16031 11759 16037
rect 11701 16028 11713 16031
rect 11572 16000 11713 16028
rect 11572 15988 11578 16000
rect 11701 15997 11713 16000
rect 11747 15997 11759 16031
rect 11701 15991 11759 15997
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 15997 12311 16031
rect 12253 15991 12311 15997
rect 12434 15988 12440 16040
rect 12492 15988 12498 16040
rect 12618 15988 12624 16040
rect 12676 16028 12682 16040
rect 13173 16031 13231 16037
rect 13173 16028 13185 16031
rect 12676 16000 13185 16028
rect 12676 15988 12682 16000
rect 13173 15997 13185 16000
rect 13219 15997 13231 16031
rect 13173 15991 13231 15997
rect 13354 15988 13360 16040
rect 13412 15988 13418 16040
rect 14185 16031 14243 16037
rect 14185 15997 14197 16031
rect 14231 16028 14243 16031
rect 14274 16028 14280 16040
rect 14231 16000 14280 16028
rect 14231 15997 14243 16000
rect 14185 15991 14243 15997
rect 14274 15988 14280 16000
rect 14332 15988 14338 16040
rect 14642 15988 14648 16040
rect 14700 15988 14706 16040
rect 14734 15988 14740 16040
rect 14792 16028 14798 16040
rect 15102 16028 15108 16040
rect 14792 16000 15108 16028
rect 14792 15988 14798 16000
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 17034 15988 17040 16040
rect 17092 16028 17098 16040
rect 17221 16031 17279 16037
rect 17221 16028 17233 16031
rect 17092 16000 17233 16028
rect 17092 15988 17098 16000
rect 17221 15997 17233 16000
rect 17267 15997 17279 16031
rect 17221 15991 17279 15997
rect 18322 15988 18328 16040
rect 18380 16028 18386 16040
rect 18693 16031 18751 16037
rect 18693 16028 18705 16031
rect 18380 16000 18705 16028
rect 18380 15988 18386 16000
rect 18693 15997 18705 16000
rect 18739 15997 18751 16031
rect 18693 15991 18751 15997
rect 21082 15988 21088 16040
rect 21140 15988 21146 16040
rect 21358 16037 21364 16040
rect 21352 16028 21364 16037
rect 21319 16000 21364 16028
rect 21352 15991 21364 16000
rect 21358 15988 21364 15991
rect 21416 15988 21422 16040
rect 22278 15988 22284 16040
rect 22336 16028 22342 16040
rect 23216 16037 23244 16068
rect 23400 16068 23612 16096
rect 23400 16037 23428 16068
rect 22695 16031 22753 16037
rect 22695 16028 22707 16031
rect 22336 16000 22707 16028
rect 22336 15988 22342 16000
rect 22695 15997 22707 16000
rect 22741 15997 22753 16031
rect 22695 15991 22753 15997
rect 22833 16031 22891 16037
rect 22833 15997 22845 16031
rect 22879 15997 22891 16031
rect 22833 15991 22891 15997
rect 23108 16031 23166 16037
rect 23108 15997 23120 16031
rect 23154 15997 23166 16031
rect 23108 15991 23166 15997
rect 23201 16031 23259 16037
rect 23201 15997 23213 16031
rect 23247 15997 23259 16031
rect 23201 15991 23259 15997
rect 23385 16031 23443 16037
rect 23385 15997 23397 16031
rect 23431 15997 23443 16031
rect 23385 15991 23443 15997
rect 23477 16031 23535 16037
rect 23477 15997 23489 16031
rect 23523 16028 23535 16031
rect 24578 16028 24584 16040
rect 23523 16000 24584 16028
rect 23523 15997 23535 16000
rect 23477 15991 23535 15997
rect 11790 15920 11796 15972
rect 11848 15960 11854 15972
rect 13541 15963 13599 15969
rect 13541 15960 13553 15963
rect 11848 15932 13553 15960
rect 11848 15920 11854 15932
rect 13541 15929 13553 15932
rect 13587 15929 13599 15963
rect 13541 15923 13599 15929
rect 18960 15963 19018 15969
rect 18960 15929 18972 15963
rect 19006 15960 19018 15963
rect 20165 15963 20223 15969
rect 20165 15960 20177 15963
rect 19006 15932 20177 15960
rect 19006 15929 19018 15932
rect 18960 15923 19018 15929
rect 20165 15929 20177 15932
rect 20211 15929 20223 15963
rect 20165 15923 20223 15929
rect 22848 15904 22876 15991
rect 22925 15963 22983 15969
rect 22925 15929 22937 15963
rect 22971 15929 22983 15963
rect 23124 15960 23152 15991
rect 24578 15988 24584 16000
rect 24636 15988 24642 16040
rect 25225 16031 25283 16037
rect 25225 16028 25237 16031
rect 24872 16000 25237 16028
rect 24872 15972 24900 16000
rect 25225 15997 25237 16000
rect 25271 15997 25283 16031
rect 25225 15991 25283 15997
rect 25869 16031 25927 16037
rect 25869 15997 25881 16031
rect 25915 15997 25927 16031
rect 25869 15991 25927 15997
rect 23124 15932 23888 15960
rect 22925 15923 22983 15929
rect 11698 15892 11704 15904
rect 11440 15864 11704 15892
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 13078 15852 13084 15904
rect 13136 15852 13142 15904
rect 14918 15852 14924 15904
rect 14976 15892 14982 15904
rect 15289 15895 15347 15901
rect 15289 15892 15301 15895
rect 14976 15864 15301 15892
rect 14976 15852 14982 15864
rect 15289 15861 15301 15864
rect 15335 15861 15347 15895
rect 15289 15855 15347 15861
rect 17865 15895 17923 15901
rect 17865 15861 17877 15895
rect 17911 15892 17923 15895
rect 18874 15892 18880 15904
rect 17911 15864 18880 15892
rect 17911 15861 17923 15864
rect 17865 15855 17923 15861
rect 18874 15852 18880 15864
rect 18932 15852 18938 15904
rect 20073 15895 20131 15901
rect 20073 15861 20085 15895
rect 20119 15892 20131 15895
rect 20898 15892 20904 15904
rect 20119 15864 20904 15892
rect 20119 15861 20131 15864
rect 20073 15855 20131 15861
rect 20898 15852 20904 15864
rect 20956 15852 20962 15904
rect 22830 15852 22836 15904
rect 22888 15852 22894 15904
rect 22940 15892 22968 15923
rect 23290 15892 23296 15904
rect 22940 15864 23296 15892
rect 23290 15852 23296 15864
rect 23348 15852 23354 15904
rect 23860 15901 23888 15932
rect 24854 15920 24860 15972
rect 24912 15920 24918 15972
rect 24946 15920 24952 15972
rect 25004 15969 25010 15972
rect 25004 15960 25016 15969
rect 25004 15932 25049 15960
rect 25004 15923 25016 15932
rect 25004 15920 25010 15923
rect 23845 15895 23903 15901
rect 23845 15861 23857 15895
rect 23891 15892 23903 15895
rect 25884 15892 25912 15991
rect 26234 15988 26240 16040
rect 26292 15988 26298 16040
rect 23891 15864 25912 15892
rect 23891 15861 23903 15864
rect 23845 15855 23903 15861
rect 26602 15852 26608 15904
rect 26660 15892 26666 15904
rect 26789 15895 26847 15901
rect 26789 15892 26801 15895
rect 26660 15864 26801 15892
rect 26660 15852 26666 15864
rect 26789 15861 26801 15864
rect 26835 15861 26847 15895
rect 26789 15855 26847 15861
rect 552 15802 27576 15824
rect 552 15750 7114 15802
rect 7166 15750 7178 15802
rect 7230 15750 7242 15802
rect 7294 15750 7306 15802
rect 7358 15750 7370 15802
rect 7422 15750 13830 15802
rect 13882 15750 13894 15802
rect 13946 15750 13958 15802
rect 14010 15750 14022 15802
rect 14074 15750 14086 15802
rect 14138 15750 20546 15802
rect 20598 15750 20610 15802
rect 20662 15750 20674 15802
rect 20726 15750 20738 15802
rect 20790 15750 20802 15802
rect 20854 15750 27262 15802
rect 27314 15750 27326 15802
rect 27378 15750 27390 15802
rect 27442 15750 27454 15802
rect 27506 15750 27518 15802
rect 27570 15750 27576 15802
rect 552 15728 27576 15750
rect 8662 15688 8668 15700
rect 5368 15660 8668 15688
rect 4614 15512 4620 15564
rect 4672 15552 4678 15564
rect 5368 15561 5396 15660
rect 8662 15648 8668 15660
rect 8720 15648 8726 15700
rect 8754 15648 8760 15700
rect 8812 15648 8818 15700
rect 8846 15648 8852 15700
rect 8904 15688 8910 15700
rect 11606 15688 11612 15700
rect 8904 15660 11612 15688
rect 8904 15648 8910 15660
rect 11606 15648 11612 15660
rect 11664 15648 11670 15700
rect 12069 15691 12127 15697
rect 12069 15657 12081 15691
rect 12115 15688 12127 15691
rect 12434 15688 12440 15700
rect 12115 15660 12440 15688
rect 12115 15657 12127 15660
rect 12069 15651 12127 15657
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 18506 15648 18512 15700
rect 18564 15688 18570 15700
rect 18601 15691 18659 15697
rect 18601 15688 18613 15691
rect 18564 15660 18613 15688
rect 18564 15648 18570 15660
rect 18601 15657 18613 15660
rect 18647 15657 18659 15691
rect 18601 15651 18659 15657
rect 22094 15648 22100 15700
rect 22152 15648 22158 15700
rect 23290 15688 23296 15700
rect 22480 15660 23296 15688
rect 22480 15632 22508 15660
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 26878 15648 26884 15700
rect 26936 15688 26942 15700
rect 27065 15691 27123 15697
rect 27065 15688 27077 15691
rect 26936 15660 27077 15688
rect 26936 15648 26942 15660
rect 27065 15657 27077 15660
rect 27111 15657 27123 15691
rect 27065 15651 27123 15657
rect 7466 15620 7472 15632
rect 5552 15592 7472 15620
rect 5552 15561 5580 15592
rect 7466 15580 7472 15592
rect 7524 15580 7530 15632
rect 7650 15580 7656 15632
rect 7708 15620 7714 15632
rect 9674 15620 9680 15632
rect 7708 15592 9680 15620
rect 7708 15580 7714 15592
rect 5353 15555 5411 15561
rect 5353 15552 5365 15555
rect 4672 15524 5365 15552
rect 4672 15512 4678 15524
rect 5353 15521 5365 15524
rect 5399 15521 5411 15555
rect 5353 15515 5411 15521
rect 5537 15555 5595 15561
rect 5537 15521 5549 15555
rect 5583 15521 5595 15555
rect 5537 15515 5595 15521
rect 5810 15512 5816 15564
rect 5868 15512 5874 15564
rect 6080 15555 6138 15561
rect 6080 15521 6092 15555
rect 6126 15552 6138 15555
rect 6362 15552 6368 15564
rect 6126 15524 6368 15552
rect 6126 15521 6138 15524
rect 6080 15515 6138 15521
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 8202 15512 8208 15564
rect 8260 15552 8266 15564
rect 8772 15561 8800 15592
rect 9674 15580 9680 15592
rect 9732 15580 9738 15632
rect 10689 15623 10747 15629
rect 10689 15589 10701 15623
rect 10735 15620 10747 15623
rect 11057 15623 11115 15629
rect 11057 15620 11069 15623
rect 10735 15592 11069 15620
rect 10735 15589 10747 15592
rect 10689 15583 10747 15589
rect 11057 15589 11069 15592
rect 11103 15620 11115 15623
rect 12618 15620 12624 15632
rect 11103 15592 12624 15620
rect 11103 15589 11115 15592
rect 11057 15583 11115 15589
rect 8573 15555 8631 15561
rect 8573 15552 8585 15555
rect 8260 15524 8585 15552
rect 8260 15512 8266 15524
rect 8573 15521 8585 15524
rect 8619 15552 8631 15555
rect 8757 15555 8815 15561
rect 8619 15524 8708 15552
rect 8619 15521 8631 15524
rect 8573 15515 8631 15521
rect 5629 15487 5687 15493
rect 5629 15453 5641 15487
rect 5675 15453 5687 15487
rect 8680 15484 8708 15524
rect 8757 15521 8769 15555
rect 8803 15521 8815 15555
rect 10597 15555 10655 15561
rect 10597 15552 10609 15555
rect 8757 15515 8815 15521
rect 10060 15524 10609 15552
rect 9858 15484 9864 15496
rect 8680 15456 9864 15484
rect 5629 15447 5687 15453
rect 5166 15308 5172 15360
rect 5224 15308 5230 15360
rect 5644 15348 5672 15447
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 10060 15428 10088 15524
rect 10597 15521 10609 15524
rect 10643 15521 10655 15555
rect 10597 15515 10655 15521
rect 10962 15512 10968 15564
rect 11020 15512 11026 15564
rect 11241 15555 11299 15561
rect 11241 15521 11253 15555
rect 11287 15552 11299 15555
rect 11330 15552 11336 15564
rect 11287 15524 11336 15552
rect 11287 15521 11299 15524
rect 11241 15515 11299 15521
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 11716 15561 11744 15592
rect 12618 15580 12624 15592
rect 12676 15580 12682 15632
rect 12796 15623 12854 15629
rect 12796 15589 12808 15623
rect 12842 15620 12854 15623
rect 13078 15620 13084 15632
rect 12842 15592 13084 15620
rect 12842 15589 12854 15592
rect 12796 15583 12854 15589
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 18322 15620 18328 15632
rect 17236 15592 18328 15620
rect 11701 15555 11759 15561
rect 11701 15521 11713 15555
rect 11747 15521 11759 15555
rect 11701 15515 11759 15521
rect 11790 15512 11796 15564
rect 11848 15512 11854 15564
rect 12342 15512 12348 15564
rect 12400 15552 12406 15564
rect 12529 15555 12587 15561
rect 12529 15552 12541 15555
rect 12400 15524 12541 15552
rect 12400 15512 12406 15524
rect 12529 15521 12541 15524
rect 12575 15521 12587 15555
rect 12529 15515 12587 15521
rect 16666 15512 16672 15564
rect 16724 15552 16730 15564
rect 17236 15561 17264 15592
rect 18322 15580 18328 15592
rect 18380 15580 18386 15632
rect 19429 15623 19487 15629
rect 19429 15620 19441 15623
rect 18432 15592 19441 15620
rect 17221 15555 17279 15561
rect 17221 15552 17233 15555
rect 16724 15524 17233 15552
rect 16724 15512 16730 15524
rect 17221 15521 17233 15524
rect 17267 15521 17279 15555
rect 17221 15515 17279 15521
rect 17488 15555 17546 15561
rect 17488 15521 17500 15555
rect 17534 15552 17546 15555
rect 18432 15552 18460 15592
rect 19429 15589 19441 15592
rect 19475 15589 19487 15623
rect 19429 15583 19487 15589
rect 22462 15580 22468 15632
rect 22520 15580 22526 15632
rect 23474 15620 23480 15632
rect 22664 15592 23480 15620
rect 17534 15524 18460 15552
rect 18693 15555 18751 15561
rect 17534 15521 17546 15524
rect 17488 15515 17546 15521
rect 18693 15521 18705 15555
rect 18739 15521 18751 15555
rect 18693 15515 18751 15521
rect 18877 15555 18935 15561
rect 18877 15521 18889 15555
rect 18923 15521 18935 15555
rect 18877 15515 18935 15521
rect 18969 15555 19027 15561
rect 18969 15521 18981 15555
rect 19015 15521 19027 15555
rect 18969 15515 19027 15521
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15453 11667 15487
rect 11609 15447 11667 15453
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15484 14795 15487
rect 15470 15484 15476 15496
rect 14783 15456 15476 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 6914 15376 6920 15428
rect 6972 15416 6978 15428
rect 7193 15419 7251 15425
rect 7193 15416 7205 15419
rect 6972 15388 7205 15416
rect 6972 15376 6978 15388
rect 7193 15385 7205 15388
rect 7239 15416 7251 15419
rect 10042 15416 10048 15428
rect 7239 15388 10048 15416
rect 7239 15385 7251 15388
rect 7193 15379 7251 15385
rect 10042 15376 10048 15388
rect 10100 15376 10106 15428
rect 10962 15376 10968 15428
rect 11020 15416 11026 15428
rect 11624 15416 11652 15447
rect 11020 15388 11652 15416
rect 11020 15376 11026 15388
rect 11790 15376 11796 15428
rect 11848 15416 11854 15428
rect 11900 15416 11928 15447
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 11848 15388 11928 15416
rect 13909 15419 13967 15425
rect 11848 15376 11854 15388
rect 13909 15385 13921 15419
rect 13955 15416 13967 15419
rect 14274 15416 14280 15428
rect 13955 15388 14280 15416
rect 13955 15385 13967 15388
rect 13909 15379 13967 15385
rect 14274 15376 14280 15388
rect 14332 15376 14338 15428
rect 7006 15348 7012 15360
rect 5644 15320 7012 15348
rect 7006 15308 7012 15320
rect 7064 15308 7070 15360
rect 8662 15308 8668 15360
rect 8720 15348 8726 15360
rect 11146 15348 11152 15360
rect 8720 15320 11152 15348
rect 8720 15308 8726 15320
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 11422 15308 11428 15360
rect 11480 15308 11486 15360
rect 14093 15351 14151 15357
rect 14093 15317 14105 15351
rect 14139 15348 14151 15351
rect 14458 15348 14464 15360
rect 14139 15320 14464 15348
rect 14139 15317 14151 15320
rect 14093 15311 14151 15317
rect 14458 15308 14464 15320
rect 14516 15308 14522 15360
rect 18708 15348 18736 15515
rect 18892 15416 18920 15515
rect 18984 15484 19012 15515
rect 19058 15512 19064 15564
rect 19116 15512 19122 15564
rect 19610 15552 19616 15564
rect 19168 15524 19616 15552
rect 19168 15496 19196 15524
rect 19610 15512 19616 15524
rect 19668 15512 19674 15564
rect 21266 15512 21272 15564
rect 21324 15552 21330 15564
rect 22278 15561 22284 15564
rect 22235 15555 22284 15561
rect 22235 15552 22247 15555
rect 21324 15524 22247 15552
rect 21324 15512 21330 15524
rect 22235 15521 22247 15524
rect 22281 15521 22284 15555
rect 22235 15515 22284 15521
rect 22278 15512 22284 15515
rect 22336 15512 22342 15564
rect 22664 15561 22692 15592
rect 23474 15580 23480 15592
rect 23532 15580 23538 15632
rect 25124 15623 25182 15629
rect 25124 15589 25136 15623
rect 25170 15620 25182 15623
rect 25590 15620 25596 15632
rect 25170 15592 25596 15620
rect 25170 15589 25182 15592
rect 25124 15583 25182 15589
rect 25590 15580 25596 15592
rect 25648 15580 25654 15632
rect 22373 15555 22431 15561
rect 22373 15521 22385 15555
rect 22419 15521 22431 15555
rect 22373 15515 22431 15521
rect 22648 15555 22706 15561
rect 22648 15521 22660 15555
rect 22694 15521 22706 15555
rect 22648 15515 22706 15521
rect 19150 15484 19156 15496
rect 18984 15456 19156 15484
rect 19150 15444 19156 15456
rect 19208 15444 19214 15496
rect 19337 15487 19395 15493
rect 19337 15453 19349 15487
rect 19383 15484 19395 15487
rect 19981 15487 20039 15493
rect 19981 15484 19993 15487
rect 19383 15456 19993 15484
rect 19383 15453 19395 15456
rect 19337 15447 19395 15453
rect 19981 15453 19993 15456
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 20070 15444 20076 15496
rect 20128 15484 20134 15496
rect 20165 15487 20223 15493
rect 20165 15484 20177 15487
rect 20128 15456 20177 15484
rect 20128 15444 20134 15456
rect 20165 15453 20177 15456
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 21358 15444 21364 15496
rect 21416 15484 21422 15496
rect 22388 15484 22416 15515
rect 22738 15512 22744 15564
rect 22796 15512 22802 15564
rect 22833 15555 22891 15561
rect 22833 15521 22845 15555
rect 22879 15521 22891 15555
rect 22833 15515 22891 15521
rect 21416 15456 22416 15484
rect 21416 15444 21422 15456
rect 19886 15416 19892 15428
rect 18892 15388 19892 15416
rect 19886 15376 19892 15388
rect 19944 15376 19950 15428
rect 22848 15416 22876 15515
rect 23014 15512 23020 15564
rect 23072 15512 23078 15564
rect 23109 15555 23167 15561
rect 23109 15521 23121 15555
rect 23155 15521 23167 15555
rect 23109 15515 23167 15521
rect 23201 15555 23259 15561
rect 23201 15521 23213 15555
rect 23247 15552 23259 15555
rect 23569 15555 23627 15561
rect 23569 15552 23581 15555
rect 23247 15524 23581 15552
rect 23247 15521 23259 15524
rect 23201 15515 23259 15521
rect 23569 15521 23581 15524
rect 23615 15521 23627 15555
rect 23569 15515 23627 15521
rect 22922 15444 22928 15496
rect 22980 15484 22986 15496
rect 23124 15484 23152 15515
rect 26418 15512 26424 15564
rect 26476 15512 26482 15564
rect 26602 15561 26608 15564
rect 26569 15555 26608 15561
rect 26569 15521 26581 15555
rect 26569 15515 26608 15521
rect 26602 15512 26608 15515
rect 26660 15512 26666 15564
rect 26694 15512 26700 15564
rect 26752 15512 26758 15564
rect 26786 15512 26792 15564
rect 26844 15512 26850 15564
rect 26878 15512 26884 15564
rect 26936 15561 26942 15564
rect 26936 15552 26944 15561
rect 26936 15524 26981 15552
rect 26936 15515 26944 15524
rect 26936 15512 26942 15515
rect 22980 15456 23152 15484
rect 24213 15487 24271 15493
rect 22980 15444 22986 15456
rect 24213 15453 24225 15487
rect 24259 15484 24271 15487
rect 24762 15484 24768 15496
rect 24259 15456 24768 15484
rect 24259 15453 24271 15456
rect 24213 15447 24271 15453
rect 24762 15444 24768 15456
rect 24820 15444 24826 15496
rect 24854 15444 24860 15496
rect 24912 15444 24918 15496
rect 23566 15416 23572 15428
rect 22848 15388 23572 15416
rect 23566 15376 23572 15388
rect 23624 15376 23630 15428
rect 19242 15348 19248 15360
rect 18708 15320 19248 15348
rect 19242 15308 19248 15320
rect 19300 15308 19306 15360
rect 20714 15308 20720 15360
rect 20772 15348 20778 15360
rect 20809 15351 20867 15357
rect 20809 15348 20821 15351
rect 20772 15320 20821 15348
rect 20772 15308 20778 15320
rect 20809 15317 20821 15320
rect 20855 15317 20867 15351
rect 20809 15311 20867 15317
rect 22005 15351 22063 15357
rect 22005 15317 22017 15351
rect 22051 15348 22063 15351
rect 22094 15348 22100 15360
rect 22051 15320 22100 15348
rect 22051 15317 22063 15320
rect 22005 15311 22063 15317
rect 22094 15308 22100 15320
rect 22152 15308 22158 15360
rect 23474 15308 23480 15360
rect 23532 15308 23538 15360
rect 26237 15351 26295 15357
rect 26237 15317 26249 15351
rect 26283 15348 26295 15351
rect 26326 15348 26332 15360
rect 26283 15320 26332 15348
rect 26283 15317 26295 15320
rect 26237 15311 26295 15317
rect 26326 15308 26332 15320
rect 26384 15308 26390 15360
rect 552 15258 27416 15280
rect 552 15206 3756 15258
rect 3808 15206 3820 15258
rect 3872 15206 3884 15258
rect 3936 15206 3948 15258
rect 4000 15206 4012 15258
rect 4064 15206 10472 15258
rect 10524 15206 10536 15258
rect 10588 15206 10600 15258
rect 10652 15206 10664 15258
rect 10716 15206 10728 15258
rect 10780 15206 17188 15258
rect 17240 15206 17252 15258
rect 17304 15206 17316 15258
rect 17368 15206 17380 15258
rect 17432 15206 17444 15258
rect 17496 15206 23904 15258
rect 23956 15206 23968 15258
rect 24020 15206 24032 15258
rect 24084 15206 24096 15258
rect 24148 15206 24160 15258
rect 24212 15206 27416 15258
rect 552 15184 27416 15206
rect 6454 15104 6460 15156
rect 6512 15104 6518 15156
rect 7466 15104 7472 15156
rect 7524 15104 7530 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10413 15147 10471 15153
rect 10413 15144 10425 15147
rect 10008 15116 10425 15144
rect 10008 15104 10014 15116
rect 10413 15113 10425 15116
rect 10459 15113 10471 15147
rect 10873 15147 10931 15153
rect 10873 15144 10885 15147
rect 10413 15107 10471 15113
rect 10520 15116 10885 15144
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 3602 15008 3608 15020
rect 3007 14980 3608 15008
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 3602 14968 3608 14980
rect 3660 14968 3666 15020
rect 6472 15008 6500 15104
rect 9677 15079 9735 15085
rect 9677 15045 9689 15079
rect 9723 15076 9735 15079
rect 9861 15079 9919 15085
rect 9861 15076 9873 15079
rect 9723 15048 9873 15076
rect 9723 15045 9735 15048
rect 9677 15039 9735 15045
rect 9861 15045 9873 15048
rect 9907 15045 9919 15079
rect 9861 15039 9919 15045
rect 10226 15036 10232 15088
rect 10284 15076 10290 15088
rect 10520 15076 10548 15116
rect 10873 15113 10885 15116
rect 10919 15113 10931 15147
rect 10873 15107 10931 15113
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11241 15147 11299 15153
rect 11241 15144 11253 15147
rect 11112 15116 11253 15144
rect 11112 15104 11118 15116
rect 11241 15113 11253 15116
rect 11287 15113 11299 15147
rect 11241 15107 11299 15113
rect 11330 15104 11336 15156
rect 11388 15144 11394 15156
rect 13354 15144 13360 15156
rect 11388 15116 13360 15144
rect 11388 15104 11394 15116
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 15470 15104 15476 15156
rect 15528 15104 15534 15156
rect 17034 15104 17040 15156
rect 17092 15104 17098 15156
rect 19058 15144 19064 15156
rect 17972 15116 19064 15144
rect 10284 15048 10548 15076
rect 10597 15079 10655 15085
rect 10284 15036 10290 15048
rect 10597 15045 10609 15079
rect 10643 15076 10655 15079
rect 10962 15076 10968 15088
rect 10643 15048 10968 15076
rect 10643 15045 10655 15048
rect 10597 15039 10655 15045
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 11146 15036 11152 15088
rect 11204 15076 11210 15088
rect 11348 15076 11376 15104
rect 11204 15048 11376 15076
rect 11204 15036 11210 15048
rect 7101 15011 7159 15017
rect 7101 15008 7113 15011
rect 6472 14980 7113 15008
rect 7101 14977 7113 14980
rect 7147 15008 7159 15011
rect 7653 15011 7711 15017
rect 7147 14980 7604 15008
rect 7147 14977 7159 14980
rect 7101 14971 7159 14977
rect 2777 14943 2835 14949
rect 2777 14909 2789 14943
rect 2823 14909 2835 14943
rect 2777 14903 2835 14909
rect 3053 14943 3111 14949
rect 3053 14909 3065 14943
rect 3099 14940 3111 14943
rect 3786 14940 3792 14952
rect 3099 14912 3792 14940
rect 3099 14909 3111 14912
rect 3053 14903 3111 14909
rect 2038 14832 2044 14884
rect 2096 14872 2102 14884
rect 2792 14872 2820 14903
rect 3786 14900 3792 14912
rect 3844 14900 3850 14952
rect 3881 14943 3939 14949
rect 3881 14909 3893 14943
rect 3927 14940 3939 14943
rect 4154 14940 4160 14952
rect 3927 14912 4160 14940
rect 3927 14909 3939 14912
rect 3881 14903 3939 14909
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14940 5135 14943
rect 5810 14940 5816 14952
rect 5123 14912 5816 14940
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 5810 14900 5816 14912
rect 5868 14940 5874 14952
rect 6822 14940 6828 14952
rect 5868 14912 6828 14940
rect 5868 14900 5874 14912
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 7006 14900 7012 14952
rect 7064 14940 7070 14952
rect 7469 14943 7527 14949
rect 7469 14940 7481 14943
rect 7064 14912 7481 14940
rect 7064 14900 7070 14912
rect 7469 14909 7481 14912
rect 7515 14909 7527 14943
rect 7576 14940 7604 14980
rect 7653 14977 7665 15011
rect 7699 15008 7711 15011
rect 8113 15011 8171 15017
rect 8113 15008 8125 15011
rect 7699 14980 8125 15008
rect 7699 14977 7711 14980
rect 7653 14971 7711 14977
rect 8113 14977 8125 14980
rect 8159 14977 8171 15011
rect 11422 15008 11428 15020
rect 8113 14971 8171 14977
rect 9508 14980 11428 15008
rect 8021 14943 8079 14949
rect 8021 14940 8033 14943
rect 7576 14912 8033 14940
rect 7469 14903 7527 14909
rect 8021 14909 8033 14912
rect 8067 14909 8079 14943
rect 8021 14903 8079 14909
rect 8205 14943 8263 14949
rect 8205 14909 8217 14943
rect 8251 14940 8263 14943
rect 8478 14940 8484 14952
rect 8251 14912 8484 14940
rect 8251 14909 8263 14912
rect 8205 14903 8263 14909
rect 8478 14900 8484 14912
rect 8536 14900 8542 14952
rect 9508 14949 9536 14980
rect 11422 14968 11428 14980
rect 11480 15008 11486 15020
rect 11480 14980 11652 15008
rect 11480 14968 11486 14980
rect 9493 14943 9551 14949
rect 9493 14909 9505 14943
rect 9539 14909 9551 14943
rect 9493 14903 9551 14909
rect 9674 14900 9680 14952
rect 9732 14940 9738 14952
rect 9769 14943 9827 14949
rect 9769 14940 9781 14943
rect 9732 14912 9781 14940
rect 9732 14900 9738 14912
rect 9769 14909 9781 14912
rect 9815 14940 9827 14943
rect 9815 14912 9996 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 3237 14875 3295 14881
rect 3237 14872 3249 14875
rect 2096 14844 2728 14872
rect 2792 14844 3249 14872
rect 2096 14832 2102 14844
rect 2314 14764 2320 14816
rect 2372 14804 2378 14816
rect 2593 14807 2651 14813
rect 2593 14804 2605 14807
rect 2372 14776 2605 14804
rect 2372 14764 2378 14776
rect 2593 14773 2605 14776
rect 2639 14773 2651 14807
rect 2700 14804 2728 14844
rect 3237 14841 3249 14844
rect 3283 14841 3295 14875
rect 3237 14835 3295 14841
rect 5166 14832 5172 14884
rect 5224 14872 5230 14884
rect 5322 14875 5380 14881
rect 5322 14872 5334 14875
rect 5224 14844 5334 14872
rect 5224 14832 5230 14844
rect 5322 14841 5334 14844
rect 5368 14841 5380 14875
rect 7650 14872 7656 14884
rect 5322 14835 5380 14841
rect 5828 14844 7656 14872
rect 5828 14804 5856 14844
rect 7650 14832 7656 14844
rect 7708 14832 7714 14884
rect 7929 14875 7987 14881
rect 7929 14841 7941 14875
rect 7975 14872 7987 14875
rect 7975 14844 9076 14872
rect 7975 14841 7987 14844
rect 7929 14835 7987 14841
rect 9048 14816 9076 14844
rect 9858 14832 9864 14884
rect 9916 14832 9922 14884
rect 9968 14872 9996 14912
rect 10042 14900 10048 14952
rect 10100 14900 10106 14952
rect 10137 14943 10195 14949
rect 10137 14909 10149 14943
rect 10183 14940 10195 14943
rect 11146 14940 11152 14952
rect 10183 14912 11152 14940
rect 10183 14909 10195 14912
rect 10137 14903 10195 14909
rect 11146 14900 11152 14912
rect 11204 14900 11210 14952
rect 11624 14949 11652 14980
rect 11698 14968 11704 15020
rect 11756 15008 11762 15020
rect 11756 14980 11836 15008
rect 11756 14968 11762 14980
rect 11808 14949 11836 14980
rect 11333 14943 11391 14949
rect 11333 14909 11345 14943
rect 11379 14909 11391 14943
rect 11333 14903 11391 14909
rect 11609 14943 11667 14949
rect 11609 14909 11621 14943
rect 11655 14909 11667 14943
rect 11609 14903 11667 14909
rect 11793 14943 11851 14949
rect 11793 14909 11805 14943
rect 11839 14909 11851 14943
rect 11793 14903 11851 14909
rect 10229 14875 10287 14881
rect 10229 14872 10241 14875
rect 9968 14844 10241 14872
rect 10229 14841 10241 14844
rect 10275 14841 10287 14875
rect 11057 14875 11115 14881
rect 11057 14872 11069 14875
rect 10229 14835 10287 14841
rect 10336 14844 11069 14872
rect 10336 14816 10364 14844
rect 11057 14841 11069 14844
rect 11103 14841 11115 14875
rect 11057 14835 11115 14841
rect 11348 14816 11376 14903
rect 11974 14900 11980 14952
rect 12032 14940 12038 14952
rect 14093 14943 14151 14949
rect 12032 14912 12388 14940
rect 12032 14900 12038 14912
rect 12360 14884 12388 14912
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 14182 14940 14188 14952
rect 14139 14912 14188 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 14182 14900 14188 14912
rect 14240 14940 14246 14952
rect 15657 14943 15715 14949
rect 15657 14940 15669 14943
rect 14240 14912 15669 14940
rect 14240 14900 14246 14912
rect 15657 14909 15669 14912
rect 15703 14940 15715 14943
rect 16666 14940 16672 14952
rect 15703 14912 16672 14940
rect 15703 14909 15715 14912
rect 15657 14903 15715 14909
rect 16666 14900 16672 14912
rect 16724 14900 16730 14952
rect 16942 14900 16948 14952
rect 17000 14940 17006 14952
rect 17589 14943 17647 14949
rect 17589 14940 17601 14943
rect 17000 14912 17601 14940
rect 17000 14900 17006 14912
rect 17589 14909 17601 14912
rect 17635 14909 17647 14943
rect 17589 14903 17647 14909
rect 17737 14943 17795 14949
rect 17737 14909 17749 14943
rect 17783 14940 17795 14943
rect 17972 14940 18000 15116
rect 19058 15104 19064 15116
rect 19116 15104 19122 15156
rect 19886 15104 19892 15156
rect 19944 15144 19950 15156
rect 20165 15147 20223 15153
rect 20165 15144 20177 15147
rect 19944 15116 20177 15144
rect 19944 15104 19950 15116
rect 20165 15113 20177 15116
rect 20211 15113 20223 15147
rect 22738 15144 22744 15156
rect 20165 15107 20223 15113
rect 21008 15116 22744 15144
rect 18233 15079 18291 15085
rect 18233 15045 18245 15079
rect 18279 15076 18291 15079
rect 18279 15048 19196 15076
rect 18279 15045 18291 15048
rect 18233 15039 18291 15045
rect 17783 14912 18000 14940
rect 18095 14943 18153 14949
rect 17783 14909 17795 14912
rect 17737 14903 17795 14909
rect 18095 14909 18107 14943
rect 18141 14940 18153 14943
rect 18598 14940 18604 14952
rect 18141 14912 18604 14940
rect 18141 14909 18153 14912
rect 18095 14903 18153 14909
rect 18598 14900 18604 14912
rect 18656 14900 18662 14952
rect 18874 14900 18880 14952
rect 18932 14940 18938 14952
rect 18969 14943 19027 14949
rect 18969 14940 18981 14943
rect 18932 14912 18981 14940
rect 18932 14900 18938 14912
rect 18969 14909 18981 14912
rect 19015 14909 19027 14943
rect 18969 14903 19027 14909
rect 19058 14900 19064 14952
rect 19116 14900 19122 14952
rect 19168 14949 19196 15048
rect 19794 14968 19800 15020
rect 19852 15008 19858 15020
rect 20254 15008 20260 15020
rect 19852 14980 20260 15008
rect 19852 14968 19858 14980
rect 20254 14968 20260 14980
rect 20312 14968 20318 15020
rect 20898 15008 20904 15020
rect 20732 14980 20904 15008
rect 19153 14943 19211 14949
rect 19153 14909 19165 14943
rect 19199 14909 19211 14943
rect 19153 14903 19211 14909
rect 19242 14900 19248 14952
rect 19300 14940 19306 14952
rect 19337 14943 19395 14949
rect 19337 14940 19349 14943
rect 19300 14912 19349 14940
rect 19300 14900 19306 14912
rect 19337 14909 19349 14912
rect 19383 14909 19395 14943
rect 19337 14903 19395 14909
rect 20073 14943 20131 14949
rect 20073 14909 20085 14943
rect 20119 14940 20131 14943
rect 20162 14940 20168 14952
rect 20119 14912 20168 14940
rect 20119 14909 20131 14912
rect 20073 14903 20131 14909
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 20346 14949 20352 14952
rect 20344 14940 20352 14949
rect 20307 14912 20352 14940
rect 20344 14903 20352 14912
rect 20346 14900 20352 14903
rect 20404 14900 20410 14952
rect 20441 14943 20499 14949
rect 20441 14909 20453 14943
rect 20487 14940 20499 14943
rect 20622 14940 20628 14952
rect 20487 14912 20628 14940
rect 20487 14909 20499 14912
rect 20441 14903 20499 14909
rect 20622 14900 20628 14912
rect 20680 14900 20686 14952
rect 20732 14949 20760 14980
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 21008 14952 21036 15116
rect 22738 15104 22744 15116
rect 22796 15104 22802 15156
rect 24486 15104 24492 15156
rect 24544 15144 24550 15156
rect 24762 15144 24768 15156
rect 24544 15116 24768 15144
rect 24544 15104 24550 15116
rect 24762 15104 24768 15116
rect 24820 15144 24826 15156
rect 25225 15147 25283 15153
rect 25225 15144 25237 15147
rect 24820 15116 25237 15144
rect 24820 15104 24826 15116
rect 25225 15113 25237 15116
rect 25271 15113 25283 15147
rect 25225 15107 25283 15113
rect 21082 14968 21088 15020
rect 21140 15008 21146 15020
rect 21177 15011 21235 15017
rect 21177 15008 21189 15011
rect 21140 14980 21189 15008
rect 21140 14968 21146 14980
rect 21177 14977 21189 14980
rect 21223 14977 21235 15011
rect 23842 15008 23848 15020
rect 21177 14971 21235 14977
rect 23124 14980 23848 15008
rect 20716 14943 20774 14949
rect 20716 14909 20728 14943
rect 20762 14909 20774 14943
rect 20716 14903 20774 14909
rect 20809 14943 20867 14949
rect 20809 14909 20821 14943
rect 20855 14940 20867 14943
rect 20990 14940 20996 14952
rect 20855 14912 20996 14940
rect 20855 14909 20867 14912
rect 20809 14903 20867 14909
rect 20990 14900 20996 14912
rect 21048 14900 21054 14952
rect 21192 14940 21220 14971
rect 21726 14940 21732 14952
rect 21192 14912 21732 14940
rect 21726 14900 21732 14912
rect 21784 14940 21790 14952
rect 22738 14940 22744 14952
rect 21784 14912 22744 14940
rect 21784 14900 21790 14912
rect 22738 14900 22744 14912
rect 22796 14940 22802 14952
rect 23124 14940 23152 14980
rect 23842 14968 23848 14980
rect 23900 14968 23906 15020
rect 26329 15011 26387 15017
rect 26329 14977 26341 15011
rect 26375 15008 26387 15011
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26375 14980 26985 15008
rect 26375 14977 26387 14980
rect 26329 14971 26387 14977
rect 26973 14977 26985 14980
rect 27019 14977 27031 15011
rect 26973 14971 27031 14977
rect 22796 14912 23152 14940
rect 22796 14900 22802 14912
rect 23198 14900 23204 14952
rect 23256 14900 23262 14952
rect 25685 14943 25743 14949
rect 25685 14940 25697 14943
rect 24964 14912 25697 14940
rect 11701 14875 11759 14881
rect 11701 14841 11713 14875
rect 11747 14872 11759 14875
rect 12222 14875 12280 14881
rect 12222 14872 12234 14875
rect 11747 14844 12234 14872
rect 11747 14841 11759 14844
rect 11701 14835 11759 14841
rect 12222 14841 12234 14844
rect 12268 14841 12280 14875
rect 12222 14835 12280 14841
rect 12342 14832 12348 14884
rect 12400 14832 12406 14884
rect 14366 14881 14372 14884
rect 14360 14835 14372 14881
rect 14366 14832 14372 14835
rect 14424 14832 14430 14884
rect 15924 14875 15982 14881
rect 15924 14841 15936 14875
rect 15970 14872 15982 14875
rect 15970 14844 17356 14872
rect 15970 14841 15982 14844
rect 15924 14835 15982 14841
rect 2700 14776 5856 14804
rect 2593 14767 2651 14773
rect 6546 14764 6552 14816
rect 6604 14764 6610 14816
rect 6638 14764 6644 14816
rect 6696 14804 6702 14816
rect 7285 14807 7343 14813
rect 7285 14804 7297 14807
rect 6696 14776 7297 14804
rect 6696 14764 6702 14776
rect 7285 14773 7297 14776
rect 7331 14773 7343 14807
rect 7285 14767 7343 14773
rect 9030 14764 9036 14816
rect 9088 14804 9094 14816
rect 9309 14807 9367 14813
rect 9309 14804 9321 14807
rect 9088 14776 9321 14804
rect 9088 14764 9094 14776
rect 9309 14773 9321 14776
rect 9355 14773 9367 14807
rect 9309 14767 9367 14773
rect 10042 14764 10048 14816
rect 10100 14804 10106 14816
rect 10318 14804 10324 14816
rect 10100 14776 10324 14804
rect 10100 14764 10106 14776
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 10439 14807 10497 14813
rect 10439 14773 10451 14807
rect 10485 14804 10497 14807
rect 10594 14804 10600 14816
rect 10485 14776 10600 14804
rect 10485 14773 10497 14776
rect 10439 14767 10497 14773
rect 10594 14764 10600 14776
rect 10652 14804 10658 14816
rect 10689 14807 10747 14813
rect 10689 14804 10701 14807
rect 10652 14776 10701 14804
rect 10652 14764 10658 14776
rect 10689 14773 10701 14776
rect 10735 14773 10747 14807
rect 10689 14767 10747 14773
rect 10857 14807 10915 14813
rect 10857 14773 10869 14807
rect 10903 14804 10915 14807
rect 11146 14804 11152 14816
rect 10903 14776 11152 14804
rect 10903 14773 10915 14776
rect 10857 14767 10915 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 13357 14807 13415 14813
rect 13357 14804 13369 14807
rect 11388 14776 13369 14804
rect 11388 14764 11394 14776
rect 13357 14773 13369 14776
rect 13403 14804 13415 14807
rect 13538 14804 13544 14816
rect 13403 14776 13544 14804
rect 13403 14773 13415 14776
rect 13357 14767 13415 14773
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 13722 14764 13728 14816
rect 13780 14804 13786 14816
rect 16114 14804 16120 14816
rect 13780 14776 16120 14804
rect 13780 14764 13786 14776
rect 16114 14764 16120 14776
rect 16172 14764 16178 14816
rect 17328 14804 17356 14844
rect 17862 14832 17868 14884
rect 17920 14832 17926 14884
rect 17957 14875 18015 14881
rect 17957 14841 17969 14875
rect 18003 14872 18015 14875
rect 18230 14872 18236 14884
rect 18003 14844 18236 14872
rect 18003 14841 18015 14844
rect 17957 14835 18015 14841
rect 18230 14832 18236 14844
rect 18288 14832 18294 14884
rect 18782 14832 18788 14884
rect 18840 14872 18846 14884
rect 20533 14875 20591 14881
rect 20533 14872 20545 14875
rect 18840 14844 20545 14872
rect 18840 14832 18846 14844
rect 20533 14841 20545 14844
rect 20579 14841 20591 14875
rect 20533 14835 20591 14841
rect 21444 14875 21502 14881
rect 21444 14841 21456 14875
rect 21490 14872 21502 14875
rect 22278 14872 22284 14884
rect 21490 14844 22284 14872
rect 21490 14841 21502 14844
rect 21444 14835 21502 14841
rect 18693 14807 18751 14813
rect 18693 14804 18705 14807
rect 17328 14776 18705 14804
rect 18693 14773 18705 14776
rect 18739 14773 18751 14807
rect 18693 14767 18751 14773
rect 19426 14764 19432 14816
rect 19484 14764 19490 14816
rect 20548 14804 20576 14835
rect 22278 14832 22284 14844
rect 22336 14832 22342 14884
rect 22370 14832 22376 14884
rect 22428 14872 22434 14884
rect 22649 14875 22707 14881
rect 22649 14872 22661 14875
rect 22428 14844 22661 14872
rect 22428 14832 22434 14844
rect 22649 14841 22661 14844
rect 22695 14841 22707 14875
rect 22649 14835 22707 14841
rect 23474 14832 23480 14884
rect 23532 14872 23538 14884
rect 24090 14875 24148 14881
rect 24090 14872 24102 14875
rect 23532 14844 24102 14872
rect 23532 14832 23538 14844
rect 24090 14841 24102 14844
rect 24136 14841 24148 14875
rect 24090 14835 24148 14841
rect 24670 14832 24676 14884
rect 24728 14872 24734 14884
rect 24964 14872 24992 14912
rect 25685 14909 25697 14912
rect 25731 14909 25743 14943
rect 25685 14903 25743 14909
rect 25866 14900 25872 14952
rect 25924 14900 25930 14952
rect 25958 14900 25964 14952
rect 26016 14900 26022 14952
rect 26053 14943 26111 14949
rect 26053 14909 26065 14943
rect 26099 14940 26111 14943
rect 26602 14940 26608 14952
rect 26099 14912 26608 14940
rect 26099 14909 26111 14912
rect 26053 14903 26111 14909
rect 26602 14900 26608 14912
rect 26660 14900 26666 14952
rect 24728 14844 24992 14872
rect 24728 14832 24734 14844
rect 25038 14832 25044 14884
rect 25096 14872 25102 14884
rect 25976 14872 26004 14900
rect 25096 14844 26004 14872
rect 25096 14832 25102 14844
rect 21174 14804 21180 14816
rect 20548 14776 21180 14804
rect 21174 14764 21180 14776
rect 21232 14804 21238 14816
rect 22462 14804 22468 14816
rect 21232 14776 22468 14804
rect 21232 14764 21238 14776
rect 22462 14764 22468 14776
rect 22520 14764 22526 14816
rect 22557 14807 22615 14813
rect 22557 14773 22569 14807
rect 22603 14804 22615 14807
rect 22830 14804 22836 14816
rect 22603 14776 22836 14804
rect 22603 14773 22615 14776
rect 22557 14767 22615 14773
rect 22830 14764 22836 14776
rect 22888 14764 22894 14816
rect 23290 14764 23296 14816
rect 23348 14804 23354 14816
rect 24394 14804 24400 14816
rect 23348 14776 24400 14804
rect 23348 14764 23354 14776
rect 24394 14764 24400 14776
rect 24452 14764 24458 14816
rect 26418 14764 26424 14816
rect 26476 14764 26482 14816
rect 552 14714 27576 14736
rect 552 14662 7114 14714
rect 7166 14662 7178 14714
rect 7230 14662 7242 14714
rect 7294 14662 7306 14714
rect 7358 14662 7370 14714
rect 7422 14662 13830 14714
rect 13882 14662 13894 14714
rect 13946 14662 13958 14714
rect 14010 14662 14022 14714
rect 14074 14662 14086 14714
rect 14138 14662 20546 14714
rect 20598 14662 20610 14714
rect 20662 14662 20674 14714
rect 20726 14662 20738 14714
rect 20790 14662 20802 14714
rect 20854 14662 27262 14714
rect 27314 14662 27326 14714
rect 27378 14662 27390 14714
rect 27442 14662 27454 14714
rect 27506 14662 27518 14714
rect 27570 14662 27576 14714
rect 552 14640 27576 14662
rect 3786 14560 3792 14612
rect 3844 14560 3850 14612
rect 6362 14560 6368 14612
rect 6420 14560 6426 14612
rect 6454 14560 6460 14612
rect 6512 14600 6518 14612
rect 10594 14600 10600 14612
rect 6512 14572 6776 14600
rect 6512 14560 6518 14572
rect 2041 14467 2099 14473
rect 2041 14433 2053 14467
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 2056 14328 2084 14427
rect 2314 14424 2320 14476
rect 2372 14424 2378 14476
rect 2676 14467 2734 14473
rect 2676 14433 2688 14467
rect 2722 14464 2734 14467
rect 3234 14464 3240 14476
rect 2722 14436 3240 14464
rect 2722 14433 2734 14436
rect 2676 14427 2734 14433
rect 3234 14424 3240 14436
rect 3292 14424 3298 14476
rect 3804 14464 3832 14560
rect 5997 14535 6055 14541
rect 5997 14501 6009 14535
rect 6043 14532 6055 14535
rect 6638 14532 6644 14544
rect 6043 14504 6644 14532
rect 6043 14501 6055 14504
rect 5997 14495 6055 14501
rect 6638 14492 6644 14504
rect 6696 14492 6702 14544
rect 4246 14464 4252 14476
rect 3804 14436 4252 14464
rect 4246 14424 4252 14436
rect 4304 14464 4310 14476
rect 4433 14467 4491 14473
rect 4433 14464 4445 14467
rect 4304 14436 4445 14464
rect 4304 14424 4310 14436
rect 4433 14433 4445 14436
rect 4479 14464 4491 14467
rect 5169 14467 5227 14473
rect 5169 14464 5181 14467
rect 4479 14436 5181 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 5169 14433 5181 14436
rect 5215 14433 5227 14467
rect 5169 14427 5227 14433
rect 6546 14424 6552 14476
rect 6604 14424 6610 14476
rect 6748 14473 6776 14572
rect 6840 14572 10600 14600
rect 6840 14473 6868 14572
rect 10594 14560 10600 14572
rect 10652 14560 10658 14612
rect 10689 14603 10747 14609
rect 10689 14569 10701 14603
rect 10735 14600 10747 14603
rect 10870 14600 10876 14612
rect 10735 14572 10876 14600
rect 10735 14569 10747 14572
rect 10689 14563 10747 14569
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 11517 14603 11575 14609
rect 11517 14569 11529 14603
rect 11563 14600 11575 14603
rect 11606 14600 11612 14612
rect 11563 14572 11612 14600
rect 11563 14569 11575 14572
rect 11517 14563 11575 14569
rect 11606 14560 11612 14572
rect 11664 14560 11670 14612
rect 13817 14603 13875 14609
rect 13817 14569 13829 14603
rect 13863 14600 13875 14603
rect 14366 14600 14372 14612
rect 13863 14572 14372 14600
rect 13863 14569 13875 14572
rect 13817 14563 13875 14569
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 14458 14560 14464 14612
rect 14516 14560 14522 14612
rect 16390 14600 16396 14612
rect 14660 14572 16396 14600
rect 7453 14535 7511 14541
rect 7453 14501 7465 14535
rect 7499 14532 7511 14535
rect 7653 14535 7711 14541
rect 7499 14504 7604 14532
rect 7499 14501 7511 14504
rect 7453 14495 7511 14501
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 6825 14467 6883 14473
rect 6825 14433 6837 14467
rect 6871 14433 6883 14467
rect 6825 14427 6883 14433
rect 7576 14464 7604 14504
rect 7653 14501 7665 14535
rect 7699 14532 7711 14535
rect 8294 14532 8300 14544
rect 7699 14504 8300 14532
rect 7699 14501 7711 14504
rect 7653 14495 7711 14501
rect 8294 14492 8300 14504
rect 8352 14492 8358 14544
rect 9582 14532 9588 14544
rect 8404 14504 9076 14532
rect 7742 14464 7748 14476
rect 7576 14436 7748 14464
rect 2406 14356 2412 14408
rect 2464 14356 2470 14408
rect 3418 14356 3424 14408
rect 3476 14396 3482 14408
rect 4614 14396 4620 14408
rect 3476 14368 4620 14396
rect 3476 14356 3482 14368
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 4893 14399 4951 14405
rect 4893 14396 4905 14399
rect 4856 14368 4905 14396
rect 4856 14356 4862 14368
rect 4893 14365 4905 14368
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 6638 14356 6644 14408
rect 6696 14356 6702 14408
rect 7576 14396 7604 14436
rect 7742 14424 7748 14436
rect 7800 14424 7806 14476
rect 8404 14473 8432 14504
rect 9048 14476 9076 14504
rect 9508 14504 9588 14532
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14433 8447 14467
rect 8389 14427 8447 14433
rect 8478 14424 8484 14476
rect 8536 14464 8542 14476
rect 8757 14467 8815 14473
rect 8757 14464 8769 14467
rect 8536 14436 8769 14464
rect 8536 14424 8542 14436
rect 6840 14368 7604 14396
rect 2056 14300 2360 14328
rect 1762 14220 1768 14272
rect 1820 14260 1826 14272
rect 1857 14263 1915 14269
rect 1857 14260 1869 14263
rect 1820 14232 1869 14260
rect 1820 14220 1826 14232
rect 1857 14229 1869 14232
rect 1903 14229 1915 14263
rect 1857 14223 1915 14229
rect 2222 14220 2228 14272
rect 2280 14220 2286 14272
rect 2332 14260 2360 14300
rect 3510 14288 3516 14340
rect 3568 14328 3574 14340
rect 3881 14331 3939 14337
rect 3881 14328 3893 14331
rect 3568 14300 3893 14328
rect 3568 14288 3574 14300
rect 3881 14297 3893 14300
rect 3927 14297 3939 14331
rect 5813 14331 5871 14337
rect 5813 14328 5825 14331
rect 3881 14291 3939 14297
rect 4540 14300 5825 14328
rect 2682 14260 2688 14272
rect 2332 14232 2688 14260
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 3602 14220 3608 14272
rect 3660 14260 3666 14272
rect 4540 14260 4568 14300
rect 3660 14232 4568 14260
rect 3660 14220 3666 14232
rect 4614 14220 4620 14272
rect 4672 14220 4678 14272
rect 4816 14269 4844 14300
rect 5813 14297 5825 14300
rect 5859 14297 5871 14331
rect 5813 14291 5871 14297
rect 5902 14288 5908 14340
rect 5960 14328 5966 14340
rect 6840 14328 6868 14368
rect 5960 14300 6868 14328
rect 5960 14288 5966 14300
rect 7006 14288 7012 14340
rect 7064 14328 7070 14340
rect 7285 14331 7343 14337
rect 7285 14328 7297 14331
rect 7064 14300 7297 14328
rect 7064 14288 7070 14300
rect 7285 14297 7297 14300
rect 7331 14297 7343 14331
rect 8588 14328 8616 14436
rect 8757 14433 8769 14436
rect 8803 14433 8815 14467
rect 8757 14427 8815 14433
rect 9030 14424 9036 14476
rect 9088 14424 9094 14476
rect 9508 14473 9536 14504
rect 9582 14492 9588 14504
rect 9640 14532 9646 14544
rect 9858 14532 9864 14544
rect 9640 14504 9864 14532
rect 9640 14492 9646 14504
rect 9858 14492 9864 14504
rect 9916 14492 9922 14544
rect 11977 14535 12035 14541
rect 9968 14504 10272 14532
rect 9493 14467 9551 14473
rect 9493 14433 9505 14467
rect 9539 14433 9551 14467
rect 9968 14464 9996 14504
rect 9493 14427 9551 14433
rect 9600 14436 9996 14464
rect 8665 14399 8723 14405
rect 8665 14365 8677 14399
rect 8711 14396 8723 14399
rect 9217 14399 9275 14405
rect 9217 14396 9229 14399
rect 8711 14368 9229 14396
rect 8711 14365 8723 14368
rect 8665 14359 8723 14365
rect 9217 14365 9229 14368
rect 9263 14365 9275 14399
rect 9217 14359 9275 14365
rect 9398 14356 9404 14408
rect 9456 14396 9462 14408
rect 9600 14396 9628 14436
rect 10134 14422 10140 14474
rect 10192 14422 10198 14474
rect 10244 14462 10272 14504
rect 11977 14501 11989 14535
rect 12023 14532 12035 14535
rect 14476 14532 14504 14560
rect 12023 14504 14504 14532
rect 12023 14501 12035 14504
rect 11977 14495 12035 14501
rect 10321 14462 10379 14463
rect 10244 14457 10379 14462
rect 10244 14434 10333 14457
rect 10321 14423 10333 14434
rect 10367 14423 10379 14457
rect 10410 14424 10416 14476
rect 10468 14464 10474 14476
rect 10597 14467 10655 14473
rect 10597 14464 10609 14467
rect 10468 14436 10609 14464
rect 10468 14424 10474 14436
rect 10597 14433 10609 14436
rect 10643 14433 10655 14467
rect 10597 14427 10655 14433
rect 10781 14467 10839 14473
rect 10781 14433 10793 14467
rect 10827 14464 10839 14467
rect 10870 14464 10876 14476
rect 10827 14436 10876 14464
rect 10827 14433 10839 14436
rect 10781 14427 10839 14433
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 11146 14424 11152 14476
rect 11204 14424 11210 14476
rect 11330 14424 11336 14476
rect 11388 14424 11394 14476
rect 11885 14467 11943 14473
rect 11885 14433 11897 14467
rect 11931 14464 11943 14467
rect 13078 14464 13084 14476
rect 11931 14436 13084 14464
rect 11931 14433 11943 14436
rect 11885 14427 11943 14433
rect 13078 14424 13084 14436
rect 13136 14424 13142 14476
rect 13354 14424 13360 14476
rect 13412 14424 13418 14476
rect 13538 14424 13544 14476
rect 13596 14424 13602 14476
rect 14108 14473 14136 14504
rect 14093 14467 14151 14473
rect 14093 14433 14105 14467
rect 14139 14433 14151 14467
rect 14093 14427 14151 14433
rect 14185 14467 14243 14473
rect 14185 14433 14197 14467
rect 14231 14433 14243 14467
rect 14185 14427 14243 14433
rect 14277 14467 14335 14473
rect 14277 14433 14289 14467
rect 14323 14433 14335 14467
rect 14277 14427 14335 14433
rect 14461 14467 14519 14473
rect 14461 14433 14473 14467
rect 14507 14464 14519 14467
rect 14553 14467 14611 14473
rect 14553 14464 14565 14467
rect 14507 14436 14565 14464
rect 14507 14433 14519 14436
rect 14461 14427 14519 14433
rect 14553 14433 14565 14436
rect 14599 14433 14611 14467
rect 14660 14462 14688 14572
rect 16390 14560 16396 14572
rect 16448 14560 16454 14612
rect 17037 14603 17095 14609
rect 17037 14569 17049 14603
rect 17083 14569 17095 14603
rect 17037 14563 17095 14569
rect 17052 14532 17080 14563
rect 17862 14560 17868 14612
rect 17920 14600 17926 14612
rect 18138 14600 18144 14612
rect 17920 14572 18144 14600
rect 17920 14560 17926 14572
rect 18138 14560 18144 14572
rect 18196 14600 18202 14612
rect 18782 14600 18788 14612
rect 18196 14572 18788 14600
rect 18196 14560 18202 14572
rect 18782 14560 18788 14572
rect 18840 14560 18846 14612
rect 19705 14603 19763 14609
rect 19705 14569 19717 14603
rect 19751 14600 19763 14603
rect 20070 14600 20076 14612
rect 19751 14572 20076 14600
rect 19751 14569 19763 14572
rect 19705 14563 19763 14569
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 20806 14560 20812 14612
rect 20864 14600 20870 14612
rect 20990 14600 20996 14612
rect 20864 14572 20996 14600
rect 20864 14560 20870 14572
rect 20990 14560 20996 14572
rect 21048 14560 21054 14612
rect 21269 14603 21327 14609
rect 21269 14569 21281 14603
rect 21315 14600 21327 14603
rect 21358 14600 21364 14612
rect 21315 14572 21364 14600
rect 21315 14569 21327 14572
rect 21269 14563 21327 14569
rect 21358 14560 21364 14572
rect 21416 14560 21422 14612
rect 22278 14560 22284 14612
rect 22336 14600 22342 14612
rect 22741 14603 22799 14609
rect 22741 14600 22753 14603
rect 22336 14572 22753 14600
rect 22336 14560 22342 14572
rect 22741 14569 22753 14572
rect 22787 14569 22799 14603
rect 22741 14563 22799 14569
rect 26234 14560 26240 14612
rect 26292 14560 26298 14612
rect 26786 14560 26792 14612
rect 26844 14600 26850 14612
rect 27065 14603 27123 14609
rect 27065 14600 27077 14603
rect 26844 14572 27077 14600
rect 26844 14560 26850 14572
rect 27065 14569 27077 14572
rect 27111 14569 27123 14603
rect 27065 14563 27123 14569
rect 18592 14535 18650 14541
rect 14844 14504 16896 14532
rect 17052 14504 18552 14532
rect 14844 14476 14872 14504
rect 14737 14467 14795 14473
rect 14737 14462 14749 14467
rect 14660 14434 14749 14462
rect 14553 14427 14611 14433
rect 14737 14433 14749 14434
rect 14783 14433 14795 14467
rect 14737 14427 14795 14433
rect 10321 14417 10379 14423
rect 9456 14368 9628 14396
rect 9456 14356 9462 14368
rect 12066 14356 12072 14408
rect 12124 14356 12130 14408
rect 13998 14356 14004 14408
rect 14056 14396 14062 14408
rect 14200 14396 14228 14427
rect 14056 14368 14228 14396
rect 14292 14396 14320 14427
rect 14366 14396 14372 14408
rect 14292 14368 14372 14396
rect 14056 14356 14062 14368
rect 14366 14356 14372 14368
rect 14424 14356 14430 14408
rect 10229 14331 10287 14337
rect 10229 14328 10241 14331
rect 8588 14300 10241 14328
rect 7285 14291 7343 14297
rect 10229 14297 10241 14300
rect 10275 14297 10287 14331
rect 13722 14328 13728 14340
rect 10229 14291 10287 14297
rect 10336 14300 11100 14328
rect 4801 14263 4859 14269
rect 4801 14229 4813 14263
rect 4847 14260 4859 14263
rect 4890 14260 4896 14272
rect 4847 14232 4896 14260
rect 4847 14229 4859 14232
rect 4801 14223 4859 14229
rect 4890 14220 4896 14232
rect 4948 14220 4954 14272
rect 7469 14263 7527 14269
rect 7469 14229 7481 14263
rect 7515 14260 7527 14263
rect 7834 14260 7840 14272
rect 7515 14232 7840 14260
rect 7515 14229 7527 14232
rect 7469 14223 7527 14229
rect 7834 14220 7840 14232
rect 7892 14220 7898 14272
rect 8849 14263 8907 14269
rect 8849 14229 8861 14263
rect 8895 14260 8907 14263
rect 9950 14260 9956 14272
rect 8895 14232 9956 14260
rect 8895 14229 8907 14232
rect 8849 14223 8907 14229
rect 9950 14220 9956 14232
rect 10008 14260 10014 14272
rect 10336 14260 10364 14300
rect 10008 14232 10364 14260
rect 10008 14220 10014 14232
rect 10962 14220 10968 14272
rect 11020 14220 11026 14272
rect 11072 14260 11100 14300
rect 12406 14300 13728 14328
rect 12406 14260 12434 14300
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 14568 14328 14596 14427
rect 14826 14424 14832 14476
rect 14884 14424 14890 14476
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14464 14979 14467
rect 16022 14464 16028 14476
rect 14967 14436 16028 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 16022 14424 16028 14436
rect 16080 14464 16086 14476
rect 16868 14473 16896 14504
rect 16117 14467 16175 14473
rect 16117 14464 16129 14467
rect 16080 14436 16129 14464
rect 16080 14424 16086 14436
rect 16117 14433 16129 14436
rect 16163 14433 16175 14467
rect 16117 14427 16175 14433
rect 16853 14467 16911 14473
rect 16853 14433 16865 14467
rect 16899 14433 16911 14467
rect 16853 14427 16911 14433
rect 18322 14424 18328 14476
rect 18380 14424 18386 14476
rect 18524 14464 18552 14504
rect 18592 14501 18604 14535
rect 18638 14532 18650 14535
rect 19426 14532 19432 14544
rect 18638 14504 19432 14532
rect 18638 14501 18650 14504
rect 18592 14495 18650 14501
rect 19426 14492 19432 14504
rect 19484 14492 19490 14544
rect 20346 14492 20352 14544
rect 20404 14492 20410 14544
rect 22830 14492 22836 14544
rect 22888 14532 22894 14544
rect 25124 14535 25182 14541
rect 22888 14504 24072 14532
rect 22888 14492 22894 14504
rect 19058 14464 19064 14476
rect 18524 14436 19064 14464
rect 19058 14424 19064 14436
rect 19116 14424 19122 14476
rect 20364 14464 20392 14492
rect 20533 14467 20591 14473
rect 20533 14464 20545 14467
rect 19444 14436 20545 14464
rect 15197 14399 15255 14405
rect 15197 14365 15209 14399
rect 15243 14396 15255 14399
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15243 14368 15853 14396
rect 15243 14365 15255 14368
rect 15197 14359 15255 14365
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 16666 14356 16672 14408
rect 16724 14356 16730 14408
rect 18046 14356 18052 14408
rect 18104 14356 18110 14408
rect 15470 14328 15476 14340
rect 14568 14300 15476 14328
rect 15470 14288 15476 14300
rect 15528 14328 15534 14340
rect 15528 14300 17724 14328
rect 15528 14288 15534 14300
rect 11072 14232 12434 14260
rect 13449 14263 13507 14269
rect 13449 14229 13461 14263
rect 13495 14260 13507 14263
rect 14826 14260 14832 14272
rect 13495 14232 14832 14260
rect 13495 14229 13507 14232
rect 13449 14223 13507 14229
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 15286 14220 15292 14272
rect 15344 14220 15350 14272
rect 16114 14220 16120 14272
rect 16172 14260 16178 14272
rect 16942 14260 16948 14272
rect 16172 14232 16948 14260
rect 16172 14220 16178 14232
rect 16942 14220 16948 14232
rect 17000 14220 17006 14272
rect 17497 14263 17555 14269
rect 17497 14229 17509 14263
rect 17543 14260 17555 14263
rect 17586 14260 17592 14272
rect 17543 14232 17592 14260
rect 17543 14229 17555 14232
rect 17497 14223 17555 14229
rect 17586 14220 17592 14232
rect 17644 14220 17650 14272
rect 17696 14260 17724 14300
rect 18506 14260 18512 14272
rect 17696 14232 18512 14260
rect 18506 14220 18512 14232
rect 18564 14220 18570 14272
rect 18598 14220 18604 14272
rect 18656 14260 18662 14272
rect 19444 14260 19472 14436
rect 20533 14433 20545 14436
rect 20579 14433 20591 14467
rect 20533 14427 20591 14433
rect 20622 14424 20628 14476
rect 20680 14464 20686 14476
rect 22002 14464 22008 14476
rect 20680 14436 22008 14464
rect 20680 14424 20686 14436
rect 22002 14424 22008 14436
rect 22060 14424 22066 14476
rect 22370 14424 22376 14476
rect 22428 14473 22434 14476
rect 22428 14464 22440 14473
rect 23017 14467 23075 14473
rect 23017 14464 23029 14467
rect 22428 14436 22473 14464
rect 22848 14436 23029 14464
rect 22428 14427 22440 14436
rect 22428 14424 22434 14427
rect 20070 14356 20076 14408
rect 20128 14396 20134 14408
rect 20349 14399 20407 14405
rect 20349 14396 20361 14399
rect 20128 14368 20361 14396
rect 20128 14356 20134 14368
rect 20349 14365 20361 14368
rect 20395 14365 20407 14399
rect 20349 14359 20407 14365
rect 22649 14399 22707 14405
rect 22649 14365 22661 14399
rect 22695 14396 22707 14399
rect 22738 14396 22744 14408
rect 22695 14368 22744 14396
rect 22695 14365 22707 14368
rect 22649 14359 22707 14365
rect 22738 14356 22744 14368
rect 22796 14356 22802 14408
rect 18656 14232 19472 14260
rect 18656 14220 18662 14232
rect 19518 14220 19524 14272
rect 19576 14260 19582 14272
rect 19797 14263 19855 14269
rect 19797 14260 19809 14263
rect 19576 14232 19809 14260
rect 19576 14220 19582 14232
rect 19797 14229 19809 14232
rect 19843 14229 19855 14263
rect 19797 14223 19855 14229
rect 20346 14220 20352 14272
rect 20404 14260 20410 14272
rect 20717 14263 20775 14269
rect 20717 14260 20729 14263
rect 20404 14232 20729 14260
rect 20404 14220 20410 14232
rect 20717 14229 20729 14232
rect 20763 14260 20775 14263
rect 21358 14260 21364 14272
rect 20763 14232 21364 14260
rect 20763 14229 20775 14232
rect 20717 14223 20775 14229
rect 21358 14220 21364 14232
rect 21416 14260 21422 14272
rect 22646 14260 22652 14272
rect 21416 14232 22652 14260
rect 21416 14220 21422 14232
rect 22646 14220 22652 14232
rect 22704 14220 22710 14272
rect 22848 14260 22876 14436
rect 23017 14433 23029 14436
rect 23063 14433 23075 14467
rect 23017 14427 23075 14433
rect 23109 14467 23167 14473
rect 23109 14433 23121 14467
rect 23155 14433 23167 14467
rect 23109 14427 23167 14433
rect 23201 14467 23259 14473
rect 23201 14433 23213 14467
rect 23247 14464 23259 14467
rect 23290 14464 23296 14476
rect 23247 14436 23296 14464
rect 23247 14433 23259 14436
rect 23201 14427 23259 14433
rect 22922 14288 22928 14340
rect 22980 14328 22986 14340
rect 23124 14328 23152 14427
rect 23290 14424 23296 14436
rect 23348 14424 23354 14476
rect 23385 14467 23443 14473
rect 23385 14433 23397 14467
rect 23431 14464 23443 14467
rect 23566 14464 23572 14476
rect 23431 14436 23572 14464
rect 23431 14433 23443 14436
rect 23385 14427 23443 14433
rect 23566 14424 23572 14436
rect 23624 14424 23630 14476
rect 24044 14473 24072 14504
rect 25124 14501 25136 14535
rect 25170 14532 25182 14535
rect 26418 14532 26424 14544
rect 25170 14504 26424 14532
rect 25170 14501 25182 14504
rect 25124 14495 25182 14501
rect 26418 14492 26424 14504
rect 26476 14492 26482 14544
rect 24029 14467 24087 14473
rect 24029 14433 24041 14467
rect 24075 14433 24087 14467
rect 24029 14427 24087 14433
rect 23842 14356 23848 14408
rect 23900 14396 23906 14408
rect 24854 14396 24860 14408
rect 23900 14368 24860 14396
rect 23900 14356 23906 14368
rect 24854 14356 24860 14368
rect 24912 14356 24918 14408
rect 26418 14356 26424 14408
rect 26476 14356 26482 14408
rect 22980 14300 23152 14328
rect 22980 14288 22986 14300
rect 23477 14263 23535 14269
rect 23477 14260 23489 14263
rect 22848 14232 23489 14260
rect 23477 14229 23489 14232
rect 23523 14229 23535 14263
rect 23477 14223 23535 14229
rect 24394 14220 24400 14272
rect 24452 14260 24458 14272
rect 26602 14260 26608 14272
rect 24452 14232 26608 14260
rect 24452 14220 24458 14232
rect 26602 14220 26608 14232
rect 26660 14220 26666 14272
rect 552 14170 27416 14192
rect 552 14118 3756 14170
rect 3808 14118 3820 14170
rect 3872 14118 3884 14170
rect 3936 14118 3948 14170
rect 4000 14118 4012 14170
rect 4064 14118 10472 14170
rect 10524 14118 10536 14170
rect 10588 14118 10600 14170
rect 10652 14118 10664 14170
rect 10716 14118 10728 14170
rect 10780 14118 17188 14170
rect 17240 14118 17252 14170
rect 17304 14118 17316 14170
rect 17368 14118 17380 14170
rect 17432 14118 17444 14170
rect 17496 14118 23904 14170
rect 23956 14118 23968 14170
rect 24020 14118 24032 14170
rect 24084 14118 24096 14170
rect 24148 14118 24160 14170
rect 24212 14118 27416 14170
rect 552 14096 27416 14118
rect 3234 14016 3240 14068
rect 3292 14016 3298 14068
rect 4154 14056 4160 14068
rect 3528 14028 4160 14056
rect 2869 13991 2927 13997
rect 2869 13957 2881 13991
rect 2915 13988 2927 13991
rect 3528 13988 3556 14028
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 4706 14016 4712 14068
rect 4764 14056 4770 14068
rect 6181 14059 6239 14065
rect 6181 14056 6193 14059
rect 4764 14028 6193 14056
rect 4764 14016 4770 14028
rect 6181 14025 6193 14028
rect 6227 14025 6239 14059
rect 6181 14019 6239 14025
rect 4801 13991 4859 13997
rect 4801 13988 4813 13991
rect 2915 13960 3556 13988
rect 3620 13960 4813 13988
rect 2915 13957 2927 13960
rect 2869 13951 2927 13957
rect 1489 13855 1547 13861
rect 1489 13821 1501 13855
rect 1535 13852 1547 13855
rect 1535 13824 2452 13852
rect 1535 13821 1547 13824
rect 1489 13815 1547 13821
rect 2424 13796 2452 13824
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 3418 13852 3424 13864
rect 2740 13824 3424 13852
rect 2740 13812 2746 13824
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 3510 13812 3516 13864
rect 3568 13812 3574 13864
rect 3620 13861 3648 13960
rect 4801 13957 4813 13960
rect 4847 13988 4859 13991
rect 5166 13988 5172 14000
rect 4847 13960 5172 13988
rect 4847 13957 4859 13960
rect 4801 13951 4859 13957
rect 5166 13948 5172 13960
rect 5224 13948 5230 14000
rect 6196 13988 6224 14019
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 6788 14028 7328 14056
rect 6788 14016 6794 14028
rect 6196 13960 7236 13988
rect 4614 13920 4620 13932
rect 3712 13892 4620 13920
rect 3712 13861 3740 13892
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 5721 13923 5779 13929
rect 5721 13920 5733 13923
rect 4724 13892 5733 13920
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13821 3663 13855
rect 3605 13815 3663 13821
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13821 3755 13855
rect 3881 13855 3939 13861
rect 3881 13852 3893 13855
rect 3697 13815 3755 13821
rect 3804 13824 3893 13852
rect 1762 13793 1768 13796
rect 1756 13784 1768 13793
rect 1723 13756 1768 13784
rect 1756 13747 1768 13756
rect 1762 13744 1768 13747
rect 1820 13744 1826 13796
rect 2406 13744 2412 13796
rect 2464 13744 2470 13796
rect 3436 13784 3464 13812
rect 3804 13784 3832 13824
rect 3881 13821 3893 13824
rect 3927 13821 3939 13855
rect 3881 13815 3939 13821
rect 3973 13855 4031 13861
rect 3973 13821 3985 13855
rect 4019 13852 4031 13855
rect 4019 13824 4108 13852
rect 4019 13821 4031 13824
rect 3973 13815 4031 13821
rect 3436 13756 3832 13784
rect 4080 13784 4108 13824
rect 4154 13812 4160 13864
rect 4212 13812 4218 13864
rect 4246 13812 4252 13864
rect 4304 13812 4310 13864
rect 4338 13812 4344 13864
rect 4396 13852 4402 13864
rect 4724 13852 4752 13892
rect 4396 13824 4752 13852
rect 4396 13812 4402 13824
rect 4890 13812 4896 13864
rect 4948 13812 4954 13864
rect 5092 13861 5120 13892
rect 5721 13889 5733 13892
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13821 5135 13855
rect 5077 13815 5135 13821
rect 5353 13855 5411 13861
rect 5353 13821 5365 13855
rect 5399 13821 5411 13855
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 5353 13815 5411 13821
rect 5736 13824 6101 13852
rect 4264 13784 4292 13812
rect 4080 13756 4292 13784
rect 4908 13784 4936 13812
rect 5368 13784 5396 13815
rect 5736 13784 5764 13824
rect 6089 13821 6101 13824
rect 6135 13852 6147 13855
rect 6178 13852 6184 13864
rect 6135 13824 6184 13852
rect 6135 13821 6147 13824
rect 6089 13815 6147 13821
rect 6178 13812 6184 13824
rect 6236 13812 6242 13864
rect 6365 13855 6423 13861
rect 6365 13852 6377 13855
rect 6288 13824 6377 13852
rect 4908 13756 5396 13784
rect 5460 13756 5764 13784
rect 5905 13787 5963 13793
rect 1946 13676 1952 13728
rect 2004 13716 2010 13728
rect 3602 13716 3608 13728
rect 2004 13688 3608 13716
rect 2004 13676 2010 13688
rect 3602 13676 3608 13688
rect 3660 13676 3666 13728
rect 4154 13676 4160 13728
rect 4212 13716 4218 13728
rect 4341 13719 4399 13725
rect 4341 13716 4353 13719
rect 4212 13688 4353 13716
rect 4212 13676 4218 13688
rect 4341 13685 4353 13688
rect 4387 13685 4399 13719
rect 4341 13679 4399 13685
rect 5074 13676 5080 13728
rect 5132 13716 5138 13728
rect 5169 13719 5227 13725
rect 5169 13716 5181 13719
rect 5132 13688 5181 13716
rect 5132 13676 5138 13688
rect 5169 13685 5181 13688
rect 5215 13685 5227 13719
rect 5169 13679 5227 13685
rect 5258 13676 5264 13728
rect 5316 13716 5322 13728
rect 5460 13716 5488 13756
rect 5905 13753 5917 13787
rect 5951 13784 5963 13787
rect 6288 13784 6316 13824
rect 6365 13821 6377 13824
rect 6411 13852 6423 13855
rect 6914 13852 6920 13864
rect 6411 13824 6920 13852
rect 6411 13821 6423 13824
rect 6365 13815 6423 13821
rect 6914 13812 6920 13824
rect 6972 13812 6978 13864
rect 7208 13852 7236 13960
rect 7300 13929 7328 14028
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 9858 14056 9864 14068
rect 7800 14028 9864 14056
rect 7800 14016 7806 14028
rect 7558 13948 7564 14000
rect 7616 13988 7622 14000
rect 7616 13960 7880 13988
rect 7616 13948 7622 13960
rect 7285 13923 7343 13929
rect 7285 13889 7297 13923
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7852 13861 7880 13960
rect 8202 13948 8208 14000
rect 8260 13948 8266 14000
rect 7837 13855 7895 13861
rect 7208 13824 7696 13852
rect 5951 13756 6316 13784
rect 7668 13784 7696 13824
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 8294 13852 8300 13864
rect 7883 13824 8300 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 8294 13812 8300 13824
rect 8352 13852 8358 13864
rect 8864 13861 8892 14028
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 10321 14059 10379 14065
rect 10321 14025 10333 14059
rect 10367 14056 10379 14059
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 10367 14028 11989 14056
rect 10367 14025 10379 14028
rect 10321 14019 10379 14025
rect 11977 14025 11989 14028
rect 12023 14056 12035 14059
rect 12066 14056 12072 14068
rect 12023 14028 12072 14056
rect 12023 14025 12035 14028
rect 11977 14019 12035 14025
rect 10336 13988 10364 14019
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 14366 14016 14372 14068
rect 14424 14056 14430 14068
rect 15473 14059 15531 14065
rect 15473 14056 15485 14059
rect 14424 14028 15485 14056
rect 14424 14016 14430 14028
rect 15473 14025 15485 14028
rect 15519 14025 15531 14059
rect 15473 14019 15531 14025
rect 16390 14016 16396 14068
rect 16448 14016 16454 14068
rect 18598 14056 18604 14068
rect 16868 14028 18604 14056
rect 8956 13960 10364 13988
rect 15381 13991 15439 13997
rect 8665 13855 8723 13861
rect 8665 13852 8677 13855
rect 8352 13824 8677 13852
rect 8352 13812 8358 13824
rect 8665 13821 8677 13824
rect 8711 13821 8723 13855
rect 8665 13815 8723 13821
rect 8849 13855 8907 13861
rect 8849 13821 8861 13855
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 8021 13787 8079 13793
rect 7668 13756 7972 13784
rect 5951 13753 5963 13756
rect 5905 13747 5963 13753
rect 5316 13688 5488 13716
rect 5316 13676 5322 13688
rect 5534 13676 5540 13728
rect 5592 13676 5598 13728
rect 7742 13676 7748 13728
rect 7800 13676 7806 13728
rect 7944 13716 7972 13756
rect 8021 13753 8033 13787
rect 8067 13784 8079 13787
rect 8386 13784 8392 13796
rect 8067 13756 8392 13784
rect 8067 13753 8079 13756
rect 8021 13747 8079 13753
rect 8386 13744 8392 13756
rect 8444 13784 8450 13796
rect 8956 13784 8984 13960
rect 15381 13957 15393 13991
rect 15427 13988 15439 13991
rect 16666 13988 16672 14000
rect 15427 13960 16672 13988
rect 15427 13957 15439 13960
rect 15381 13951 15439 13957
rect 16666 13948 16672 13960
rect 16724 13948 16730 14000
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13920 10011 13923
rect 16868 13920 16896 14028
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 20162 14016 20168 14068
rect 20220 14016 20226 14068
rect 22002 14016 22008 14068
rect 22060 14056 22066 14068
rect 22922 14056 22928 14068
rect 22060 14028 22928 14056
rect 22060 14016 22066 14028
rect 17034 13948 17040 14000
rect 17092 13948 17098 14000
rect 18509 13991 18567 13997
rect 18509 13957 18521 13991
rect 18555 13988 18567 13991
rect 20898 13988 20904 14000
rect 18555 13960 19288 13988
rect 18555 13957 18567 13960
rect 18509 13951 18567 13957
rect 17052 13920 17080 13948
rect 9999 13892 10364 13920
rect 9999 13889 10011 13892
rect 9953 13883 10011 13889
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13852 9091 13855
rect 9674 13852 9680 13864
rect 9079 13824 9680 13852
rect 9079 13821 9091 13824
rect 9033 13815 9091 13821
rect 9674 13812 9680 13824
rect 9732 13812 9738 13864
rect 9858 13812 9864 13864
rect 9916 13812 9922 13864
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 8444 13756 8984 13784
rect 8444 13744 8450 13756
rect 9766 13744 9772 13796
rect 9824 13784 9830 13796
rect 10060 13784 10088 13815
rect 9824 13756 10088 13784
rect 9824 13744 9830 13756
rect 10134 13744 10140 13796
rect 10192 13744 10198 13796
rect 10336 13793 10364 13892
rect 15856 13892 16896 13920
rect 16960 13892 17080 13920
rect 10597 13855 10655 13861
rect 10597 13821 10609 13855
rect 10643 13852 10655 13855
rect 11974 13852 11980 13864
rect 10643 13824 11980 13852
rect 10643 13821 10655 13824
rect 10597 13815 10655 13821
rect 11532 13796 11560 13824
rect 11974 13812 11980 13824
rect 12032 13812 12038 13864
rect 14001 13855 14059 13861
rect 12406 13824 13952 13852
rect 10870 13793 10876 13796
rect 10336 13787 10395 13793
rect 10336 13756 10349 13787
rect 10337 13753 10349 13756
rect 10383 13753 10395 13787
rect 10337 13747 10395 13753
rect 10428 13756 10640 13784
rect 8478 13716 8484 13728
rect 7944 13688 8484 13716
rect 8478 13676 8484 13688
rect 8536 13716 8542 13728
rect 9398 13716 9404 13728
rect 8536 13688 9404 13716
rect 8536 13676 8542 13688
rect 9398 13676 9404 13688
rect 9456 13716 9462 13728
rect 10428 13716 10456 13756
rect 9456 13688 10456 13716
rect 9456 13676 9462 13688
rect 10502 13676 10508 13728
rect 10560 13676 10566 13728
rect 10612 13716 10640 13756
rect 10864 13747 10876 13793
rect 10870 13744 10876 13747
rect 10928 13744 10934 13796
rect 11514 13744 11520 13796
rect 11572 13744 11578 13796
rect 12406 13784 12434 13824
rect 11624 13756 12434 13784
rect 13924 13784 13952 13824
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 14090 13852 14096 13864
rect 14047 13824 14096 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 14268 13855 14326 13861
rect 14268 13821 14280 13855
rect 14314 13852 14326 13855
rect 15286 13852 15292 13864
rect 14314 13824 15292 13852
rect 14314 13821 14326 13824
rect 14268 13815 14326 13821
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 15611 13855 15669 13861
rect 15611 13852 15623 13855
rect 15396 13824 15623 13852
rect 15396 13784 15424 13824
rect 15611 13821 15623 13824
rect 15657 13852 15669 13855
rect 15856 13852 15884 13892
rect 16022 13852 16028 13864
rect 15657 13824 15884 13852
rect 15983 13824 16028 13852
rect 15657 13821 15669 13824
rect 15611 13815 15669 13821
rect 16022 13812 16028 13824
rect 16080 13812 16086 13864
rect 16114 13812 16120 13864
rect 16172 13812 16178 13864
rect 16546 13861 16574 13892
rect 16531 13855 16589 13861
rect 16531 13821 16543 13855
rect 16577 13821 16589 13855
rect 16531 13815 16589 13821
rect 16666 13812 16672 13864
rect 16724 13812 16730 13864
rect 16960 13861 16988 13892
rect 18230 13880 18236 13932
rect 18288 13920 18294 13932
rect 19260 13929 19288 13960
rect 20548 13960 20904 13988
rect 18693 13923 18751 13929
rect 18693 13920 18705 13923
rect 18288 13892 18705 13920
rect 18288 13880 18294 13892
rect 18693 13889 18705 13892
rect 18739 13889 18751 13923
rect 18693 13883 18751 13889
rect 19245 13923 19303 13929
rect 19245 13889 19257 13923
rect 19291 13889 19303 13923
rect 20548 13920 20576 13960
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 22388 13920 22416 14028
rect 22922 14016 22928 14028
rect 22980 14016 22986 14068
rect 24029 14059 24087 14065
rect 24029 14025 24041 14059
rect 24075 14056 24087 14059
rect 24302 14056 24308 14068
rect 24075 14028 24308 14056
rect 24075 14025 24087 14028
rect 24029 14019 24087 14025
rect 24302 14016 24308 14028
rect 24360 14016 24366 14068
rect 25866 14016 25872 14068
rect 25924 14056 25930 14068
rect 26973 14059 27031 14065
rect 26973 14056 26985 14059
rect 25924 14028 26985 14056
rect 25924 14016 25930 14028
rect 26973 14025 26985 14028
rect 27019 14025 27031 14059
rect 26973 14019 27031 14025
rect 26326 13988 26332 14000
rect 24596 13960 26332 13988
rect 23198 13920 23204 13932
rect 19245 13883 19303 13889
rect 19352 13892 20392 13920
rect 16761 13855 16819 13861
rect 16761 13821 16773 13855
rect 16807 13821 16819 13855
rect 16761 13815 16819 13821
rect 16944 13855 17002 13861
rect 16944 13821 16956 13855
rect 16990 13821 17002 13855
rect 16944 13815 17002 13821
rect 13924 13756 15424 13784
rect 11054 13716 11060 13728
rect 10612 13688 11060 13716
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 11330 13676 11336 13728
rect 11388 13716 11394 13728
rect 11624 13716 11652 13756
rect 15746 13744 15752 13796
rect 15804 13744 15810 13796
rect 15841 13787 15899 13793
rect 15841 13753 15853 13787
rect 15887 13753 15899 13787
rect 16776 13784 16804 13815
rect 17034 13812 17040 13864
rect 17092 13812 17098 13864
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17954 13852 17960 13864
rect 17175 13824 17960 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17954 13812 17960 13824
rect 18012 13852 18018 13864
rect 18322 13852 18328 13864
rect 18012 13824 18328 13852
rect 18012 13812 18018 13824
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 18506 13812 18512 13864
rect 18564 13852 18570 13864
rect 19352 13852 19380 13892
rect 18564 13824 19380 13852
rect 18564 13812 18570 13824
rect 19518 13812 19524 13864
rect 19576 13852 19582 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19576 13824 19717 13852
rect 19576 13812 19582 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 19794 13812 19800 13864
rect 19852 13812 19858 13864
rect 19886 13812 19892 13864
rect 19944 13812 19950 13864
rect 20073 13855 20131 13861
rect 20073 13821 20085 13855
rect 20119 13852 20131 13855
rect 20254 13852 20260 13864
rect 20119 13824 20260 13852
rect 20119 13821 20131 13824
rect 20073 13815 20131 13821
rect 20254 13812 20260 13824
rect 20312 13812 20318 13864
rect 17218 13784 17224 13796
rect 15841 13747 15899 13753
rect 16408 13756 17224 13784
rect 11388 13688 11652 13716
rect 11388 13676 11394 13688
rect 12066 13676 12072 13728
rect 12124 13716 12130 13728
rect 15856 13716 15884 13747
rect 16408 13716 16436 13756
rect 17218 13744 17224 13756
rect 17276 13744 17282 13796
rect 17396 13787 17454 13793
rect 17396 13753 17408 13787
rect 17442 13784 17454 13787
rect 17586 13784 17592 13796
rect 17442 13756 17592 13784
rect 17442 13753 17454 13756
rect 17396 13747 17454 13753
rect 17586 13744 17592 13756
rect 17644 13744 17650 13796
rect 18598 13744 18604 13796
rect 18656 13784 18662 13796
rect 19242 13784 19248 13796
rect 18656 13756 19248 13784
rect 18656 13744 18662 13756
rect 19242 13744 19248 13756
rect 19300 13744 19306 13796
rect 20364 13784 20392 13892
rect 20456 13892 20576 13920
rect 21928 13892 22416 13920
rect 22664 13892 23204 13920
rect 20456 13861 20484 13892
rect 20441 13855 20499 13861
rect 20441 13821 20453 13855
rect 20487 13821 20499 13855
rect 20441 13815 20499 13821
rect 20530 13812 20536 13864
rect 20588 13812 20594 13864
rect 20625 13855 20683 13861
rect 20625 13821 20637 13855
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 20640 13784 20668 13815
rect 20714 13812 20720 13864
rect 20772 13852 20778 13864
rect 21082 13861 21088 13864
rect 20809 13855 20867 13861
rect 20809 13852 20821 13855
rect 20772 13824 20821 13852
rect 20772 13812 20778 13824
rect 20809 13821 20821 13824
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 20901 13855 20959 13861
rect 20901 13821 20913 13855
rect 20947 13821 20959 13855
rect 20901 13815 20959 13821
rect 21049 13855 21088 13861
rect 21049 13821 21061 13855
rect 21049 13815 21088 13821
rect 20364 13756 20668 13784
rect 12124 13688 16436 13716
rect 12124 13676 12130 13688
rect 19426 13676 19432 13728
rect 19484 13676 19490 13728
rect 20254 13676 20260 13728
rect 20312 13716 20318 13728
rect 20806 13716 20812 13728
rect 20312 13688 20812 13716
rect 20312 13676 20318 13688
rect 20806 13676 20812 13688
rect 20864 13716 20870 13728
rect 20916 13716 20944 13815
rect 21082 13812 21088 13815
rect 21140 13812 21146 13864
rect 21174 13812 21180 13864
rect 21232 13812 21238 13864
rect 21266 13812 21272 13864
rect 21324 13812 21330 13864
rect 21358 13812 21364 13864
rect 21416 13861 21422 13864
rect 21416 13852 21424 13861
rect 21637 13855 21695 13861
rect 21416 13824 21461 13852
rect 21416 13815 21424 13824
rect 21637 13821 21649 13855
rect 21683 13852 21695 13855
rect 21726 13852 21732 13864
rect 21683 13824 21732 13852
rect 21683 13821 21695 13824
rect 21637 13815 21695 13821
rect 21416 13812 21422 13815
rect 21726 13812 21732 13824
rect 21784 13812 21790 13864
rect 21818 13812 21824 13864
rect 21876 13812 21882 13864
rect 21928 13861 21956 13892
rect 21913 13855 21971 13861
rect 21913 13821 21925 13855
rect 21959 13821 21971 13855
rect 21913 13815 21971 13821
rect 22005 13855 22063 13861
rect 22005 13821 22017 13855
rect 22051 13852 22063 13855
rect 22094 13852 22100 13864
rect 22051 13824 22100 13852
rect 22051 13821 22063 13824
rect 22005 13815 22063 13821
rect 22094 13812 22100 13824
rect 22152 13812 22158 13864
rect 22664 13852 22692 13892
rect 23198 13880 23204 13892
rect 23256 13880 23262 13932
rect 24486 13920 24492 13932
rect 24320 13892 24492 13920
rect 22296 13824 22692 13852
rect 22296 13793 22324 13824
rect 22738 13812 22744 13864
rect 22796 13852 22802 13864
rect 24210 13861 24216 13864
rect 22925 13855 22983 13861
rect 22925 13852 22937 13855
rect 22796 13824 22937 13852
rect 22796 13812 22802 13824
rect 22925 13821 22937 13824
rect 22971 13821 22983 13855
rect 24167 13855 24216 13861
rect 24167 13852 24179 13855
rect 22925 13815 22983 13821
rect 23124 13824 24179 13852
rect 22281 13787 22339 13793
rect 22281 13753 22293 13787
rect 22327 13753 22339 13787
rect 22281 13747 22339 13753
rect 22646 13744 22652 13796
rect 22704 13784 22710 13796
rect 23124 13784 23152 13824
rect 24167 13821 24179 13824
rect 24213 13821 24216 13855
rect 24167 13815 24216 13821
rect 24210 13812 24216 13815
rect 24268 13812 24274 13864
rect 24320 13861 24348 13892
rect 24486 13880 24492 13892
rect 24544 13880 24550 13932
rect 24305 13855 24363 13861
rect 24305 13821 24317 13855
rect 24351 13821 24363 13855
rect 24305 13815 24363 13821
rect 24394 13812 24400 13864
rect 24452 13812 24458 13864
rect 24596 13861 24624 13960
rect 26326 13948 26332 13960
rect 26384 13948 26390 14000
rect 26510 13948 26516 14000
rect 26568 13948 26574 14000
rect 26528 13920 26556 13948
rect 25608 13892 26556 13920
rect 24580 13855 24638 13861
rect 24580 13821 24592 13855
rect 24626 13821 24638 13855
rect 24580 13815 24638 13821
rect 24673 13855 24731 13861
rect 24673 13821 24685 13855
rect 24719 13821 24731 13855
rect 24673 13815 24731 13821
rect 22704 13756 23152 13784
rect 22704 13744 22710 13756
rect 20864 13688 20944 13716
rect 21545 13719 21603 13725
rect 20864 13676 20870 13688
rect 21545 13685 21557 13719
rect 21591 13716 21603 13719
rect 21726 13716 21732 13728
rect 21591 13688 21732 13716
rect 21591 13685 21603 13688
rect 21545 13679 21603 13685
rect 21726 13676 21732 13688
rect 21784 13676 21790 13728
rect 22370 13676 22376 13728
rect 22428 13676 22434 13728
rect 23198 13676 23204 13728
rect 23256 13716 23262 13728
rect 24688 13716 24716 13815
rect 24946 13812 24952 13864
rect 25004 13812 25010 13864
rect 25608 13861 25636 13892
rect 25593 13855 25651 13861
rect 25593 13852 25605 13855
rect 25056 13824 25605 13852
rect 25056 13716 25084 13824
rect 25593 13821 25605 13824
rect 25639 13821 25651 13855
rect 25593 13815 25651 13821
rect 25686 13855 25744 13861
rect 25686 13821 25698 13855
rect 25732 13821 25744 13855
rect 25686 13815 25744 13821
rect 25869 13855 25927 13861
rect 25869 13821 25881 13855
rect 25915 13821 25927 13855
rect 25869 13815 25927 13821
rect 25700 13784 25728 13815
rect 25516 13756 25728 13784
rect 25884 13784 25912 13815
rect 25958 13812 25964 13864
rect 26016 13812 26022 13864
rect 26050 13812 26056 13864
rect 26108 13861 26114 13864
rect 26344 13861 26372 13892
rect 26510 13861 26516 13864
rect 26108 13852 26116 13861
rect 26329 13855 26387 13861
rect 26108 13824 26153 13852
rect 26108 13815 26116 13824
rect 26329 13821 26341 13855
rect 26375 13821 26387 13855
rect 26329 13815 26387 13821
rect 26477 13855 26516 13861
rect 26477 13821 26489 13855
rect 26477 13815 26516 13821
rect 26108 13812 26114 13815
rect 26510 13812 26516 13815
rect 26568 13812 26574 13864
rect 26602 13812 26608 13864
rect 26660 13812 26666 13864
rect 26694 13812 26700 13864
rect 26752 13812 26758 13864
rect 26786 13812 26792 13864
rect 26844 13861 26850 13864
rect 26844 13852 26852 13861
rect 26844 13824 26889 13852
rect 26844 13815 26852 13824
rect 26844 13812 26850 13815
rect 26620 13784 26648 13812
rect 25884 13756 26648 13784
rect 23256 13688 25084 13716
rect 23256 13676 23262 13688
rect 25406 13676 25412 13728
rect 25464 13716 25470 13728
rect 25516 13725 25544 13756
rect 25501 13719 25559 13725
rect 25501 13716 25513 13719
rect 25464 13688 25513 13716
rect 25464 13676 25470 13688
rect 25501 13685 25513 13688
rect 25547 13685 25559 13719
rect 25501 13679 25559 13685
rect 26234 13676 26240 13728
rect 26292 13676 26298 13728
rect 552 13626 27576 13648
rect 552 13574 7114 13626
rect 7166 13574 7178 13626
rect 7230 13574 7242 13626
rect 7294 13574 7306 13626
rect 7358 13574 7370 13626
rect 7422 13574 13830 13626
rect 13882 13574 13894 13626
rect 13946 13574 13958 13626
rect 14010 13574 14022 13626
rect 14074 13574 14086 13626
rect 14138 13574 20546 13626
rect 20598 13574 20610 13626
rect 20662 13574 20674 13626
rect 20726 13574 20738 13626
rect 20790 13574 20802 13626
rect 20854 13574 27262 13626
rect 27314 13574 27326 13626
rect 27378 13574 27390 13626
rect 27442 13574 27454 13626
rect 27506 13574 27518 13626
rect 27570 13574 27576 13626
rect 552 13552 27576 13574
rect 1765 13515 1823 13521
rect 1765 13481 1777 13515
rect 1811 13512 1823 13515
rect 4154 13512 4160 13524
rect 1811 13484 4160 13512
rect 1811 13481 1823 13484
rect 1765 13475 1823 13481
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 5902 13512 5908 13524
rect 5368 13484 5908 13512
rect 1946 13404 1952 13456
rect 2004 13404 2010 13456
rect 2777 13447 2835 13453
rect 2777 13444 2789 13447
rect 2332 13416 2789 13444
rect 2332 13385 2360 13416
rect 2777 13413 2789 13416
rect 2823 13413 2835 13447
rect 2777 13407 2835 13413
rect 3602 13404 3608 13456
rect 3660 13444 3666 13456
rect 3973 13447 4031 13453
rect 3973 13444 3985 13447
rect 3660 13416 3985 13444
rect 3660 13404 3666 13416
rect 3973 13413 3985 13416
rect 4019 13413 4031 13447
rect 3973 13407 4031 13413
rect 5258 13404 5264 13456
rect 5316 13404 5322 13456
rect 5368 13453 5396 13484
rect 5902 13472 5908 13484
rect 5960 13472 5966 13524
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 6972 13484 8248 13512
rect 6972 13472 6978 13484
rect 5534 13453 5540 13456
rect 5353 13447 5411 13453
rect 5353 13413 5365 13447
rect 5399 13413 5411 13447
rect 5353 13407 5411 13413
rect 5491 13447 5540 13453
rect 5491 13413 5503 13447
rect 5537 13413 5540 13447
rect 5491 13407 5540 13413
rect 5534 13404 5540 13407
rect 5592 13404 5598 13456
rect 7558 13444 7564 13456
rect 6564 13416 7564 13444
rect 1673 13379 1731 13385
rect 1673 13345 1685 13379
rect 1719 13345 1731 13379
rect 1673 13339 1731 13345
rect 2317 13379 2375 13385
rect 2317 13345 2329 13379
rect 2363 13345 2375 13379
rect 2317 13339 2375 13345
rect 2409 13379 2467 13385
rect 2409 13345 2421 13379
rect 2455 13345 2467 13379
rect 2409 13339 2467 13345
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 2547 13348 2636 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 1688 13240 1716 13339
rect 1876 13311 1934 13317
rect 1876 13277 1888 13311
rect 1922 13308 1934 13311
rect 2222 13308 2228 13320
rect 1922 13280 2228 13308
rect 1922 13277 1934 13280
rect 1876 13271 1934 13277
rect 2222 13268 2228 13280
rect 2280 13308 2286 13320
rect 2424 13308 2452 13339
rect 2280 13280 2452 13308
rect 2280 13268 2286 13280
rect 2608 13240 2636 13348
rect 2682 13336 2688 13388
rect 2740 13336 2746 13388
rect 2958 13336 2964 13388
rect 3016 13376 3022 13388
rect 3697 13379 3755 13385
rect 3697 13376 3709 13379
rect 3016 13348 3709 13376
rect 3016 13336 3022 13348
rect 3697 13345 3709 13348
rect 3743 13345 3755 13379
rect 3697 13339 3755 13345
rect 5166 13336 5172 13388
rect 5224 13336 5230 13388
rect 6564 13385 6592 13416
rect 7558 13404 7564 13416
rect 7616 13404 7622 13456
rect 8220 13444 8248 13484
rect 8294 13472 8300 13524
rect 8352 13472 8358 13524
rect 10781 13515 10839 13521
rect 10244 13484 10640 13512
rect 8220 13416 8524 13444
rect 5813 13379 5871 13385
rect 5813 13376 5825 13379
rect 5644 13348 5825 13376
rect 5644 13320 5672 13348
rect 5813 13345 5825 13348
rect 5859 13345 5871 13379
rect 5813 13339 5871 13345
rect 5997 13379 6055 13385
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 6549 13379 6607 13385
rect 6043 13348 6408 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 3418 13268 3424 13320
rect 3476 13268 3482 13320
rect 3881 13311 3939 13317
rect 3881 13277 3893 13311
rect 3927 13308 3939 13311
rect 4798 13308 4804 13320
rect 3927 13280 4804 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 5626 13268 5632 13320
rect 5684 13308 5690 13320
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 5684 13280 6285 13308
rect 5684 13268 5690 13280
rect 6273 13277 6285 13280
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 3513 13243 3571 13249
rect 3513 13240 3525 13243
rect 1688 13212 2544 13240
rect 2608 13212 3525 13240
rect 2038 13132 2044 13184
rect 2096 13132 2102 13184
rect 2516 13172 2544 13212
rect 3513 13209 3525 13212
rect 3559 13209 3571 13243
rect 3513 13203 3571 13209
rect 5074 13200 5080 13252
rect 5132 13240 5138 13252
rect 6380 13249 6408 13348
rect 6549 13345 6561 13379
rect 6595 13345 6607 13379
rect 6549 13339 6607 13345
rect 6822 13336 6828 13388
rect 6880 13376 6886 13388
rect 7190 13385 7196 13388
rect 6917 13379 6975 13385
rect 6917 13376 6929 13379
rect 6880 13348 6929 13376
rect 6880 13336 6886 13348
rect 6917 13345 6929 13348
rect 6963 13345 6975 13379
rect 6917 13339 6975 13345
rect 7184 13339 7196 13385
rect 7190 13336 7196 13339
rect 7248 13336 7254 13388
rect 8496 13385 8524 13416
rect 8389 13379 8447 13385
rect 8389 13376 8401 13379
rect 7944 13348 8401 13376
rect 6365 13243 6423 13249
rect 6365 13240 6377 13243
rect 5132 13212 6377 13240
rect 5132 13200 5138 13212
rect 6365 13209 6377 13212
rect 6411 13209 6423 13243
rect 6365 13203 6423 13209
rect 3326 13172 3332 13184
rect 2516 13144 3332 13172
rect 3326 13132 3332 13144
rect 3384 13132 3390 13184
rect 3973 13175 4031 13181
rect 3973 13141 3985 13175
rect 4019 13172 4031 13175
rect 4154 13172 4160 13184
rect 4019 13144 4160 13172
rect 4019 13141 4031 13144
rect 3973 13135 4031 13141
rect 4154 13132 4160 13144
rect 4212 13132 4218 13184
rect 4982 13132 4988 13184
rect 5040 13132 5046 13184
rect 6733 13175 6791 13181
rect 6733 13141 6745 13175
rect 6779 13172 6791 13175
rect 7558 13172 7564 13184
rect 6779 13144 7564 13172
rect 6779 13141 6791 13144
rect 6733 13135 6791 13141
rect 7558 13132 7564 13144
rect 7616 13172 7622 13184
rect 7944 13172 7972 13348
rect 8389 13345 8401 13348
rect 8435 13345 8447 13379
rect 8389 13339 8447 13345
rect 8481 13379 8539 13385
rect 8481 13345 8493 13379
rect 8527 13345 8539 13379
rect 8481 13339 8539 13345
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 9953 13379 10011 13385
rect 9953 13376 9965 13379
rect 9732 13348 9965 13376
rect 9732 13336 9738 13348
rect 9953 13345 9965 13348
rect 9999 13376 10011 13379
rect 10244 13376 10272 13484
rect 10502 13444 10508 13456
rect 10336 13416 10508 13444
rect 10336 13385 10364 13416
rect 10502 13404 10508 13416
rect 10560 13404 10566 13456
rect 10612 13444 10640 13484
rect 10781 13481 10793 13515
rect 10827 13512 10839 13515
rect 10870 13512 10876 13524
rect 10827 13484 10876 13512
rect 10827 13481 10839 13484
rect 10781 13475 10839 13481
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 11330 13512 11336 13524
rect 10980 13484 11336 13512
rect 10980 13444 11008 13484
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 15470 13512 15476 13524
rect 15304 13484 15476 13512
rect 12713 13447 12771 13453
rect 12713 13444 12725 13447
rect 10612 13416 11008 13444
rect 11256 13416 12725 13444
rect 9999 13348 10272 13376
rect 10321 13379 10379 13385
rect 9999 13345 10011 13348
rect 9953 13339 10011 13345
rect 10321 13345 10333 13379
rect 10367 13345 10379 13379
rect 10321 13339 10379 13345
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13376 10471 13379
rect 10870 13376 10876 13388
rect 10459 13348 10876 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 11054 13336 11060 13388
rect 11112 13336 11118 13388
rect 11256 13385 11284 13416
rect 12713 13413 12725 13416
rect 12759 13413 12771 13447
rect 15304 13444 15332 13484
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 15746 13472 15752 13524
rect 15804 13512 15810 13524
rect 16117 13515 16175 13521
rect 16117 13512 16129 13515
rect 15804 13484 16129 13512
rect 15804 13472 15810 13484
rect 16117 13481 16129 13484
rect 16163 13481 16175 13515
rect 16117 13475 16175 13481
rect 17681 13515 17739 13521
rect 17681 13481 17693 13515
rect 17727 13512 17739 13515
rect 18046 13512 18052 13524
rect 17727 13484 18052 13512
rect 17727 13481 17739 13484
rect 17681 13475 17739 13481
rect 18046 13472 18052 13484
rect 18104 13472 18110 13524
rect 18138 13472 18144 13524
rect 18196 13512 18202 13524
rect 18601 13515 18659 13521
rect 18601 13512 18613 13515
rect 18196 13484 18613 13512
rect 18196 13472 18202 13484
rect 18601 13481 18613 13484
rect 18647 13481 18659 13515
rect 18601 13475 18659 13481
rect 21082 13472 21088 13524
rect 21140 13472 21146 13524
rect 24857 13515 24915 13521
rect 24857 13481 24869 13515
rect 24903 13512 24915 13515
rect 24946 13512 24952 13524
rect 24903 13484 24952 13512
rect 24903 13481 24915 13484
rect 24857 13475 24915 13481
rect 24946 13472 24952 13484
rect 25004 13472 25010 13524
rect 18230 13444 18236 13456
rect 12713 13407 12771 13413
rect 15212 13416 15332 13444
rect 17972 13416 18236 13444
rect 11205 13379 11284 13385
rect 11205 13345 11217 13379
rect 11251 13348 11284 13379
rect 11251 13345 11263 13348
rect 11205 13339 11263 13345
rect 11330 13336 11336 13388
rect 11388 13336 11394 13388
rect 11425 13379 11483 13385
rect 11425 13345 11437 13379
rect 11471 13345 11483 13379
rect 11425 13339 11483 13345
rect 11563 13379 11621 13385
rect 11563 13345 11575 13379
rect 11609 13376 11621 13379
rect 12158 13376 12164 13388
rect 11609 13348 12164 13376
rect 11609 13345 11621 13348
rect 11563 13339 11621 13345
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 10505 13311 10563 13317
rect 10505 13308 10517 13311
rect 9824 13280 10517 13308
rect 9824 13268 9830 13280
rect 10505 13277 10517 13280
rect 10551 13277 10563 13311
rect 10505 13271 10563 13277
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13277 10655 13311
rect 10597 13271 10655 13277
rect 8757 13243 8815 13249
rect 8757 13209 8769 13243
rect 8803 13240 8815 13243
rect 9674 13240 9680 13252
rect 8803 13212 9680 13240
rect 8803 13209 8815 13212
rect 8757 13203 8815 13209
rect 9674 13200 9680 13212
rect 9732 13200 9738 13252
rect 10612 13240 10640 13271
rect 10686 13268 10692 13320
rect 10744 13308 10750 13320
rect 11440 13308 11468 13339
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 14829 13379 14887 13385
rect 14829 13345 14841 13379
rect 14875 13345 14887 13379
rect 14829 13339 14887 13345
rect 14921 13379 14979 13385
rect 14921 13345 14933 13379
rect 14967 13345 14979 13379
rect 14921 13339 14979 13345
rect 10744 13280 11468 13308
rect 10744 13268 10750 13280
rect 13354 13268 13360 13320
rect 13412 13268 13418 13320
rect 14274 13268 14280 13320
rect 14332 13268 14338 13320
rect 9784 13212 10640 13240
rect 14844 13240 14872 13339
rect 14936 13308 14964 13339
rect 15010 13336 15016 13388
rect 15068 13336 15074 13388
rect 15212 13385 15240 13416
rect 17972 13385 18000 13416
rect 18230 13404 18236 13416
rect 18288 13404 18294 13456
rect 19334 13444 19340 13456
rect 18340 13416 19340 13444
rect 18340 13388 18368 13416
rect 19334 13404 19340 13416
rect 19392 13404 19398 13456
rect 21904 13447 21962 13453
rect 19720 13416 21220 13444
rect 15197 13379 15255 13385
rect 15197 13345 15209 13379
rect 15243 13345 15255 13379
rect 15197 13339 15255 13345
rect 17957 13379 18015 13385
rect 17957 13345 17969 13379
rect 18003 13345 18015 13379
rect 17957 13339 18015 13345
rect 18046 13336 18052 13388
rect 18104 13336 18110 13388
rect 18138 13336 18144 13388
rect 18196 13336 18202 13388
rect 18322 13336 18328 13388
rect 18380 13336 18386 13388
rect 18417 13379 18475 13385
rect 18417 13345 18429 13379
rect 18463 13345 18475 13379
rect 18417 13339 18475 13345
rect 15102 13308 15108 13320
rect 14936 13280 15108 13308
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 15841 13311 15899 13317
rect 15841 13308 15853 13311
rect 15528 13280 15853 13308
rect 15528 13268 15534 13280
rect 15841 13277 15853 13280
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 16666 13268 16672 13320
rect 16724 13268 16730 13320
rect 16942 13268 16948 13320
rect 17000 13268 17006 13320
rect 17218 13268 17224 13320
rect 17276 13308 17282 13320
rect 18432 13308 18460 13339
rect 19426 13336 19432 13388
rect 19484 13376 19490 13388
rect 19720 13385 19748 13416
rect 21192 13388 21220 13416
rect 21904 13413 21916 13447
rect 21950 13444 21962 13447
rect 22370 13444 22376 13456
rect 21950 13416 22376 13444
rect 21950 13413 21962 13416
rect 21904 13407 21962 13413
rect 22370 13404 22376 13416
rect 22428 13404 22434 13456
rect 19978 13385 19984 13388
rect 19521 13379 19579 13385
rect 19521 13376 19533 13379
rect 19484 13348 19533 13376
rect 19484 13336 19490 13348
rect 19521 13345 19533 13348
rect 19567 13345 19579 13379
rect 19521 13339 19579 13345
rect 19705 13379 19763 13385
rect 19705 13345 19717 13379
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 19972 13339 19984 13385
rect 19978 13336 19984 13339
rect 20036 13336 20042 13388
rect 21174 13336 21180 13388
rect 21232 13376 21238 13388
rect 21634 13376 21640 13388
rect 21232 13348 21640 13376
rect 21232 13336 21238 13348
rect 21634 13336 21640 13348
rect 21692 13376 21698 13388
rect 22830 13376 22836 13388
rect 21692 13348 22836 13376
rect 21692 13336 21698 13348
rect 22830 13336 22836 13348
rect 22888 13376 22894 13388
rect 23744 13379 23802 13385
rect 22888 13348 23520 13376
rect 22888 13336 22894 13348
rect 23492 13317 23520 13348
rect 23744 13345 23756 13379
rect 23790 13376 23802 13379
rect 24949 13379 25007 13385
rect 24949 13376 24961 13379
rect 23790 13348 24961 13376
rect 23790 13345 23802 13348
rect 23744 13339 23802 13345
rect 24949 13345 24961 13348
rect 24995 13345 25007 13379
rect 24949 13339 25007 13345
rect 26510 13336 26516 13388
rect 26568 13376 26574 13388
rect 26973 13379 27031 13385
rect 26973 13376 26985 13379
rect 26568 13348 26985 13376
rect 26568 13336 26574 13348
rect 26973 13345 26985 13348
rect 27019 13345 27031 13379
rect 26973 13339 27031 13345
rect 17276 13280 18460 13308
rect 23477 13311 23535 13317
rect 17276 13268 17282 13280
rect 23477 13277 23489 13311
rect 23523 13277 23535 13311
rect 23477 13271 23535 13277
rect 25222 13268 25228 13320
rect 25280 13308 25286 13320
rect 25501 13311 25559 13317
rect 25501 13308 25513 13311
rect 25280 13280 25513 13308
rect 25280 13268 25286 13280
rect 25501 13277 25513 13280
rect 25547 13277 25559 13311
rect 25501 13271 25559 13277
rect 14844 13212 14964 13240
rect 7616 13144 7972 13172
rect 7616 13132 7622 13144
rect 8386 13132 8392 13184
rect 8444 13132 8450 13184
rect 8846 13132 8852 13184
rect 8904 13172 8910 13184
rect 9784 13181 9812 13212
rect 9769 13175 9827 13181
rect 9769 13172 9781 13175
rect 8904 13144 9781 13172
rect 8904 13132 8910 13144
rect 9769 13141 9781 13144
rect 9815 13141 9827 13175
rect 9769 13135 9827 13141
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10778 13172 10784 13184
rect 10100 13144 10784 13172
rect 10100 13132 10106 13144
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 11698 13132 11704 13184
rect 11756 13132 11762 13184
rect 13630 13132 13636 13184
rect 13688 13132 13694 13184
rect 14366 13132 14372 13184
rect 14424 13172 14430 13184
rect 14553 13175 14611 13181
rect 14553 13172 14565 13175
rect 14424 13144 14565 13172
rect 14424 13132 14430 13144
rect 14553 13141 14565 13144
rect 14599 13141 14611 13175
rect 14936 13172 14964 13212
rect 15289 13175 15347 13181
rect 15289 13172 15301 13175
rect 14936 13144 15301 13172
rect 14553 13135 14611 13141
rect 15289 13141 15301 13144
rect 15335 13141 15347 13175
rect 15289 13135 15347 13141
rect 17586 13132 17592 13184
rect 17644 13132 17650 13184
rect 18966 13132 18972 13184
rect 19024 13132 19030 13184
rect 23017 13175 23075 13181
rect 23017 13141 23029 13175
rect 23063 13172 23075 13175
rect 23474 13172 23480 13184
rect 23063 13144 23480 13172
rect 23063 13141 23075 13144
rect 23017 13135 23075 13141
rect 23474 13132 23480 13144
rect 23532 13132 23538 13184
rect 25774 13132 25780 13184
rect 25832 13172 25838 13184
rect 26421 13175 26479 13181
rect 26421 13172 26433 13175
rect 25832 13144 26433 13172
rect 25832 13132 25838 13144
rect 26421 13141 26433 13144
rect 26467 13141 26479 13175
rect 26421 13135 26479 13141
rect 552 13082 27416 13104
rect 552 13030 3756 13082
rect 3808 13030 3820 13082
rect 3872 13030 3884 13082
rect 3936 13030 3948 13082
rect 4000 13030 4012 13082
rect 4064 13030 10472 13082
rect 10524 13030 10536 13082
rect 10588 13030 10600 13082
rect 10652 13030 10664 13082
rect 10716 13030 10728 13082
rect 10780 13030 17188 13082
rect 17240 13030 17252 13082
rect 17304 13030 17316 13082
rect 17368 13030 17380 13082
rect 17432 13030 17444 13082
rect 17496 13030 23904 13082
rect 23956 13030 23968 13082
rect 24020 13030 24032 13082
rect 24084 13030 24096 13082
rect 24148 13030 24160 13082
rect 24212 13030 27416 13082
rect 552 13008 27416 13030
rect 2958 12928 2964 12980
rect 3016 12928 3022 12980
rect 3418 12928 3424 12980
rect 3476 12968 3482 12980
rect 4157 12971 4215 12977
rect 4157 12968 4169 12971
rect 3476 12940 4169 12968
rect 3476 12928 3482 12940
rect 4157 12937 4169 12940
rect 4203 12968 4215 12971
rect 4341 12971 4399 12977
rect 4203 12940 4292 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 2777 12903 2835 12909
rect 2777 12869 2789 12903
rect 2823 12900 2835 12903
rect 3436 12900 3464 12928
rect 2823 12872 3464 12900
rect 4264 12900 4292 12940
rect 4341 12937 4353 12971
rect 4387 12968 4399 12971
rect 5074 12968 5080 12980
rect 4387 12940 5080 12968
rect 4387 12937 4399 12940
rect 4341 12931 4399 12937
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 7190 12928 7196 12980
rect 7248 12968 7254 12980
rect 7377 12971 7435 12977
rect 7377 12968 7389 12971
rect 7248 12940 7389 12968
rect 7248 12928 7254 12940
rect 7377 12937 7389 12940
rect 7423 12937 7435 12971
rect 10870 12968 10876 12980
rect 7377 12931 7435 12937
rect 7484 12940 10876 12968
rect 4264 12872 4476 12900
rect 2823 12869 2835 12872
rect 2777 12863 2835 12869
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 2406 12764 2412 12776
rect 1443 12736 2412 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 2406 12724 2412 12736
rect 2464 12724 2470 12776
rect 2884 12773 2912 12872
rect 3602 12792 3608 12844
rect 3660 12832 3666 12844
rect 4448 12841 4476 12872
rect 4706 12860 4712 12912
rect 4764 12860 4770 12912
rect 6454 12860 6460 12912
rect 6512 12900 6518 12912
rect 6822 12900 6828 12912
rect 6512 12872 6828 12900
rect 6512 12860 6518 12872
rect 6822 12860 6828 12872
rect 6880 12900 6886 12912
rect 7484 12900 7512 12940
rect 10870 12928 10876 12940
rect 10928 12968 10934 12980
rect 11057 12971 11115 12977
rect 11057 12968 11069 12971
rect 10928 12940 11069 12968
rect 10928 12928 10934 12940
rect 11057 12937 11069 12940
rect 11103 12968 11115 12971
rect 11790 12968 11796 12980
rect 11103 12940 11796 12968
rect 11103 12937 11115 12940
rect 11057 12931 11115 12937
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 13170 12928 13176 12980
rect 13228 12968 13234 12980
rect 13228 12940 15148 12968
rect 13228 12928 13234 12940
rect 6880 12872 7512 12900
rect 7653 12903 7711 12909
rect 6880 12860 6886 12872
rect 7653 12869 7665 12903
rect 7699 12900 7711 12903
rect 7742 12900 7748 12912
rect 7699 12872 7748 12900
rect 7699 12869 7711 12872
rect 7653 12863 7711 12869
rect 7742 12860 7748 12872
rect 7800 12860 7806 12912
rect 8386 12860 8392 12912
rect 8444 12860 8450 12912
rect 10962 12900 10968 12912
rect 9140 12872 10968 12900
rect 4065 12835 4123 12841
rect 4065 12832 4077 12835
rect 3660 12804 4077 12832
rect 3660 12792 3666 12804
rect 4065 12801 4077 12804
rect 4111 12801 4123 12835
rect 4065 12795 4123 12801
rect 4433 12835 4491 12841
rect 4433 12801 4445 12835
rect 4479 12801 4491 12835
rect 8404 12832 8432 12860
rect 8662 12832 8668 12844
rect 4433 12795 4491 12801
rect 7852 12804 8668 12832
rect 2869 12767 2927 12773
rect 2869 12733 2881 12767
rect 2915 12733 2927 12767
rect 3418 12764 3424 12776
rect 2869 12727 2927 12733
rect 2976 12736 3424 12764
rect 1664 12699 1722 12705
rect 1664 12665 1676 12699
rect 1710 12696 1722 12699
rect 2038 12696 2044 12708
rect 1710 12668 2044 12696
rect 1710 12665 1722 12668
rect 1664 12659 1722 12665
rect 2038 12656 2044 12668
rect 2096 12656 2102 12708
rect 2682 12656 2688 12708
rect 2740 12696 2746 12708
rect 2976 12696 3004 12736
rect 3418 12724 3424 12736
rect 3476 12724 3482 12776
rect 3694 12724 3700 12776
rect 3752 12764 3758 12776
rect 3789 12767 3847 12773
rect 3789 12764 3801 12767
rect 3752 12736 3801 12764
rect 3752 12724 3758 12736
rect 3789 12733 3801 12736
rect 3835 12733 3847 12767
rect 3789 12727 3847 12733
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12733 3939 12767
rect 3881 12727 3939 12733
rect 3973 12767 4031 12773
rect 3973 12733 3985 12767
rect 4019 12764 4031 12767
rect 4154 12764 4160 12776
rect 4019 12736 4160 12764
rect 4019 12733 4031 12736
rect 3973 12727 4031 12733
rect 2740 12668 3004 12696
rect 2740 12656 2746 12668
rect 3326 12656 3332 12708
rect 3384 12696 3390 12708
rect 3896 12696 3924 12727
rect 4154 12724 4160 12736
rect 4212 12764 4218 12776
rect 4617 12767 4675 12773
rect 4617 12764 4629 12767
rect 4212 12736 4629 12764
rect 4212 12724 4218 12736
rect 4617 12733 4629 12736
rect 4663 12733 4675 12767
rect 4617 12727 4675 12733
rect 4709 12767 4767 12773
rect 4709 12733 4721 12767
rect 4755 12733 4767 12767
rect 4709 12727 4767 12733
rect 4893 12767 4951 12773
rect 4893 12733 4905 12767
rect 4939 12764 4951 12767
rect 6086 12764 6092 12776
rect 4939 12736 6092 12764
rect 4939 12733 4951 12736
rect 4893 12727 4951 12733
rect 4338 12696 4344 12708
rect 3384 12668 4344 12696
rect 3384 12656 3390 12668
rect 4338 12656 4344 12668
rect 4396 12656 4402 12708
rect 3234 12588 3240 12640
rect 3292 12588 3298 12640
rect 3418 12588 3424 12640
rect 3476 12588 3482 12640
rect 3694 12588 3700 12640
rect 3752 12628 3758 12640
rect 4724 12628 4752 12727
rect 6086 12724 6092 12736
rect 6144 12764 6150 12776
rect 6730 12764 6736 12776
rect 6144 12736 6736 12764
rect 6144 12724 6150 12736
rect 6730 12724 6736 12736
rect 6788 12724 6794 12776
rect 7558 12724 7564 12776
rect 7616 12724 7622 12776
rect 7852 12773 7880 12804
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 5160 12699 5218 12705
rect 5160 12665 5172 12699
rect 5206 12696 5218 12699
rect 5258 12696 5264 12708
rect 5206 12668 5264 12696
rect 5206 12665 5218 12668
rect 5160 12659 5218 12665
rect 5258 12656 5264 12668
rect 5316 12656 5322 12708
rect 7760 12696 7788 12727
rect 8110 12724 8116 12776
rect 8168 12764 8174 12776
rect 8389 12767 8447 12773
rect 8389 12764 8401 12767
rect 8168 12736 8401 12764
rect 8168 12724 8174 12736
rect 8389 12733 8401 12736
rect 8435 12764 8447 12767
rect 9140 12764 9168 12872
rect 10962 12860 10968 12872
rect 11020 12860 11026 12912
rect 15120 12900 15148 12940
rect 15470 12928 15476 12980
rect 15528 12928 15534 12980
rect 16577 12971 16635 12977
rect 16577 12937 16589 12971
rect 16623 12968 16635 12971
rect 16942 12968 16948 12980
rect 16623 12940 16948 12968
rect 16623 12937 16635 12940
rect 16577 12931 16635 12937
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 17310 12968 17316 12980
rect 17052 12940 17316 12968
rect 17052 12900 17080 12940
rect 17310 12928 17316 12940
rect 17368 12968 17374 12980
rect 18046 12968 18052 12980
rect 17368 12940 18052 12968
rect 17368 12928 17374 12940
rect 18046 12928 18052 12940
rect 18104 12968 18110 12980
rect 20438 12968 20444 12980
rect 18104 12940 20444 12968
rect 18104 12928 18110 12940
rect 20438 12928 20444 12940
rect 20496 12928 20502 12980
rect 22830 12928 22836 12980
rect 22888 12968 22894 12980
rect 22925 12971 22983 12977
rect 22925 12968 22937 12971
rect 22888 12940 22937 12968
rect 22888 12928 22894 12940
rect 22925 12937 22937 12940
rect 22971 12937 22983 12971
rect 22925 12931 22983 12937
rect 25222 12928 25228 12980
rect 25280 12928 25286 12980
rect 26510 12928 26516 12980
rect 26568 12968 26574 12980
rect 26697 12971 26755 12977
rect 26697 12968 26709 12971
rect 26568 12940 26709 12968
rect 26568 12928 26574 12940
rect 26697 12937 26709 12940
rect 26743 12937 26755 12971
rect 26697 12931 26755 12937
rect 15120 12872 17080 12900
rect 24394 12860 24400 12912
rect 24452 12860 24458 12912
rect 24854 12860 24860 12912
rect 24912 12900 24918 12912
rect 24912 12872 25360 12900
rect 24912 12860 24918 12872
rect 9674 12832 9680 12844
rect 9600 12804 9680 12832
rect 9600 12773 9628 12804
rect 9674 12792 9680 12804
rect 9732 12832 9738 12844
rect 9858 12832 9864 12844
rect 9732 12804 9864 12832
rect 9732 12792 9738 12804
rect 9858 12792 9864 12804
rect 9916 12832 9922 12844
rect 12066 12832 12072 12844
rect 9916 12804 12072 12832
rect 9916 12792 9922 12804
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 17954 12792 17960 12844
rect 18012 12832 18018 12844
rect 18690 12832 18696 12844
rect 18012 12804 18696 12832
rect 18012 12792 18018 12804
rect 18690 12792 18696 12804
rect 18748 12792 18754 12844
rect 21082 12792 21088 12844
rect 21140 12792 21146 12844
rect 23474 12792 23480 12844
rect 23532 12832 23538 12844
rect 24412 12832 24440 12860
rect 25038 12832 25044 12844
rect 23532 12804 23980 12832
rect 23532 12792 23538 12804
rect 8435 12736 9168 12764
rect 9585 12767 9643 12773
rect 8435 12733 8447 12736
rect 8389 12727 8447 12733
rect 9585 12733 9597 12767
rect 9631 12733 9643 12767
rect 9585 12727 9643 12733
rect 9950 12724 9956 12776
rect 10008 12724 10014 12776
rect 10134 12724 10140 12776
rect 10192 12764 10198 12776
rect 10873 12767 10931 12773
rect 10873 12764 10885 12767
rect 10192 12736 10885 12764
rect 10192 12724 10198 12736
rect 10873 12733 10885 12736
rect 10919 12764 10931 12767
rect 11974 12764 11980 12776
rect 10919 12736 11980 12764
rect 10919 12733 10931 12736
rect 10873 12727 10931 12733
rect 11974 12724 11980 12736
rect 12032 12724 12038 12776
rect 14093 12767 14151 12773
rect 14093 12733 14105 12767
rect 14139 12764 14151 12767
rect 14182 12764 14188 12776
rect 14139 12736 14188 12764
rect 14139 12733 14151 12736
rect 14093 12727 14151 12733
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 14366 12773 14372 12776
rect 14360 12764 14372 12773
rect 14327 12736 14372 12764
rect 14360 12727 14372 12736
rect 14366 12724 14372 12727
rect 14424 12724 14430 12776
rect 14826 12724 14832 12776
rect 14884 12764 14890 12776
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 14884 12736 15669 12764
rect 14884 12724 14890 12736
rect 15657 12733 15669 12736
rect 15703 12764 15715 12767
rect 16114 12764 16120 12776
rect 15703 12736 16120 12764
rect 15703 12733 15715 12736
rect 15657 12727 15715 12733
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 17126 12724 17132 12776
rect 17184 12764 17190 12776
rect 18233 12767 18291 12773
rect 18233 12764 18245 12767
rect 17184 12736 18245 12764
rect 17184 12724 17190 12736
rect 18233 12733 18245 12736
rect 18279 12733 18291 12767
rect 18233 12727 18291 12733
rect 20254 12724 20260 12776
rect 20312 12764 20318 12776
rect 23198 12764 23204 12776
rect 20312 12736 23204 12764
rect 20312 12724 20318 12736
rect 23198 12724 23204 12736
rect 23256 12764 23262 12776
rect 23952 12773 23980 12804
rect 24136 12804 24440 12832
rect 24872 12804 25044 12832
rect 24136 12773 24164 12804
rect 23845 12767 23903 12773
rect 23845 12764 23857 12767
rect 23256 12736 23857 12764
rect 23256 12724 23262 12736
rect 23845 12733 23857 12736
rect 23891 12733 23903 12767
rect 23845 12727 23903 12733
rect 23938 12767 23996 12773
rect 23938 12733 23950 12767
rect 23984 12733 23996 12767
rect 23938 12727 23996 12733
rect 24121 12767 24179 12773
rect 24121 12733 24133 12767
rect 24167 12733 24179 12767
rect 24121 12727 24179 12733
rect 24302 12724 24308 12776
rect 24360 12773 24366 12776
rect 24360 12764 24368 12773
rect 24581 12767 24639 12773
rect 24360 12736 24405 12764
rect 24360 12727 24368 12736
rect 24581 12733 24593 12767
rect 24627 12764 24639 12767
rect 24670 12764 24676 12776
rect 24627 12736 24676 12764
rect 24627 12733 24639 12736
rect 24581 12727 24639 12733
rect 24360 12724 24366 12727
rect 24670 12724 24676 12736
rect 24728 12724 24734 12776
rect 24872 12773 24900 12804
rect 25038 12792 25044 12804
rect 25096 12792 25102 12844
rect 25332 12841 25360 12872
rect 25317 12835 25375 12841
rect 25317 12801 25329 12835
rect 25363 12801 25375 12835
rect 25317 12795 25375 12801
rect 24765 12767 24823 12773
rect 24765 12733 24777 12767
rect 24811 12733 24823 12767
rect 24765 12727 24823 12733
rect 24857 12767 24915 12773
rect 24857 12733 24869 12767
rect 24903 12733 24915 12767
rect 24857 12727 24915 12733
rect 24949 12767 25007 12773
rect 24949 12733 24961 12767
rect 24995 12764 25007 12767
rect 25406 12764 25412 12776
rect 24995 12736 25412 12764
rect 24995 12733 25007 12736
rect 24949 12727 25007 12733
rect 13170 12696 13176 12708
rect 7760 12668 13176 12696
rect 3752 12600 4752 12628
rect 3752 12588 3758 12600
rect 6270 12588 6276 12640
rect 6328 12588 6334 12640
rect 8588 12637 8616 12668
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 14108 12668 15608 12696
rect 8573 12631 8631 12637
rect 8573 12597 8585 12631
rect 8619 12597 8631 12631
rect 8573 12591 8631 12597
rect 8662 12588 8668 12640
rect 8720 12628 8726 12640
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 8720 12600 9413 12628
rect 8720 12588 8726 12600
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 9401 12591 9459 12597
rect 9766 12588 9772 12640
rect 9824 12588 9830 12640
rect 10042 12588 10048 12640
rect 10100 12628 10106 12640
rect 14108 12628 14136 12668
rect 10100 12600 14136 12628
rect 15580 12628 15608 12668
rect 16942 12656 16948 12708
rect 17000 12696 17006 12708
rect 17690 12699 17748 12705
rect 17690 12696 17702 12699
rect 17000 12668 17702 12696
rect 17000 12656 17006 12668
rect 17690 12665 17702 12668
rect 17736 12665 17748 12699
rect 17690 12659 17748 12665
rect 20441 12699 20499 12705
rect 20441 12665 20453 12699
rect 20487 12696 20499 12699
rect 21634 12696 21640 12708
rect 20487 12668 21640 12696
rect 20487 12665 20499 12668
rect 20441 12659 20499 12665
rect 21634 12656 21640 12668
rect 21692 12656 21698 12708
rect 22922 12656 22928 12708
rect 22980 12696 22986 12708
rect 23382 12696 23388 12708
rect 22980 12668 23388 12696
rect 22980 12656 22986 12668
rect 23382 12656 23388 12668
rect 23440 12656 23446 12708
rect 24213 12699 24271 12705
rect 24213 12665 24225 12699
rect 24259 12696 24271 12699
rect 24780 12696 24808 12727
rect 25406 12724 25412 12736
rect 25464 12724 25470 12776
rect 25590 12705 25596 12708
rect 24259 12668 24440 12696
rect 24259 12665 24271 12668
rect 24213 12659 24271 12665
rect 24412 12640 24440 12668
rect 24504 12668 24808 12696
rect 15749 12631 15807 12637
rect 15749 12628 15761 12631
rect 15580 12600 15761 12628
rect 10100 12588 10106 12600
rect 15749 12597 15761 12600
rect 15795 12597 15807 12631
rect 15749 12591 15807 12597
rect 18417 12631 18475 12637
rect 18417 12597 18429 12631
rect 18463 12628 18475 12631
rect 19426 12628 19432 12640
rect 18463 12600 19432 12628
rect 18463 12597 18475 12600
rect 18417 12591 18475 12597
rect 19426 12588 19432 12600
rect 19484 12628 19490 12640
rect 20254 12628 20260 12640
rect 19484 12600 20260 12628
rect 19484 12588 19490 12600
rect 20254 12588 20260 12600
rect 20312 12588 20318 12640
rect 20346 12588 20352 12640
rect 20404 12628 20410 12640
rect 20533 12631 20591 12637
rect 20533 12628 20545 12631
rect 20404 12600 20545 12628
rect 20404 12588 20410 12600
rect 20533 12597 20545 12600
rect 20579 12597 20591 12631
rect 20533 12591 20591 12597
rect 23566 12588 23572 12640
rect 23624 12628 23630 12640
rect 24302 12628 24308 12640
rect 23624 12600 24308 12628
rect 23624 12588 23630 12600
rect 24302 12588 24308 12600
rect 24360 12588 24366 12640
rect 24394 12588 24400 12640
rect 24452 12588 24458 12640
rect 24504 12637 24532 12668
rect 25584 12659 25596 12705
rect 25590 12656 25596 12659
rect 25648 12656 25654 12708
rect 24489 12631 24547 12637
rect 24489 12597 24501 12631
rect 24535 12597 24547 12631
rect 24489 12591 24547 12597
rect 25038 12588 25044 12640
rect 25096 12628 25102 12640
rect 25866 12628 25872 12640
rect 25096 12600 25872 12628
rect 25096 12588 25102 12600
rect 25866 12588 25872 12600
rect 25924 12588 25930 12640
rect 552 12538 27576 12560
rect 552 12486 7114 12538
rect 7166 12486 7178 12538
rect 7230 12486 7242 12538
rect 7294 12486 7306 12538
rect 7358 12486 7370 12538
rect 7422 12486 13830 12538
rect 13882 12486 13894 12538
rect 13946 12486 13958 12538
rect 14010 12486 14022 12538
rect 14074 12486 14086 12538
rect 14138 12486 20546 12538
rect 20598 12486 20610 12538
rect 20662 12486 20674 12538
rect 20726 12486 20738 12538
rect 20790 12486 20802 12538
rect 20854 12486 27262 12538
rect 27314 12486 27326 12538
rect 27378 12486 27390 12538
rect 27442 12486 27454 12538
rect 27506 12486 27518 12538
rect 27570 12486 27576 12538
rect 552 12464 27576 12486
rect 3418 12384 3424 12436
rect 3476 12424 3482 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3476 12396 3801 12424
rect 3476 12384 3482 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 3789 12387 3847 12393
rect 5258 12384 5264 12436
rect 5316 12384 5322 12436
rect 7190 12384 7196 12436
rect 7248 12424 7254 12436
rect 8110 12424 8116 12436
rect 7248 12396 8116 12424
rect 7248 12384 7254 12396
rect 8110 12384 8116 12396
rect 8168 12384 8174 12436
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 12158 12424 12164 12436
rect 9732 12396 12164 12424
rect 9732 12384 9738 12396
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 12406 12396 12848 12424
rect 3234 12356 3240 12368
rect 2792 12328 3240 12356
rect 2593 12291 2651 12297
rect 2593 12257 2605 12291
rect 2639 12257 2651 12291
rect 2593 12251 2651 12257
rect 2608 12220 2636 12251
rect 2682 12248 2688 12300
rect 2740 12248 2746 12300
rect 2792 12297 2820 12328
rect 3234 12316 3240 12328
rect 3292 12316 3298 12368
rect 5626 12356 5632 12368
rect 4264 12328 5632 12356
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12257 2835 12291
rect 2777 12251 2835 12257
rect 2961 12291 3019 12297
rect 2961 12257 2973 12291
rect 3007 12288 3019 12291
rect 3510 12288 3516 12300
rect 3007 12260 3516 12288
rect 3007 12257 3019 12260
rect 2961 12251 3019 12257
rect 3510 12248 3516 12260
rect 3568 12248 3574 12300
rect 4264 12297 4292 12328
rect 5626 12316 5632 12328
rect 5684 12356 5690 12368
rect 6270 12356 6276 12368
rect 5684 12328 6276 12356
rect 5684 12316 5690 12328
rect 6270 12316 6276 12328
rect 6328 12316 6334 12368
rect 7009 12359 7067 12365
rect 7009 12325 7021 12359
rect 7055 12356 7067 12359
rect 8662 12356 8668 12368
rect 7055 12328 8668 12356
rect 7055 12325 7067 12328
rect 7009 12319 7067 12325
rect 8662 12316 8668 12328
rect 8720 12316 8726 12368
rect 9769 12359 9827 12365
rect 9769 12356 9781 12359
rect 9140 12328 9781 12356
rect 4249 12291 4307 12297
rect 4249 12257 4261 12291
rect 4295 12257 4307 12291
rect 4249 12251 4307 12257
rect 4982 12248 4988 12300
rect 5040 12248 5046 12300
rect 5169 12291 5227 12297
rect 5169 12257 5181 12291
rect 5215 12288 5227 12291
rect 5445 12291 5503 12297
rect 5445 12288 5457 12291
rect 5215 12260 5457 12288
rect 5215 12257 5227 12260
rect 5169 12251 5227 12257
rect 5445 12257 5457 12260
rect 5491 12257 5503 12291
rect 5445 12251 5503 12257
rect 7190 12248 7196 12300
rect 7248 12248 7254 12300
rect 7466 12248 7472 12300
rect 7524 12248 7530 12300
rect 7745 12291 7803 12297
rect 7745 12257 7757 12291
rect 7791 12257 7803 12291
rect 7745 12251 7803 12257
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 3053 12223 3111 12229
rect 3053 12220 3065 12223
rect 2608 12192 3065 12220
rect 3053 12189 3065 12192
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 3602 12180 3608 12232
rect 3660 12180 3666 12232
rect 4798 12180 4804 12232
rect 4856 12180 4862 12232
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12220 6883 12223
rect 7760 12220 7788 12251
rect 6871 12192 7788 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 6638 12112 6644 12164
rect 6696 12152 6702 12164
rect 6696 12124 7512 12152
rect 6696 12112 6702 12124
rect 2314 12044 2320 12096
rect 2372 12044 2378 12096
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 3973 12087 4031 12093
rect 3973 12084 3985 12087
rect 3660 12056 3985 12084
rect 3660 12044 3666 12056
rect 3973 12053 3985 12056
rect 4019 12053 4031 12087
rect 3973 12047 4031 12053
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 7285 12087 7343 12093
rect 7285 12084 7297 12087
rect 6972 12056 7297 12084
rect 6972 12044 6978 12056
rect 7285 12053 7297 12056
rect 7331 12053 7343 12087
rect 7484 12084 7512 12124
rect 7558 12112 7564 12164
rect 7616 12112 7622 12164
rect 7650 12112 7656 12164
rect 7708 12112 7714 12164
rect 7944 12084 7972 12251
rect 8938 12248 8944 12300
rect 8996 12248 9002 12300
rect 9140 12297 9168 12328
rect 9769 12325 9781 12328
rect 9815 12325 9827 12359
rect 12406 12356 12434 12396
rect 9769 12319 9827 12325
rect 11164 12328 12434 12356
rect 9125 12291 9183 12297
rect 9125 12257 9137 12291
rect 9171 12257 9183 12291
rect 9125 12251 9183 12257
rect 9398 12248 9404 12300
rect 9456 12288 9462 12300
rect 9493 12291 9551 12297
rect 9493 12288 9505 12291
rect 9456 12260 9505 12288
rect 9456 12248 9462 12260
rect 9493 12257 9505 12260
rect 9539 12257 9551 12291
rect 9493 12251 9551 12257
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 11164 12297 11192 12328
rect 9953 12291 10011 12297
rect 9953 12288 9965 12291
rect 9916 12260 9965 12288
rect 9916 12248 9922 12260
rect 9953 12257 9965 12260
rect 9999 12257 10011 12291
rect 10229 12291 10287 12297
rect 10229 12288 10241 12291
rect 9953 12251 10011 12257
rect 10060 12260 10241 12288
rect 8018 12180 8024 12232
rect 8076 12180 8082 12232
rect 9214 12180 9220 12232
rect 9272 12180 9278 12232
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12220 9367 12223
rect 9582 12220 9588 12232
rect 9355 12192 9588 12220
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 9582 12180 9588 12192
rect 9640 12220 9646 12232
rect 10060 12220 10088 12260
rect 10229 12257 10241 12260
rect 10275 12288 10287 12291
rect 10965 12291 11023 12297
rect 10965 12288 10977 12291
rect 10275 12260 10977 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 10965 12257 10977 12260
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12257 11207 12291
rect 11149 12251 11207 12257
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12288 11483 12291
rect 11514 12288 11520 12300
rect 11471 12260 11520 12288
rect 11471 12257 11483 12260
rect 11425 12251 11483 12257
rect 9640 12192 10088 12220
rect 9640 12180 9646 12192
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 11164 12220 11192 12251
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 11692 12291 11750 12297
rect 11692 12257 11704 12291
rect 11738 12288 11750 12291
rect 12066 12288 12072 12300
rect 11738 12260 12072 12288
rect 11738 12257 11750 12260
rect 11692 12251 11750 12257
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 10192 12192 11192 12220
rect 10192 12180 10198 12192
rect 8754 12112 8760 12164
rect 8812 12152 8818 12164
rect 10413 12155 10471 12161
rect 10413 12152 10425 12155
rect 8812 12124 10425 12152
rect 8812 12112 8818 12124
rect 10413 12121 10425 12124
rect 10459 12121 10471 12155
rect 10413 12115 10471 12121
rect 7484 12056 7972 12084
rect 7285 12047 7343 12053
rect 9674 12044 9680 12096
rect 9732 12044 9738 12096
rect 11333 12087 11391 12093
rect 11333 12053 11345 12087
rect 11379 12084 11391 12087
rect 11606 12084 11612 12096
rect 11379 12056 11612 12084
rect 11379 12053 11391 12056
rect 11333 12047 11391 12053
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 12158 12044 12164 12096
rect 12216 12084 12222 12096
rect 12710 12084 12716 12096
rect 12216 12056 12716 12084
rect 12216 12044 12222 12056
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 12820 12093 12848 12396
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 14274 12424 14280 12436
rect 13872 12396 14280 12424
rect 13872 12384 13878 12396
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 14737 12427 14795 12433
rect 14737 12393 14749 12427
rect 14783 12393 14795 12427
rect 14737 12387 14795 12393
rect 14182 12356 14188 12368
rect 13372 12328 14188 12356
rect 13372 12297 13400 12328
rect 14182 12316 14188 12328
rect 14240 12316 14246 12368
rect 14752 12356 14780 12387
rect 16206 12384 16212 12436
rect 16264 12384 16270 12436
rect 16942 12384 16948 12436
rect 17000 12384 17006 12436
rect 17586 12424 17592 12436
rect 17144 12396 17592 12424
rect 16666 12356 16672 12368
rect 14752 12328 16672 12356
rect 13630 12297 13636 12300
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12257 13415 12291
rect 13624 12288 13636 12297
rect 13591 12260 13636 12288
rect 13357 12251 13415 12257
rect 13624 12251 13636 12260
rect 13630 12248 13636 12251
rect 13688 12248 13694 12300
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 15488 12297 15516 12328
rect 16666 12316 16672 12328
rect 16724 12316 16730 12368
rect 14829 12291 14887 12297
rect 14829 12288 14841 12291
rect 13964 12260 14841 12288
rect 13964 12248 13970 12260
rect 14829 12257 14841 12260
rect 14875 12257 14887 12291
rect 14829 12251 14887 12257
rect 15473 12291 15531 12297
rect 15473 12257 15485 12291
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 14458 12180 14464 12232
rect 14516 12220 14522 12232
rect 14918 12220 14924 12232
rect 14516 12192 14924 12220
rect 14516 12180 14522 12192
rect 14918 12180 14924 12192
rect 14976 12220 14982 12232
rect 15672 12220 15700 12251
rect 15930 12248 15936 12300
rect 15988 12248 15994 12300
rect 16117 12291 16175 12297
rect 16117 12257 16129 12291
rect 16163 12257 16175 12291
rect 16117 12251 16175 12257
rect 16301 12291 16359 12297
rect 16301 12257 16313 12291
rect 16347 12257 16359 12291
rect 17144 12288 17172 12396
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 19978 12384 19984 12436
rect 20036 12424 20042 12436
rect 20073 12427 20131 12433
rect 20073 12424 20085 12427
rect 20036 12396 20085 12424
rect 20036 12384 20042 12396
rect 20073 12393 20085 12396
rect 20119 12393 20131 12427
rect 20073 12387 20131 12393
rect 22738 12384 22744 12436
rect 22796 12384 22802 12436
rect 25038 12424 25044 12436
rect 23308 12396 25044 12424
rect 18868 12359 18926 12365
rect 18868 12325 18880 12359
rect 18914 12356 18926 12359
rect 18966 12356 18972 12368
rect 18914 12328 18972 12356
rect 18914 12325 18926 12328
rect 18868 12319 18926 12325
rect 18966 12316 18972 12328
rect 19024 12316 19030 12368
rect 19794 12316 19800 12368
rect 19852 12356 19858 12368
rect 19852 12328 20484 12356
rect 19852 12316 19858 12328
rect 19996 12300 20024 12328
rect 17221 12291 17279 12297
rect 17221 12288 17233 12291
rect 17144 12260 17233 12288
rect 16301 12251 16359 12257
rect 17221 12257 17233 12260
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 16132 12220 16160 12251
rect 14976 12192 15700 12220
rect 15856 12192 16160 12220
rect 16316 12220 16344 12251
rect 17310 12248 17316 12300
rect 17368 12248 17374 12300
rect 17405 12291 17463 12297
rect 17405 12257 17417 12291
rect 17451 12257 17463 12291
rect 17405 12251 17463 12257
rect 17589 12291 17647 12297
rect 17589 12257 17601 12291
rect 17635 12288 17647 12291
rect 18322 12288 18328 12300
rect 17635 12260 18328 12288
rect 17635 12257 17647 12260
rect 17589 12251 17647 12257
rect 17328 12220 17356 12248
rect 16316 12192 17356 12220
rect 14976 12180 14982 12192
rect 15856 12096 15884 12192
rect 17420 12152 17448 12251
rect 18322 12248 18328 12260
rect 18380 12248 18386 12300
rect 18601 12291 18659 12297
rect 18601 12257 18613 12291
rect 18647 12288 18659 12291
rect 18690 12288 18696 12300
rect 18647 12260 18696 12288
rect 18647 12257 18659 12260
rect 18601 12251 18659 12257
rect 18690 12248 18696 12260
rect 18748 12248 18754 12300
rect 19978 12248 19984 12300
rect 20036 12248 20042 12300
rect 20346 12248 20352 12300
rect 20404 12248 20410 12300
rect 20456 12297 20484 12328
rect 21726 12316 21732 12368
rect 21784 12356 21790 12368
rect 23308 12356 23336 12396
rect 25038 12384 25044 12396
rect 25096 12384 25102 12436
rect 25501 12427 25559 12433
rect 25501 12393 25513 12427
rect 25547 12424 25559 12427
rect 25590 12424 25596 12436
rect 25547 12396 25596 12424
rect 25547 12393 25559 12396
rect 25501 12387 25559 12393
rect 25590 12384 25596 12396
rect 25648 12384 25654 12436
rect 25958 12424 25964 12436
rect 25700 12396 25964 12424
rect 21784 12328 22324 12356
rect 21784 12316 21790 12328
rect 20441 12291 20499 12297
rect 20441 12257 20453 12291
rect 20487 12257 20499 12291
rect 20441 12251 20499 12257
rect 20530 12248 20536 12300
rect 20588 12248 20594 12300
rect 22296 12297 22324 12328
rect 22388 12328 23336 12356
rect 22388 12297 22416 12328
rect 23382 12316 23388 12368
rect 23440 12356 23446 12368
rect 23440 12328 23612 12356
rect 23440 12316 23446 12328
rect 20717 12291 20775 12297
rect 20717 12257 20729 12291
rect 20763 12288 20775 12291
rect 22097 12291 22155 12297
rect 22097 12288 22109 12291
rect 20763 12260 22109 12288
rect 20763 12257 20775 12260
rect 20717 12251 20775 12257
rect 22097 12257 22109 12260
rect 22143 12257 22155 12291
rect 22097 12251 22155 12257
rect 22281 12291 22339 12297
rect 22281 12257 22293 12291
rect 22327 12257 22339 12291
rect 22281 12251 22339 12257
rect 22373 12291 22431 12297
rect 22373 12257 22385 12291
rect 22419 12257 22431 12291
rect 22373 12251 22431 12257
rect 22465 12291 22523 12297
rect 22465 12257 22477 12291
rect 22511 12288 22523 12291
rect 22833 12291 22891 12297
rect 22833 12288 22845 12291
rect 22511 12260 22845 12288
rect 22511 12257 22523 12260
rect 22465 12251 22523 12257
rect 22833 12257 22845 12260
rect 22879 12257 22891 12291
rect 22833 12251 22891 12257
rect 21266 12180 21272 12232
rect 21324 12220 21330 12232
rect 21913 12223 21971 12229
rect 21913 12220 21925 12223
rect 21324 12192 21925 12220
rect 21324 12180 21330 12192
rect 21913 12189 21925 12192
rect 21959 12189 21971 12223
rect 21913 12183 21971 12189
rect 17586 12152 17592 12164
rect 17420 12124 17592 12152
rect 17586 12112 17592 12124
rect 17644 12112 17650 12164
rect 19981 12155 20039 12161
rect 19981 12121 19993 12155
rect 20027 12152 20039 12155
rect 20070 12152 20076 12164
rect 20027 12124 20076 12152
rect 20027 12121 20039 12124
rect 19981 12115 20039 12121
rect 20070 12112 20076 12124
rect 20128 12112 20134 12164
rect 22112 12152 22140 12251
rect 23474 12248 23480 12300
rect 23532 12248 23538 12300
rect 23584 12297 23612 12328
rect 23953 12328 25084 12356
rect 23569 12291 23627 12297
rect 23569 12257 23581 12291
rect 23615 12257 23627 12291
rect 23569 12251 23627 12257
rect 23474 12152 23480 12164
rect 22112 12124 23480 12152
rect 23474 12112 23480 12124
rect 23532 12112 23538 12164
rect 23753 12155 23811 12161
rect 23753 12121 23765 12155
rect 23799 12152 23811 12155
rect 23953 12152 23981 12328
rect 25056 12300 25084 12328
rect 24302 12248 24308 12300
rect 24360 12288 24366 12300
rect 24765 12291 24823 12297
rect 24765 12288 24777 12291
rect 24360 12260 24777 12288
rect 24360 12248 24366 12260
rect 24765 12257 24777 12260
rect 24811 12257 24823 12291
rect 24765 12251 24823 12257
rect 24949 12291 25007 12297
rect 24949 12257 24961 12291
rect 24995 12257 25007 12291
rect 24949 12251 25007 12257
rect 23799 12124 23981 12152
rect 23799 12121 23811 12124
rect 23753 12115 23811 12121
rect 24762 12112 24768 12164
rect 24820 12152 24826 12164
rect 24964 12152 24992 12251
rect 25038 12248 25044 12300
rect 25096 12248 25102 12300
rect 25133 12291 25191 12297
rect 25133 12257 25145 12291
rect 25179 12288 25191 12291
rect 25700 12288 25728 12396
rect 25958 12384 25964 12396
rect 26016 12424 26022 12436
rect 26421 12427 26479 12433
rect 26421 12424 26433 12427
rect 26016 12396 26433 12424
rect 26016 12384 26022 12396
rect 26421 12393 26433 12396
rect 26467 12393 26479 12427
rect 26421 12387 26479 12393
rect 26234 12356 26240 12368
rect 25976 12328 26240 12356
rect 25179 12260 25728 12288
rect 25179 12257 25191 12260
rect 25133 12251 25191 12257
rect 25774 12248 25780 12300
rect 25832 12248 25838 12300
rect 25866 12248 25872 12300
rect 25924 12248 25930 12300
rect 25976 12297 26004 12328
rect 26234 12316 26240 12328
rect 26292 12316 26298 12368
rect 25961 12291 26019 12297
rect 25961 12257 25973 12291
rect 26007 12257 26019 12291
rect 25961 12251 26019 12257
rect 26145 12291 26203 12297
rect 26145 12257 26157 12291
rect 26191 12257 26203 12291
rect 26145 12251 26203 12257
rect 26160 12152 26188 12251
rect 26234 12180 26240 12232
rect 26292 12220 26298 12232
rect 26973 12223 27031 12229
rect 26973 12220 26985 12223
rect 26292 12192 26985 12220
rect 26292 12180 26298 12192
rect 26973 12189 26985 12192
rect 27019 12189 27031 12223
rect 26973 12183 27031 12189
rect 24820 12124 24992 12152
rect 25056 12124 26188 12152
rect 24820 12112 24826 12124
rect 12805 12087 12863 12093
rect 12805 12053 12817 12087
rect 12851 12084 12863 12087
rect 15010 12084 15016 12096
rect 12851 12056 15016 12084
rect 12851 12053 12863 12056
rect 12805 12047 12863 12053
rect 15010 12044 15016 12056
rect 15068 12044 15074 12096
rect 15838 12044 15844 12096
rect 15896 12044 15902 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 18966 12084 18972 12096
rect 16080 12056 18972 12084
rect 16080 12044 16086 12056
rect 18966 12044 18972 12056
rect 19024 12044 19030 12096
rect 21358 12044 21364 12096
rect 21416 12044 21422 12096
rect 24670 12044 24676 12096
rect 24728 12084 24734 12096
rect 25056 12084 25084 12124
rect 24728 12056 25084 12084
rect 24728 12044 24734 12056
rect 25406 12044 25412 12096
rect 25464 12044 25470 12096
rect 552 11994 27416 12016
rect 552 11942 3756 11994
rect 3808 11942 3820 11994
rect 3872 11942 3884 11994
rect 3936 11942 3948 11994
rect 4000 11942 4012 11994
rect 4064 11942 10472 11994
rect 10524 11942 10536 11994
rect 10588 11942 10600 11994
rect 10652 11942 10664 11994
rect 10716 11942 10728 11994
rect 10780 11942 17188 11994
rect 17240 11942 17252 11994
rect 17304 11942 17316 11994
rect 17368 11942 17380 11994
rect 17432 11942 17444 11994
rect 17496 11942 23904 11994
rect 23956 11942 23968 11994
rect 24020 11942 24032 11994
rect 24084 11942 24096 11994
rect 24148 11942 24160 11994
rect 24212 11942 27416 11994
rect 552 11920 27416 11942
rect 3053 11883 3111 11889
rect 3053 11849 3065 11883
rect 3099 11880 3111 11883
rect 3602 11880 3608 11892
rect 3099 11852 3608 11880
rect 3099 11849 3111 11852
rect 3053 11843 3111 11849
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 7834 11880 7840 11892
rect 7616 11852 7840 11880
rect 7616 11840 7622 11852
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 8941 11883 8999 11889
rect 8941 11849 8953 11883
rect 8987 11880 8999 11883
rect 9214 11880 9220 11892
rect 8987 11852 9220 11880
rect 8987 11849 8999 11852
rect 8941 11843 8999 11849
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 12066 11840 12072 11892
rect 12124 11840 12130 11892
rect 13357 11883 13415 11889
rect 13357 11849 13369 11883
rect 13403 11880 13415 11883
rect 13814 11880 13820 11892
rect 13403 11852 13820 11880
rect 13403 11849 13415 11852
rect 13357 11843 13415 11849
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 14642 11840 14648 11892
rect 14700 11880 14706 11892
rect 15105 11883 15163 11889
rect 14700 11852 14964 11880
rect 14700 11840 14706 11852
rect 4798 11772 4804 11824
rect 4856 11812 4862 11824
rect 12434 11812 12440 11824
rect 4856 11784 12440 11812
rect 4856 11772 4862 11784
rect 12434 11772 12440 11784
rect 12492 11772 12498 11824
rect 12710 11772 12716 11824
rect 12768 11812 12774 11824
rect 14936 11812 14964 11852
rect 15105 11849 15117 11883
rect 15151 11880 15163 11883
rect 15562 11880 15568 11892
rect 15151 11852 15568 11880
rect 15151 11849 15163 11852
rect 15105 11843 15163 11849
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 17405 11883 17463 11889
rect 17405 11849 17417 11883
rect 17451 11880 17463 11883
rect 17586 11880 17592 11892
rect 17451 11852 17592 11880
rect 17451 11849 17463 11852
rect 17405 11843 17463 11849
rect 17586 11840 17592 11852
rect 17644 11840 17650 11892
rect 18138 11840 18144 11892
rect 18196 11880 18202 11892
rect 18233 11883 18291 11889
rect 18233 11880 18245 11883
rect 18196 11852 18245 11880
rect 18196 11840 18202 11852
rect 18233 11849 18245 11852
rect 18279 11849 18291 11883
rect 18233 11843 18291 11849
rect 19337 11883 19395 11889
rect 19337 11849 19349 11883
rect 19383 11880 19395 11883
rect 19886 11880 19892 11892
rect 19383 11852 19892 11880
rect 19383 11849 19395 11852
rect 19337 11843 19395 11849
rect 19886 11840 19892 11852
rect 19944 11840 19950 11892
rect 20073 11883 20131 11889
rect 20073 11849 20085 11883
rect 20119 11880 20131 11883
rect 20530 11880 20536 11892
rect 20119 11852 20536 11880
rect 20119 11849 20131 11852
rect 20073 11843 20131 11849
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 21450 11840 21456 11892
rect 21508 11880 21514 11892
rect 22557 11883 22615 11889
rect 22557 11880 22569 11883
rect 21508 11852 22569 11880
rect 21508 11840 21514 11852
rect 22557 11849 22569 11852
rect 22603 11849 22615 11883
rect 22557 11843 22615 11849
rect 23474 11840 23480 11892
rect 23532 11880 23538 11892
rect 24670 11880 24676 11892
rect 23532 11852 24676 11880
rect 23532 11840 23538 11852
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 26234 11840 26240 11892
rect 26292 11840 26298 11892
rect 15197 11815 15255 11821
rect 15197 11812 15209 11815
rect 12768 11784 14688 11812
rect 14936 11784 15209 11812
rect 12768 11772 12774 11784
rect 9950 11744 9956 11756
rect 8404 11716 9956 11744
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11676 1731 11679
rect 2406 11676 2412 11688
rect 1719 11648 2412 11676
rect 1719 11645 1731 11648
rect 1673 11639 1731 11645
rect 2406 11636 2412 11648
rect 2464 11636 2470 11688
rect 8404 11685 8432 11716
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 11333 11747 11391 11753
rect 11333 11713 11345 11747
rect 11379 11744 11391 11747
rect 11514 11744 11520 11756
rect 11379 11716 11520 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 13170 11744 13176 11756
rect 13004 11716 13176 11744
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11645 8447 11679
rect 8389 11639 8447 11645
rect 8478 11636 8484 11688
rect 8536 11636 8542 11688
rect 8662 11636 8668 11688
rect 8720 11636 8726 11688
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 8846 11676 8852 11688
rect 8803 11648 8852 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 8846 11636 8852 11648
rect 8904 11636 8910 11688
rect 9306 11636 9312 11688
rect 9364 11676 9370 11688
rect 11425 11679 11483 11685
rect 11425 11676 11437 11679
rect 9364 11648 11437 11676
rect 9364 11636 9370 11648
rect 11425 11645 11437 11648
rect 11471 11645 11483 11679
rect 11425 11639 11483 11645
rect 11606 11636 11612 11688
rect 11664 11636 11670 11688
rect 11698 11636 11704 11688
rect 11756 11636 11762 11688
rect 11793 11679 11851 11685
rect 11793 11645 11805 11679
rect 11839 11676 11851 11679
rect 12158 11676 12164 11688
rect 11839 11648 12164 11676
rect 11839 11645 11851 11648
rect 11793 11639 11851 11645
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 13004 11685 13032 11716
rect 13170 11704 13176 11716
rect 13228 11704 13234 11756
rect 13722 11704 13728 11756
rect 13780 11744 13786 11756
rect 14090 11744 14096 11756
rect 13780 11716 14096 11744
rect 13780 11704 13786 11716
rect 14090 11704 14096 11716
rect 14148 11704 14154 11756
rect 14366 11704 14372 11756
rect 14424 11744 14430 11756
rect 14461 11747 14519 11753
rect 14461 11744 14473 11747
rect 14424 11716 14473 11744
rect 14424 11704 14430 11716
rect 14461 11713 14473 11716
rect 14507 11713 14519 11747
rect 14660 11744 14688 11784
rect 15197 11781 15209 11784
rect 15243 11781 15255 11815
rect 15197 11775 15255 11781
rect 15304 11784 18736 11812
rect 15304 11744 15332 11784
rect 14660 11716 15332 11744
rect 15749 11747 15807 11753
rect 14461 11707 14519 11713
rect 15749 11713 15761 11747
rect 15795 11744 15807 11747
rect 15795 11716 16528 11744
rect 15795 11713 15807 11716
rect 15749 11707 15807 11713
rect 12713 11679 12771 11685
rect 12713 11676 12725 11679
rect 12360 11648 12725 11676
rect 1940 11611 1998 11617
rect 1940 11577 1952 11611
rect 1986 11608 1998 11611
rect 2314 11608 2320 11620
rect 1986 11580 2320 11608
rect 1986 11577 1998 11580
rect 1940 11571 1998 11577
rect 2314 11568 2320 11580
rect 2372 11568 2378 11620
rect 5810 11568 5816 11620
rect 5868 11608 5874 11620
rect 6086 11608 6092 11620
rect 5868 11580 6092 11608
rect 5868 11568 5874 11580
rect 6086 11568 6092 11580
rect 6144 11608 6150 11620
rect 6273 11611 6331 11617
rect 6273 11608 6285 11611
rect 6144 11580 6285 11608
rect 6144 11568 6150 11580
rect 6273 11577 6285 11580
rect 6319 11577 6331 11611
rect 6273 11571 6331 11577
rect 8021 11611 8079 11617
rect 8021 11577 8033 11611
rect 8067 11608 8079 11611
rect 9582 11608 9588 11620
rect 8067 11580 9588 11608
rect 8067 11577 8079 11580
rect 8021 11571 8079 11577
rect 9582 11568 9588 11580
rect 9640 11568 9646 11620
rect 12066 11568 12072 11620
rect 12124 11608 12130 11620
rect 12253 11611 12311 11617
rect 12253 11608 12265 11611
rect 12124 11580 12265 11608
rect 12124 11568 12130 11580
rect 12253 11577 12265 11580
rect 12299 11577 12311 11611
rect 12253 11571 12311 11577
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 8938 11540 8944 11552
rect 4856 11512 8944 11540
rect 4856 11500 4862 11512
rect 8938 11500 8944 11512
rect 8996 11540 9002 11552
rect 9950 11540 9956 11552
rect 8996 11512 9956 11540
rect 8996 11500 9002 11512
rect 9950 11500 9956 11512
rect 10008 11540 10014 11552
rect 12360 11540 12388 11648
rect 12713 11645 12725 11648
rect 12759 11645 12771 11679
rect 12713 11639 12771 11645
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 12989 11679 13047 11685
rect 12989 11645 13001 11679
rect 13035 11645 13047 11679
rect 12989 11639 13047 11645
rect 13081 11679 13139 11685
rect 13081 11645 13093 11679
rect 13127 11676 13139 11679
rect 13906 11676 13912 11688
rect 13127 11648 13912 11676
rect 13127 11645 13139 11648
rect 13081 11639 13139 11645
rect 12434 11568 12440 11620
rect 12492 11608 12498 11620
rect 12802 11608 12808 11620
rect 12492 11580 12808 11608
rect 12492 11568 12498 11580
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 12912 11608 12940 11639
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 14476 11676 14504 11707
rect 15764 11676 15792 11707
rect 14476 11648 15792 11676
rect 16114 11636 16120 11688
rect 16172 11676 16178 11688
rect 16500 11685 16528 11716
rect 17236 11716 18092 11744
rect 16209 11679 16267 11685
rect 16209 11676 16221 11679
rect 16172 11648 16221 11676
rect 16172 11636 16178 11648
rect 16209 11645 16221 11648
rect 16255 11645 16267 11679
rect 16209 11639 16267 11645
rect 16485 11679 16543 11685
rect 16485 11645 16497 11679
rect 16531 11676 16543 11679
rect 16945 11679 17003 11685
rect 16945 11676 16957 11679
rect 16531 11648 16957 11676
rect 16531 11645 16543 11648
rect 16485 11639 16543 11645
rect 16945 11645 16957 11648
rect 16991 11676 17003 11679
rect 17126 11676 17132 11688
rect 16991 11648 17132 11676
rect 16991 11645 17003 11648
rect 16945 11639 17003 11645
rect 16025 11611 16083 11617
rect 16025 11608 16037 11611
rect 12912 11580 16037 11608
rect 16025 11577 16037 11580
rect 16071 11577 16083 11611
rect 16224 11608 16252 11639
rect 17126 11636 17132 11648
rect 17184 11636 17190 11688
rect 17236 11685 17264 11716
rect 18064 11688 18092 11716
rect 17221 11679 17279 11685
rect 17221 11645 17233 11679
rect 17267 11645 17279 11679
rect 17763 11657 17821 11663
rect 17763 11654 17775 11657
rect 17221 11639 17279 11645
rect 17236 11608 17264 11639
rect 16224 11580 17264 11608
rect 17705 11626 17775 11654
rect 16025 11571 16083 11577
rect 10008 11512 12388 11540
rect 10008 11500 10014 11512
rect 12618 11500 12624 11552
rect 12676 11540 12682 11552
rect 13541 11543 13599 11549
rect 13541 11540 13553 11543
rect 12676 11512 13553 11540
rect 12676 11500 12682 11512
rect 13541 11509 13553 11512
rect 13587 11509 13599 11543
rect 13541 11503 13599 11509
rect 14642 11500 14648 11552
rect 14700 11500 14706 11552
rect 14737 11543 14795 11549
rect 14737 11509 14749 11543
rect 14783 11540 14795 11543
rect 15010 11540 15016 11552
rect 14783 11512 15016 11540
rect 14783 11509 14795 11512
rect 14737 11503 14795 11509
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 15562 11500 15568 11552
rect 15620 11500 15626 11552
rect 15654 11500 15660 11552
rect 15712 11500 15718 11552
rect 16393 11543 16451 11549
rect 16393 11509 16405 11543
rect 16439 11540 16451 11543
rect 16942 11540 16948 11552
rect 16439 11512 16948 11540
rect 16439 11509 16451 11512
rect 16393 11503 16451 11509
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17034 11500 17040 11552
rect 17092 11500 17098 11552
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 17705 11540 17733 11626
rect 17763 11623 17775 11626
rect 17809 11623 17821 11657
rect 18046 11636 18052 11688
rect 18104 11636 18110 11688
rect 18708 11685 18736 11784
rect 18966 11772 18972 11824
rect 19024 11812 19030 11824
rect 22465 11815 22523 11821
rect 19024 11784 19334 11812
rect 19024 11772 19030 11784
rect 18693 11679 18751 11685
rect 18693 11645 18705 11679
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 18782 11636 18788 11688
rect 18840 11636 18846 11688
rect 18984 11685 19012 11772
rect 19306 11744 19334 11784
rect 22465 11781 22477 11815
rect 22511 11812 22523 11815
rect 22511 11784 23152 11812
rect 22511 11781 22523 11784
rect 22465 11775 22523 11781
rect 23124 11753 23152 11784
rect 23109 11747 23167 11753
rect 19306 11716 19656 11744
rect 18969 11679 19027 11685
rect 18969 11645 18981 11679
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 19199 11679 19257 11685
rect 19199 11645 19211 11679
rect 19245 11676 19257 11679
rect 19334 11676 19340 11688
rect 19245 11648 19340 11676
rect 19245 11645 19257 11648
rect 19199 11639 19257 11645
rect 19334 11636 19340 11648
rect 19392 11636 19398 11688
rect 19426 11636 19432 11688
rect 19484 11636 19490 11688
rect 19518 11636 19524 11688
rect 19576 11636 19582 11688
rect 17763 11617 17821 11623
rect 19061 11611 19119 11617
rect 19061 11577 19073 11611
rect 19107 11577 19119 11611
rect 19628 11608 19656 11716
rect 23109 11713 23121 11747
rect 23155 11713 23167 11747
rect 23109 11707 23167 11713
rect 24394 11704 24400 11756
rect 24452 11704 24458 11756
rect 24854 11704 24860 11756
rect 24912 11704 24918 11756
rect 19886 11636 19892 11688
rect 19944 11685 19950 11688
rect 19944 11676 19952 11685
rect 20438 11676 20444 11688
rect 19944 11648 20444 11676
rect 19944 11639 19952 11648
rect 19944 11636 19950 11639
rect 20438 11636 20444 11648
rect 20496 11636 20502 11688
rect 21085 11679 21143 11685
rect 21085 11645 21097 11679
rect 21131 11676 21143 11679
rect 21174 11676 21180 11688
rect 21131 11648 21180 11676
rect 21131 11645 21143 11648
rect 21085 11639 21143 11645
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 22830 11636 22836 11688
rect 22888 11676 22894 11688
rect 23293 11679 23351 11685
rect 23293 11676 23305 11679
rect 22888 11648 23305 11676
rect 22888 11636 22894 11648
rect 23293 11645 23305 11648
rect 23339 11645 23351 11679
rect 23293 11639 23351 11645
rect 25124 11679 25182 11685
rect 25124 11645 25136 11679
rect 25170 11676 25182 11679
rect 25406 11676 25412 11688
rect 25170 11648 25412 11676
rect 25170 11645 25182 11648
rect 25124 11639 25182 11645
rect 25406 11636 25412 11648
rect 25464 11636 25470 11688
rect 26234 11636 26240 11688
rect 26292 11676 26298 11688
rect 26694 11676 26700 11688
rect 26292 11648 26700 11676
rect 26292 11636 26298 11648
rect 26694 11636 26700 11648
rect 26752 11676 26758 11688
rect 26881 11679 26939 11685
rect 26881 11676 26893 11679
rect 26752 11648 26893 11676
rect 26752 11636 26758 11648
rect 26881 11645 26893 11648
rect 26927 11645 26939 11679
rect 26881 11639 26939 11645
rect 19705 11611 19763 11617
rect 19705 11608 19717 11611
rect 19628 11580 19717 11608
rect 19061 11571 19119 11577
rect 19705 11577 19717 11580
rect 19751 11577 19763 11611
rect 19705 11571 19763 11577
rect 17184 11512 17733 11540
rect 17865 11543 17923 11549
rect 17184 11500 17190 11512
rect 17865 11509 17877 11543
rect 17911 11540 17923 11543
rect 18966 11540 18972 11552
rect 17911 11512 18972 11540
rect 17911 11509 17923 11512
rect 17865 11503 17923 11509
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 19076 11540 19104 11571
rect 19794 11568 19800 11620
rect 19852 11568 19858 11620
rect 21358 11617 21364 11620
rect 21352 11608 21364 11617
rect 21319 11580 21364 11608
rect 21352 11571 21364 11580
rect 21358 11568 21364 11571
rect 21416 11568 21422 11620
rect 20254 11540 20260 11552
rect 19076 11512 20260 11540
rect 20254 11500 20260 11512
rect 20312 11500 20318 11552
rect 23658 11500 23664 11552
rect 23716 11540 23722 11552
rect 23845 11543 23903 11549
rect 23845 11540 23857 11543
rect 23716 11512 23857 11540
rect 23716 11500 23722 11512
rect 23845 11509 23857 11512
rect 23891 11509 23903 11543
rect 23845 11503 23903 11509
rect 25130 11500 25136 11552
rect 25188 11540 25194 11552
rect 26329 11543 26387 11549
rect 26329 11540 26341 11543
rect 25188 11512 26341 11540
rect 25188 11500 25194 11512
rect 26329 11509 26341 11512
rect 26375 11509 26387 11543
rect 26329 11503 26387 11509
rect 552 11450 27576 11472
rect 552 11398 7114 11450
rect 7166 11398 7178 11450
rect 7230 11398 7242 11450
rect 7294 11398 7306 11450
rect 7358 11398 7370 11450
rect 7422 11398 13830 11450
rect 13882 11398 13894 11450
rect 13946 11398 13958 11450
rect 14010 11398 14022 11450
rect 14074 11398 14086 11450
rect 14138 11398 20546 11450
rect 20598 11398 20610 11450
rect 20662 11398 20674 11450
rect 20726 11398 20738 11450
rect 20790 11398 20802 11450
rect 20854 11398 27262 11450
rect 27314 11398 27326 11450
rect 27378 11398 27390 11450
rect 27442 11398 27454 11450
rect 27506 11398 27518 11450
rect 27570 11398 27576 11450
rect 552 11376 27576 11398
rect 3510 11296 3516 11348
rect 3568 11336 3574 11348
rect 7193 11339 7251 11345
rect 3568 11308 7144 11336
rect 3568 11296 3574 11308
rect 6080 11271 6138 11277
rect 6080 11237 6092 11271
rect 6126 11268 6138 11271
rect 6914 11268 6920 11280
rect 6126 11240 6920 11268
rect 6126 11237 6138 11240
rect 6080 11231 6138 11237
rect 6914 11228 6920 11240
rect 6972 11228 6978 11280
rect 3329 11203 3387 11209
rect 3329 11169 3341 11203
rect 3375 11200 3387 11203
rect 3418 11200 3424 11212
rect 3375 11172 3424 11200
rect 3375 11169 3387 11172
rect 3329 11163 3387 11169
rect 3418 11160 3424 11172
rect 3476 11200 3482 11212
rect 4617 11203 4675 11209
rect 4617 11200 4629 11203
rect 3476 11172 4629 11200
rect 3476 11160 3482 11172
rect 4617 11169 4629 11172
rect 4663 11169 4675 11203
rect 7116 11200 7144 11308
rect 7193 11305 7205 11339
rect 7239 11336 7251 11339
rect 8018 11336 8024 11348
rect 7239 11308 8024 11336
rect 7239 11305 7251 11308
rect 7193 11299 7251 11305
rect 8018 11296 8024 11308
rect 8076 11296 8082 11348
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 9398 11336 9404 11348
rect 9088 11308 9404 11336
rect 9088 11296 9094 11308
rect 9398 11296 9404 11308
rect 9456 11336 9462 11348
rect 10597 11339 10655 11345
rect 10597 11336 10609 11339
rect 9456 11308 10609 11336
rect 9456 11296 9462 11308
rect 10597 11305 10609 11308
rect 10643 11305 10655 11339
rect 10597 11299 10655 11305
rect 12253 11339 12311 11345
rect 12253 11305 12265 11339
rect 12299 11336 12311 11339
rect 12299 11308 12480 11336
rect 12299 11305 12311 11308
rect 12253 11299 12311 11305
rect 8110 11228 8116 11280
rect 8168 11268 8174 11280
rect 8389 11271 8447 11277
rect 8389 11268 8401 11271
rect 8168 11240 8401 11268
rect 8168 11228 8174 11240
rect 8389 11237 8401 11240
rect 8435 11237 8447 11271
rect 9306 11268 9312 11280
rect 8389 11231 8447 11237
rect 8496 11240 9312 11268
rect 7116 11172 8156 11200
rect 4617 11163 4675 11169
rect 5810 11092 5816 11144
rect 5868 11092 5874 11144
rect 7282 11092 7288 11144
rect 7340 11092 7346 11144
rect 8128 11132 8156 11172
rect 8202 11160 8208 11212
rect 8260 11160 8266 11212
rect 8496 11209 8524 11240
rect 9306 11228 9312 11240
rect 9364 11228 9370 11280
rect 9484 11271 9542 11277
rect 9484 11237 9496 11271
rect 9530 11268 9542 11271
rect 9674 11268 9680 11280
rect 9530 11240 9680 11268
rect 9530 11237 9542 11240
rect 9484 11231 9542 11237
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11169 8539 11203
rect 8481 11163 8539 11169
rect 8294 11132 8300 11144
rect 8128 11104 8300 11132
rect 8294 11092 8300 11104
rect 8352 11132 8358 11144
rect 8496 11132 8524 11163
rect 8662 11160 8668 11212
rect 8720 11160 8726 11212
rect 8754 11160 8760 11212
rect 8812 11160 8818 11212
rect 8849 11203 8907 11209
rect 8849 11169 8861 11203
rect 8895 11169 8907 11203
rect 8849 11163 8907 11169
rect 8352 11104 8524 11132
rect 8352 11092 8358 11104
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 8864 11132 8892 11163
rect 8628 11104 8892 11132
rect 9217 11135 9275 11141
rect 8628 11092 8634 11104
rect 9217 11101 9229 11135
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 4798 11024 4804 11076
rect 4856 11024 4862 11076
rect 6822 11024 6828 11076
rect 6880 11064 6886 11076
rect 8021 11067 8079 11073
rect 8021 11064 8033 11067
rect 6880 11036 8033 11064
rect 6880 11024 6886 11036
rect 8021 11033 8033 11036
rect 8067 11033 8079 11067
rect 8021 11027 8079 11033
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 7466 10996 7472 11008
rect 6788 10968 7472 10996
rect 6788 10956 6794 10968
rect 7466 10956 7472 10968
rect 7524 10956 7530 11008
rect 7926 10956 7932 11008
rect 7984 10956 7990 11008
rect 9122 10956 9128 11008
rect 9180 10956 9186 11008
rect 9232 10996 9260 11095
rect 10612 11064 10640 11299
rect 12452 11268 12480 11308
rect 13722 11296 13728 11348
rect 13780 11296 13786 11348
rect 18046 11296 18052 11348
rect 18104 11336 18110 11348
rect 18104 11308 18460 11336
rect 18104 11296 18110 11308
rect 12590 11271 12648 11277
rect 12590 11268 12602 11271
rect 12452 11240 12602 11268
rect 12590 11237 12602 11240
rect 12636 11237 12648 11271
rect 12590 11231 12648 11237
rect 12710 11228 12716 11280
rect 12768 11228 12774 11280
rect 13909 11271 13967 11277
rect 13909 11237 13921 11271
rect 13955 11268 13967 11271
rect 18432 11268 18460 11308
rect 18506 11296 18512 11348
rect 18564 11296 18570 11348
rect 19242 11296 19248 11348
rect 19300 11336 19306 11348
rect 19702 11336 19708 11348
rect 19300 11308 19708 11336
rect 19300 11296 19306 11308
rect 19702 11296 19708 11308
rect 19760 11296 19766 11348
rect 19794 11296 19800 11348
rect 19852 11336 19858 11348
rect 20073 11339 20131 11345
rect 20073 11336 20085 11339
rect 19852 11308 20085 11336
rect 19852 11296 19858 11308
rect 20073 11305 20085 11308
rect 20119 11305 20131 11339
rect 20073 11299 20131 11305
rect 21266 11296 21272 11348
rect 21324 11296 21330 11348
rect 24121 11339 24179 11345
rect 24121 11305 24133 11339
rect 24167 11336 24179 11339
rect 24394 11336 24400 11348
rect 24167 11308 24400 11336
rect 24167 11305 24179 11308
rect 24121 11299 24179 11305
rect 24394 11296 24400 11308
rect 24452 11296 24458 11348
rect 26234 11296 26240 11348
rect 26292 11296 26298 11348
rect 19426 11268 19432 11280
rect 13955 11240 14136 11268
rect 13955 11237 13967 11240
rect 13909 11231 13967 11237
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 12345 11203 12403 11209
rect 12345 11200 12357 11203
rect 11572 11172 12357 11200
rect 11572 11160 11578 11172
rect 12345 11169 12357 11172
rect 12391 11169 12403 11203
rect 12728 11200 12756 11228
rect 14108 11209 14136 11240
rect 18432 11240 19432 11268
rect 12345 11163 12403 11169
rect 12452 11172 12756 11200
rect 14001 11203 14059 11209
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11132 11759 11135
rect 12452 11132 12480 11172
rect 14001 11169 14013 11203
rect 14047 11169 14059 11203
rect 14001 11163 14059 11169
rect 14093 11203 14151 11209
rect 14093 11169 14105 11203
rect 14139 11200 14151 11203
rect 14182 11200 14188 11212
rect 14139 11172 14188 11200
rect 14139 11169 14151 11172
rect 14093 11163 14151 11169
rect 11747 11104 12480 11132
rect 14016 11132 14044 11163
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 14826 11160 14832 11212
rect 14884 11200 14890 11212
rect 15105 11203 15163 11209
rect 15105 11200 15117 11203
rect 14884 11172 15117 11200
rect 14884 11160 14890 11172
rect 15105 11169 15117 11172
rect 15151 11169 15163 11203
rect 15105 11163 15163 11169
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11200 15347 11203
rect 15562 11200 15568 11212
rect 15335 11172 15568 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 15562 11160 15568 11172
rect 15620 11160 15626 11212
rect 17126 11160 17132 11212
rect 17184 11200 17190 11212
rect 18049 11203 18107 11209
rect 18049 11200 18061 11203
rect 17184 11172 18061 11200
rect 17184 11160 17190 11172
rect 18049 11169 18061 11172
rect 18095 11169 18107 11203
rect 18049 11163 18107 11169
rect 18141 11203 18199 11209
rect 18141 11169 18153 11203
rect 18187 11169 18199 11203
rect 18141 11163 18199 11169
rect 18325 11203 18383 11209
rect 18325 11169 18337 11203
rect 18371 11200 18383 11203
rect 18432 11200 18460 11240
rect 19426 11228 19432 11240
rect 19484 11228 19490 11280
rect 18371 11172 18460 11200
rect 18371 11169 18383 11172
rect 18325 11163 18383 11169
rect 14458 11132 14464 11144
rect 14016 11104 14464 11132
rect 11747 11101 11759 11104
rect 11701 11095 11759 11101
rect 14458 11092 14464 11104
rect 14516 11092 14522 11144
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11132 14795 11135
rect 14918 11132 14924 11144
rect 14783 11104 14924 11132
rect 14783 11101 14795 11104
rect 14737 11095 14795 11101
rect 14918 11092 14924 11104
rect 14976 11092 14982 11144
rect 15746 11132 15752 11144
rect 15028 11104 15752 11132
rect 15028 11064 15056 11104
rect 15746 11092 15752 11104
rect 15804 11132 15810 11144
rect 16206 11132 16212 11144
rect 15804 11104 16212 11132
rect 15804 11092 15810 11104
rect 16206 11092 16212 11104
rect 16264 11092 16270 11144
rect 16942 11092 16948 11144
rect 17000 11132 17006 11144
rect 17957 11135 18015 11141
rect 17957 11132 17969 11135
rect 17000 11104 17969 11132
rect 17000 11092 17006 11104
rect 17957 11101 17969 11104
rect 18003 11101 18015 11135
rect 17957 11095 18015 11101
rect 10612 11036 12388 11064
rect 9582 10996 9588 11008
rect 9232 10968 9588 10996
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 12360 10996 12388 11036
rect 13280 11036 15056 11064
rect 15473 11067 15531 11073
rect 13280 10996 13308 11036
rect 15473 11033 15485 11067
rect 15519 11064 15531 11067
rect 18046 11064 18052 11076
rect 15519 11036 18052 11064
rect 15519 11033 15531 11036
rect 15473 11027 15531 11033
rect 18046 11024 18052 11036
rect 18104 11024 18110 11076
rect 18156 11064 18184 11163
rect 18598 11160 18604 11212
rect 18656 11160 18662 11212
rect 18782 11160 18788 11212
rect 18840 11160 18846 11212
rect 18874 11160 18880 11212
rect 18932 11160 18938 11212
rect 18969 11203 19027 11209
rect 18969 11169 18981 11203
rect 19015 11200 19027 11203
rect 19812 11200 19840 11296
rect 19886 11228 19892 11280
rect 19944 11268 19950 11280
rect 19944 11240 22048 11268
rect 19944 11228 19950 11240
rect 19015 11172 19840 11200
rect 19015 11169 19027 11172
rect 18969 11163 19027 11169
rect 20438 11160 20444 11212
rect 20496 11200 20502 11212
rect 20496 11172 20852 11200
rect 20496 11160 20502 11172
rect 19245 11135 19303 11141
rect 19245 11101 19257 11135
rect 19291 11132 19303 11135
rect 19889 11135 19947 11141
rect 19889 11132 19901 11135
rect 19291 11104 19901 11132
rect 19291 11101 19303 11104
rect 19245 11095 19303 11101
rect 19889 11101 19901 11104
rect 19935 11101 19947 11135
rect 19889 11095 19947 11101
rect 20714 11092 20720 11144
rect 20772 11092 20778 11144
rect 20824 11132 20852 11172
rect 21450 11160 21456 11212
rect 21508 11200 21514 11212
rect 21652 11209 21680 11240
rect 21545 11203 21603 11209
rect 21545 11200 21557 11203
rect 21508 11172 21557 11200
rect 21508 11160 21514 11172
rect 21545 11169 21557 11172
rect 21591 11169 21603 11203
rect 21545 11163 21603 11169
rect 21637 11203 21695 11209
rect 21637 11169 21649 11203
rect 21683 11169 21695 11203
rect 21637 11163 21695 11169
rect 21726 11160 21732 11212
rect 21784 11160 21790 11212
rect 21913 11203 21971 11209
rect 21913 11169 21925 11203
rect 21959 11169 21971 11203
rect 21913 11163 21971 11169
rect 21928 11132 21956 11163
rect 20824 11104 21956 11132
rect 21358 11064 21364 11076
rect 18156 11036 21364 11064
rect 21358 11024 21364 11036
rect 21416 11024 21422 11076
rect 22020 11064 22048 11240
rect 22097 11203 22155 11209
rect 22097 11169 22109 11203
rect 22143 11200 22155 11203
rect 22278 11200 22284 11212
rect 22143 11172 22284 11200
rect 22143 11169 22155 11172
rect 22097 11163 22155 11169
rect 22278 11160 22284 11172
rect 22336 11200 22342 11212
rect 22830 11200 22836 11212
rect 22336 11172 22836 11200
rect 22336 11160 22342 11172
rect 22830 11160 22836 11172
rect 22888 11160 22894 11212
rect 23008 11203 23066 11209
rect 23008 11169 23020 11203
rect 23054 11200 23066 11203
rect 23750 11200 23756 11212
rect 23054 11172 23756 11200
rect 23054 11169 23066 11172
rect 23008 11163 23066 11169
rect 23750 11160 23756 11172
rect 23808 11160 23814 11212
rect 24854 11160 24860 11212
rect 24912 11160 24918 11212
rect 25124 11203 25182 11209
rect 25124 11169 25136 11203
rect 25170 11200 25182 11203
rect 26421 11203 26479 11209
rect 26421 11200 26433 11203
rect 25170 11172 26433 11200
rect 25170 11169 25182 11172
rect 25124 11163 25182 11169
rect 26421 11169 26433 11172
rect 26467 11169 26479 11203
rect 26421 11163 26479 11169
rect 22738 11092 22744 11144
rect 22796 11092 22802 11144
rect 25866 11092 25872 11144
rect 25924 11132 25930 11144
rect 26973 11135 27031 11141
rect 26973 11132 26985 11135
rect 25924 11104 26985 11132
rect 25924 11092 25930 11104
rect 26973 11101 26985 11104
rect 27019 11101 27031 11135
rect 26973 11095 27031 11101
rect 22646 11064 22652 11076
rect 22020 11036 22652 11064
rect 22646 11024 22652 11036
rect 22704 11024 22710 11076
rect 12360 10968 13308 10996
rect 14277 10999 14335 11005
rect 14277 10965 14289 10999
rect 14323 10996 14335 10999
rect 14366 10996 14372 11008
rect 14323 10968 14372 10996
rect 14323 10965 14335 10968
rect 14277 10959 14335 10965
rect 14366 10956 14372 10968
rect 14424 10956 14430 11008
rect 17313 10999 17371 11005
rect 17313 10965 17325 10999
rect 17359 10996 17371 10999
rect 17586 10996 17592 11008
rect 17359 10968 17592 10996
rect 17359 10965 17371 10968
rect 17313 10959 17371 10965
rect 17586 10956 17592 10968
rect 17644 10956 17650 11008
rect 19334 10956 19340 11008
rect 19392 10956 19398 11008
rect 22281 10999 22339 11005
rect 22281 10965 22293 10999
rect 22327 10996 22339 10999
rect 22922 10996 22928 11008
rect 22327 10968 22928 10996
rect 22327 10965 22339 10968
rect 22281 10959 22339 10965
rect 22922 10956 22928 10968
rect 22980 10956 22986 11008
rect 552 10906 27416 10928
rect 552 10854 3756 10906
rect 3808 10854 3820 10906
rect 3872 10854 3884 10906
rect 3936 10854 3948 10906
rect 4000 10854 4012 10906
rect 4064 10854 10472 10906
rect 10524 10854 10536 10906
rect 10588 10854 10600 10906
rect 10652 10854 10664 10906
rect 10716 10854 10728 10906
rect 10780 10854 17188 10906
rect 17240 10854 17252 10906
rect 17304 10854 17316 10906
rect 17368 10854 17380 10906
rect 17432 10854 17444 10906
rect 17496 10854 23904 10906
rect 23956 10854 23968 10906
rect 24020 10854 24032 10906
rect 24084 10854 24096 10906
rect 24148 10854 24160 10906
rect 24212 10854 27416 10906
rect 552 10832 27416 10854
rect 7193 10795 7251 10801
rect 7193 10761 7205 10795
rect 7239 10792 7251 10795
rect 7282 10792 7288 10804
rect 7239 10764 7288 10792
rect 7239 10761 7251 10764
rect 7193 10755 7251 10761
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 8205 10795 8263 10801
rect 8205 10761 8217 10795
rect 8251 10792 8263 10795
rect 8662 10792 8668 10804
rect 8251 10764 8668 10792
rect 8251 10761 8263 10764
rect 8205 10755 8263 10761
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 8772 10764 10977 10792
rect 8772 10724 8800 10764
rect 7760 10696 8800 10724
rect 7760 10600 7788 10696
rect 8846 10684 8852 10736
rect 8904 10684 8910 10736
rect 8864 10656 8892 10684
rect 8128 10628 8892 10656
rect 9140 10656 9168 10764
rect 10965 10761 10977 10764
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 12437 10795 12495 10801
rect 12437 10761 12449 10795
rect 12483 10792 12495 10795
rect 12710 10792 12716 10804
rect 12483 10764 12716 10792
rect 12483 10761 12495 10764
rect 12437 10755 12495 10761
rect 9140 10628 9260 10656
rect 2406 10548 2412 10600
rect 2464 10588 2470 10600
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 2464 10560 4353 10588
rect 2464 10548 2470 10560
rect 4341 10557 4353 10560
rect 4387 10588 4399 10591
rect 5810 10588 5816 10600
rect 4387 10560 5816 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 5810 10548 5816 10560
rect 5868 10548 5874 10600
rect 7742 10597 7748 10600
rect 7561 10591 7619 10597
rect 7561 10557 7573 10591
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7709 10591 7748 10597
rect 7709 10557 7721 10591
rect 7709 10551 7748 10557
rect 4608 10523 4666 10529
rect 4608 10489 4620 10523
rect 4654 10520 4666 10523
rect 5626 10520 5632 10532
rect 4654 10492 5632 10520
rect 4654 10489 4666 10492
rect 4608 10483 4666 10489
rect 5626 10480 5632 10492
rect 5684 10480 5690 10532
rect 6086 10529 6092 10532
rect 6080 10483 6092 10529
rect 6086 10480 6092 10483
rect 6144 10480 6150 10532
rect 5718 10412 5724 10464
rect 5776 10412 5782 10464
rect 7576 10452 7604 10551
rect 7742 10548 7748 10551
rect 7800 10548 7806 10600
rect 7926 10548 7932 10600
rect 7984 10548 7990 10600
rect 8026 10591 8084 10597
rect 8026 10557 8038 10591
rect 8072 10588 8084 10591
rect 8128 10588 8156 10628
rect 8072 10560 8156 10588
rect 8072 10557 8084 10560
rect 8026 10551 8084 10557
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 8570 10588 8576 10600
rect 8352 10560 8576 10588
rect 8352 10548 8358 10560
rect 8570 10548 8576 10560
rect 8628 10588 8634 10600
rect 8849 10591 8907 10597
rect 8849 10588 8861 10591
rect 8628 10560 8861 10588
rect 8628 10548 8634 10560
rect 8849 10557 8861 10560
rect 8895 10557 8907 10591
rect 8849 10551 8907 10557
rect 8938 10548 8944 10600
rect 8996 10588 9002 10600
rect 9232 10597 9260 10628
rect 9033 10591 9091 10597
rect 9033 10588 9045 10591
rect 8996 10560 9045 10588
rect 8996 10548 9002 10560
rect 9033 10557 9045 10560
rect 9079 10557 9091 10591
rect 9033 10551 9091 10557
rect 9125 10591 9183 10597
rect 9125 10557 9137 10591
rect 9171 10557 9183 10591
rect 9125 10551 9183 10557
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10557 9275 10591
rect 9217 10551 9275 10557
rect 7837 10523 7895 10529
rect 7837 10489 7849 10523
rect 7883 10520 7895 10523
rect 8478 10520 8484 10532
rect 7883 10492 8484 10520
rect 7883 10489 7895 10492
rect 7837 10483 7895 10489
rect 8478 10480 8484 10492
rect 8536 10480 8542 10532
rect 8754 10480 8760 10532
rect 8812 10520 8818 10532
rect 9140 10520 9168 10551
rect 9582 10548 9588 10600
rect 9640 10548 9646 10600
rect 9493 10523 9551 10529
rect 8812 10492 9260 10520
rect 8812 10480 8818 10492
rect 9232 10464 9260 10492
rect 9493 10489 9505 10523
rect 9539 10520 9551 10523
rect 9830 10523 9888 10529
rect 9830 10520 9842 10523
rect 9539 10492 9842 10520
rect 9539 10489 9551 10492
rect 9493 10483 9551 10489
rect 9830 10489 9842 10492
rect 9876 10489 9888 10523
rect 10980 10520 11008 10755
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 14829 10795 14887 10801
rect 14829 10761 14841 10795
rect 14875 10792 14887 10795
rect 15194 10792 15200 10804
rect 14875 10764 15200 10792
rect 14875 10761 14887 10764
rect 14829 10755 14887 10761
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 15304 10764 16804 10792
rect 12526 10684 12532 10736
rect 12584 10724 12590 10736
rect 15304 10724 15332 10764
rect 12584 10696 15332 10724
rect 16776 10724 16804 10764
rect 16942 10752 16948 10804
rect 17000 10792 17006 10804
rect 17221 10795 17279 10801
rect 17221 10792 17233 10795
rect 17000 10764 17233 10792
rect 17000 10752 17006 10764
rect 17221 10761 17233 10764
rect 17267 10761 17279 10795
rect 19978 10792 19984 10804
rect 17221 10755 17279 10761
rect 17328 10764 19984 10792
rect 17328 10724 17356 10764
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 20073 10795 20131 10801
rect 20073 10761 20085 10795
rect 20119 10792 20131 10795
rect 20714 10792 20720 10804
rect 20119 10764 20720 10792
rect 20119 10761 20131 10764
rect 20073 10755 20131 10761
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 21726 10752 21732 10804
rect 21784 10792 21790 10804
rect 22005 10795 22063 10801
rect 22005 10792 22017 10795
rect 21784 10764 22017 10792
rect 21784 10752 21790 10764
rect 22005 10761 22017 10764
rect 22051 10761 22063 10795
rect 23566 10792 23572 10804
rect 22005 10755 22063 10761
rect 22388 10764 23572 10792
rect 16776 10696 17356 10724
rect 12584 10684 12590 10696
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 12820 10597 12848 10696
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10656 14335 10659
rect 14366 10656 14372 10668
rect 14323 10628 14372 10656
rect 14323 10625 14335 10628
rect 14277 10619 14335 10625
rect 14366 10616 14372 10628
rect 14424 10656 14430 10668
rect 14826 10656 14832 10668
rect 14424 10628 14832 10656
rect 14424 10616 14430 10628
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 15102 10616 15108 10668
rect 15160 10656 15166 10668
rect 18690 10656 18696 10668
rect 15160 10628 15332 10656
rect 15160 10616 15166 10628
rect 15304 10600 15332 10628
rect 17788 10628 18696 10656
rect 12713 10591 12771 10597
rect 12713 10588 12725 10591
rect 12676 10560 12725 10588
rect 12676 10548 12682 10560
rect 12713 10557 12725 10560
rect 12759 10557 12771 10591
rect 12713 10551 12771 10557
rect 12805 10591 12863 10597
rect 12805 10557 12817 10591
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 12894 10548 12900 10600
rect 12952 10548 12958 10600
rect 13078 10548 13084 10600
rect 13136 10548 13142 10600
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 15028 10520 15056 10551
rect 15194 10548 15200 10600
rect 15252 10548 15258 10600
rect 15286 10548 15292 10600
rect 15344 10548 15350 10600
rect 15378 10548 15384 10600
rect 15436 10548 15442 10600
rect 15841 10591 15899 10597
rect 15841 10557 15853 10591
rect 15887 10588 15899 10591
rect 17788 10588 17816 10628
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 15887 10560 17816 10588
rect 15887 10557 15899 10560
rect 15841 10551 15899 10557
rect 17862 10548 17868 10600
rect 17920 10548 17926 10600
rect 18960 10591 19018 10597
rect 18960 10557 18972 10591
rect 19006 10588 19018 10591
rect 19334 10588 19340 10600
rect 19006 10560 19340 10588
rect 19006 10557 19018 10560
rect 18960 10551 19018 10557
rect 19334 10548 19340 10560
rect 19392 10548 19398 10600
rect 19426 10548 19432 10600
rect 19484 10588 19490 10600
rect 20165 10591 20223 10597
rect 20165 10588 20177 10591
rect 19484 10560 20177 10588
rect 19484 10548 19490 10560
rect 20165 10557 20177 10560
rect 20211 10557 20223 10591
rect 22186 10588 22192 10600
rect 20165 10551 20223 10557
rect 21744 10560 22192 10588
rect 15746 10520 15752 10532
rect 10980 10492 14504 10520
rect 15028 10492 15752 10520
rect 9830 10483 9888 10489
rect 8294 10452 8300 10464
rect 7576 10424 8300 10452
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 9214 10412 9220 10464
rect 9272 10412 9278 10464
rect 14366 10412 14372 10464
rect 14424 10412 14430 10464
rect 14476 10461 14504 10492
rect 15746 10480 15752 10492
rect 15804 10480 15810 10532
rect 15930 10480 15936 10532
rect 15988 10520 15994 10532
rect 16086 10523 16144 10529
rect 16086 10520 16098 10523
rect 15988 10492 16098 10520
rect 15988 10480 15994 10492
rect 16086 10489 16098 10492
rect 16132 10489 16144 10523
rect 16086 10483 16144 10489
rect 21744 10464 21772 10560
rect 22186 10548 22192 10560
rect 22244 10548 22250 10600
rect 22388 10597 22416 10764
rect 23566 10752 23572 10764
rect 23624 10752 23630 10804
rect 23750 10752 23756 10804
rect 23808 10792 23814 10804
rect 23845 10795 23903 10801
rect 23845 10792 23857 10795
rect 23808 10764 23857 10792
rect 23808 10752 23814 10764
rect 23845 10761 23857 10764
rect 23891 10761 23903 10795
rect 23845 10755 23903 10761
rect 26418 10752 26424 10804
rect 26476 10792 26482 10804
rect 26605 10795 26663 10801
rect 26605 10792 26617 10795
rect 26476 10764 26617 10792
rect 26476 10752 26482 10764
rect 26605 10761 26617 10764
rect 26651 10761 26663 10795
rect 26605 10755 26663 10761
rect 22646 10684 22652 10736
rect 22704 10724 22710 10736
rect 25038 10724 25044 10736
rect 22704 10696 25044 10724
rect 22704 10684 22710 10696
rect 22373 10591 22431 10597
rect 22373 10557 22385 10591
rect 22419 10557 22431 10591
rect 22373 10551 22431 10557
rect 22465 10591 22523 10597
rect 22465 10557 22477 10591
rect 22511 10557 22523 10591
rect 22465 10551 22523 10557
rect 22002 10480 22008 10532
rect 22060 10520 22066 10532
rect 22480 10520 22508 10551
rect 22922 10548 22928 10600
rect 22980 10548 22986 10600
rect 23216 10597 23244 10696
rect 25038 10684 25044 10696
rect 25096 10684 25102 10736
rect 23569 10659 23627 10665
rect 23569 10625 23581 10659
rect 23615 10656 23627 10659
rect 24397 10659 24455 10665
rect 24397 10656 24409 10659
rect 23615 10628 24409 10656
rect 23615 10625 23627 10628
rect 23569 10619 23627 10625
rect 24397 10625 24409 10628
rect 24443 10625 24455 10659
rect 24397 10619 24455 10625
rect 24854 10616 24860 10668
rect 24912 10656 24918 10668
rect 25225 10659 25283 10665
rect 25225 10656 25237 10659
rect 24912 10628 25237 10656
rect 24912 10616 24918 10628
rect 25225 10625 25237 10628
rect 25271 10625 25283 10659
rect 25225 10619 25283 10625
rect 23109 10591 23167 10597
rect 23109 10557 23121 10591
rect 23155 10557 23167 10591
rect 23109 10551 23167 10557
rect 23201 10591 23259 10597
rect 23201 10557 23213 10591
rect 23247 10557 23259 10591
rect 23201 10551 23259 10557
rect 23293 10591 23351 10597
rect 23293 10557 23305 10591
rect 23339 10588 23351 10591
rect 23658 10588 23664 10600
rect 23339 10560 23664 10588
rect 23339 10557 23351 10560
rect 23293 10551 23351 10557
rect 22060 10492 22508 10520
rect 22060 10480 22066 10492
rect 14461 10455 14519 10461
rect 14461 10421 14473 10455
rect 14507 10452 14519 10455
rect 15010 10452 15016 10464
rect 14507 10424 15016 10452
rect 14507 10421 14519 10424
rect 14461 10415 14519 10421
rect 15010 10412 15016 10424
rect 15068 10412 15074 10464
rect 15657 10455 15715 10461
rect 15657 10421 15669 10455
rect 15703 10452 15715 10455
rect 16666 10452 16672 10464
rect 15703 10424 16672 10452
rect 15703 10421 15715 10424
rect 15657 10415 15715 10421
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 17310 10412 17316 10464
rect 17368 10412 17374 10464
rect 19886 10412 19892 10464
rect 19944 10452 19950 10464
rect 20349 10455 20407 10461
rect 20349 10452 20361 10455
rect 19944 10424 20361 10452
rect 19944 10412 19950 10424
rect 20349 10421 20361 10424
rect 20395 10452 20407 10455
rect 21726 10452 21732 10464
rect 20395 10424 21732 10452
rect 20395 10421 20407 10424
rect 20349 10415 20407 10421
rect 21726 10412 21732 10424
rect 21784 10412 21790 10464
rect 22940 10452 22968 10548
rect 23124 10520 23152 10551
rect 23658 10548 23664 10560
rect 23716 10548 23722 10600
rect 24486 10548 24492 10600
rect 24544 10588 24550 10600
rect 24765 10591 24823 10597
rect 24765 10588 24777 10591
rect 24544 10560 24777 10588
rect 24544 10548 24550 10560
rect 24765 10557 24777 10560
rect 24811 10557 24823 10591
rect 24765 10551 24823 10557
rect 24946 10548 24952 10600
rect 25004 10588 25010 10600
rect 25041 10591 25099 10597
rect 25041 10588 25053 10591
rect 25004 10560 25053 10588
rect 25004 10548 25010 10560
rect 25041 10557 25053 10560
rect 25087 10557 25099 10591
rect 25041 10551 25099 10557
rect 24581 10523 24639 10529
rect 24581 10520 24593 10523
rect 23124 10492 24593 10520
rect 24581 10489 24593 10492
rect 24627 10489 24639 10523
rect 24581 10483 24639 10489
rect 24670 10480 24676 10532
rect 24728 10520 24734 10532
rect 25470 10523 25528 10529
rect 25470 10520 25482 10523
rect 24728 10492 25482 10520
rect 24728 10480 24734 10492
rect 25470 10489 25482 10492
rect 25516 10489 25528 10523
rect 25470 10483 25528 10489
rect 24118 10452 24124 10464
rect 22940 10424 24124 10452
rect 24118 10412 24124 10424
rect 24176 10412 24182 10464
rect 24949 10455 25007 10461
rect 24949 10421 24961 10455
rect 24995 10452 25007 10455
rect 25314 10452 25320 10464
rect 24995 10424 25320 10452
rect 24995 10421 25007 10424
rect 24949 10415 25007 10421
rect 25314 10412 25320 10424
rect 25372 10412 25378 10464
rect 552 10362 27576 10384
rect 552 10310 7114 10362
rect 7166 10310 7178 10362
rect 7230 10310 7242 10362
rect 7294 10310 7306 10362
rect 7358 10310 7370 10362
rect 7422 10310 13830 10362
rect 13882 10310 13894 10362
rect 13946 10310 13958 10362
rect 14010 10310 14022 10362
rect 14074 10310 14086 10362
rect 14138 10310 20546 10362
rect 20598 10310 20610 10362
rect 20662 10310 20674 10362
rect 20726 10310 20738 10362
rect 20790 10310 20802 10362
rect 20854 10310 27262 10362
rect 27314 10310 27326 10362
rect 27378 10310 27390 10362
rect 27442 10310 27454 10362
rect 27506 10310 27518 10362
rect 27570 10310 27576 10362
rect 552 10288 27576 10310
rect 2133 10251 2191 10257
rect 2133 10217 2145 10251
rect 2179 10248 2191 10251
rect 3602 10248 3608 10260
rect 2179 10220 3608 10248
rect 2179 10217 2191 10220
rect 2133 10211 2191 10217
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 5997 10251 6055 10257
rect 5997 10217 6009 10251
rect 6043 10248 6055 10251
rect 6086 10248 6092 10260
rect 6043 10220 6092 10248
rect 6043 10217 6055 10220
rect 5997 10211 6055 10217
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 7929 10251 7987 10257
rect 7929 10217 7941 10251
rect 7975 10248 7987 10251
rect 8202 10248 8208 10260
rect 7975 10220 8208 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 8754 10248 8760 10260
rect 8628 10220 8760 10248
rect 8628 10208 8634 10220
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 8938 10208 8944 10260
rect 8996 10208 9002 10260
rect 12158 10208 12164 10260
rect 12216 10208 12222 10260
rect 12805 10251 12863 10257
rect 12805 10217 12817 10251
rect 12851 10248 12863 10251
rect 12894 10248 12900 10260
rect 12851 10220 12900 10248
rect 12851 10217 12863 10220
rect 12805 10211 12863 10217
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 12986 10208 12992 10260
rect 13044 10248 13050 10260
rect 13357 10251 13415 10257
rect 13357 10248 13369 10251
rect 13044 10220 13369 10248
rect 13044 10208 13050 10220
rect 13357 10217 13369 10220
rect 13403 10217 13415 10251
rect 13357 10211 13415 10217
rect 14185 10251 14243 10257
rect 14185 10217 14197 10251
rect 14231 10248 14243 10251
rect 14550 10248 14556 10260
rect 14231 10220 14556 10248
rect 14231 10217 14243 10220
rect 14185 10211 14243 10217
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 15378 10208 15384 10260
rect 15436 10248 15442 10260
rect 15657 10251 15715 10257
rect 15657 10248 15669 10251
rect 15436 10220 15669 10248
rect 15436 10208 15442 10220
rect 15657 10217 15669 10220
rect 15703 10217 15715 10251
rect 15657 10211 15715 10217
rect 15841 10251 15899 10257
rect 15841 10217 15853 10251
rect 15887 10248 15899 10251
rect 15930 10248 15936 10260
rect 15887 10220 15936 10248
rect 15887 10217 15899 10220
rect 15841 10211 15899 10217
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 17310 10208 17316 10260
rect 17368 10208 17374 10260
rect 20254 10208 20260 10260
rect 20312 10208 20318 10260
rect 21818 10208 21824 10260
rect 21876 10248 21882 10260
rect 21913 10251 21971 10257
rect 21913 10248 21925 10251
rect 21876 10220 21925 10248
rect 21876 10208 21882 10220
rect 21913 10217 21925 10220
rect 21959 10217 21971 10251
rect 21913 10211 21971 10217
rect 22094 10208 22100 10260
rect 22152 10208 22158 10260
rect 22925 10251 22983 10257
rect 22925 10217 22937 10251
rect 22971 10248 22983 10251
rect 23014 10248 23020 10260
rect 22971 10220 23020 10248
rect 22971 10217 22983 10220
rect 22925 10211 22983 10217
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 23290 10208 23296 10260
rect 23348 10208 23354 10260
rect 25409 10251 25467 10257
rect 25409 10217 25421 10251
rect 25455 10248 25467 10251
rect 25866 10248 25872 10260
rect 25455 10220 25872 10248
rect 25455 10217 25467 10220
rect 25409 10211 25467 10217
rect 25866 10208 25872 10220
rect 25924 10208 25930 10260
rect 2676 10183 2734 10189
rect 2676 10149 2688 10183
rect 2722 10180 2734 10183
rect 2866 10180 2872 10192
rect 2722 10152 2872 10180
rect 2722 10149 2734 10152
rect 2676 10143 2734 10149
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 5718 10140 5724 10192
rect 5776 10180 5782 10192
rect 8220 10180 8248 10208
rect 8665 10183 8723 10189
rect 8665 10180 8677 10183
rect 5776 10152 7328 10180
rect 8220 10152 8677 10180
rect 5776 10140 5782 10152
rect 2406 10072 2412 10124
rect 2464 10072 2470 10124
rect 3418 10112 3424 10124
rect 2516 10084 3424 10112
rect 2516 10044 2544 10084
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 4985 10115 5043 10121
rect 4985 10081 4997 10115
rect 5031 10112 5043 10115
rect 5442 10112 5448 10124
rect 5031 10084 5448 10112
rect 5031 10081 5043 10084
rect 4985 10075 5043 10081
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 6086 10072 6092 10124
rect 6144 10112 6150 10124
rect 6181 10115 6239 10121
rect 6181 10112 6193 10115
rect 6144 10084 6193 10112
rect 6144 10072 6150 10084
rect 6181 10081 6193 10084
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 6457 10115 6515 10121
rect 6457 10081 6469 10115
rect 6503 10112 6515 10115
rect 6503 10084 6592 10112
rect 6503 10081 6515 10084
rect 6457 10075 6515 10081
rect 4801 10047 4859 10053
rect 4801 10044 4813 10047
rect 2148 10016 2544 10044
rect 4172 10016 4813 10044
rect 1765 9979 1823 9985
rect 1765 9945 1777 9979
rect 1811 9976 1823 9979
rect 1854 9976 1860 9988
rect 1811 9948 1860 9976
rect 1811 9945 1823 9948
rect 1765 9939 1823 9945
rect 1854 9936 1860 9948
rect 1912 9936 1918 9988
rect 2148 9917 2176 10016
rect 4172 9920 4200 10016
rect 4801 10013 4813 10016
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10013 5319 10047
rect 5261 10007 5319 10013
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10044 5687 10047
rect 6564 10044 6592 10084
rect 6638 10072 6644 10124
rect 6696 10072 6702 10124
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10081 7067 10115
rect 7009 10075 7067 10081
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 5675 10016 6500 10044
rect 6564 10016 6837 10044
rect 5675 10013 5687 10016
rect 5629 10007 5687 10013
rect 4982 9936 4988 9988
rect 5040 9976 5046 9988
rect 5276 9976 5304 10007
rect 5040 9948 5304 9976
rect 6273 9979 6331 9985
rect 5040 9936 5046 9948
rect 6273 9945 6285 9979
rect 6319 9945 6331 9979
rect 6273 9939 6331 9945
rect 2133 9911 2191 9917
rect 2133 9877 2145 9911
rect 2179 9877 2191 9911
rect 2133 9871 2191 9877
rect 2317 9911 2375 9917
rect 2317 9877 2329 9911
rect 2363 9908 2375 9911
rect 3050 9908 3056 9920
rect 2363 9880 3056 9908
rect 2363 9877 2375 9880
rect 2317 9871 2375 9877
rect 3050 9868 3056 9880
rect 3108 9868 3114 9920
rect 3789 9911 3847 9917
rect 3789 9877 3801 9911
rect 3835 9908 3847 9911
rect 4154 9908 4160 9920
rect 3835 9880 4160 9908
rect 3835 9877 3847 9880
rect 3789 9871 3847 9877
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 5169 9911 5227 9917
rect 5169 9877 5181 9911
rect 5215 9908 5227 9911
rect 5534 9908 5540 9920
rect 5215 9880 5540 9908
rect 5215 9877 5227 9880
rect 5169 9871 5227 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 6288 9908 6316 9939
rect 6362 9936 6368 9988
rect 6420 9936 6426 9988
rect 6472 9976 6500 10016
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 7024 10044 7052 10075
rect 7190 10072 7196 10124
rect 7248 10072 7254 10124
rect 7300 10121 7328 10152
rect 8665 10149 8677 10152
rect 8711 10149 8723 10183
rect 9582 10180 9588 10192
rect 8665 10143 8723 10149
rect 9048 10152 9588 10180
rect 7285 10115 7343 10121
rect 7285 10081 7297 10115
rect 7331 10081 7343 10115
rect 7285 10075 7343 10081
rect 8294 10072 8300 10124
rect 8352 10072 8358 10124
rect 8445 10115 8503 10121
rect 8445 10081 8457 10115
rect 8491 10112 8503 10115
rect 8491 10081 8524 10112
rect 8445 10075 8524 10081
rect 7926 10044 7932 10056
rect 7024 10016 7932 10044
rect 6825 10007 6883 10013
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 7650 9976 7656 9988
rect 6472 9948 7656 9976
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 8496 9976 8524 10075
rect 8570 10072 8576 10124
rect 8628 10072 8634 10124
rect 8846 10121 8852 10124
rect 8803 10115 8852 10121
rect 8803 10081 8815 10115
rect 8849 10081 8852 10115
rect 8803 10075 8852 10081
rect 8846 10072 8852 10075
rect 8904 10072 8910 10124
rect 9048 10121 9076 10152
rect 9582 10140 9588 10152
rect 9640 10140 9646 10192
rect 12176 10180 12204 10208
rect 12342 10180 12348 10192
rect 12176 10152 12348 10180
rect 9033 10115 9091 10121
rect 9033 10081 9045 10115
rect 9079 10081 9091 10115
rect 9033 10075 9091 10081
rect 9122 10072 9128 10124
rect 9180 10112 9186 10124
rect 12176 10121 12204 10152
rect 12342 10140 12348 10152
rect 12400 10140 12406 10192
rect 12529 10183 12587 10189
rect 12529 10149 12541 10183
rect 12575 10180 12587 10183
rect 14274 10180 14280 10192
rect 12575 10152 14280 10180
rect 12575 10149 12587 10152
rect 12529 10143 12587 10149
rect 14274 10140 14280 10152
rect 14332 10180 14338 10192
rect 17328 10180 17356 10208
rect 14332 10152 15056 10180
rect 14332 10140 14338 10152
rect 9289 10115 9347 10121
rect 9289 10112 9301 10115
rect 9180 10084 9301 10112
rect 9180 10072 9186 10084
rect 9289 10081 9301 10084
rect 9335 10081 9347 10115
rect 9289 10075 9347 10081
rect 12161 10115 12219 10121
rect 12161 10081 12173 10115
rect 12207 10081 12219 10115
rect 12161 10075 12219 10081
rect 12250 10072 12256 10124
rect 12308 10112 12314 10124
rect 12437 10115 12495 10121
rect 12308 10084 12353 10112
rect 12308 10072 12314 10084
rect 12437 10081 12449 10115
rect 12483 10081 12495 10115
rect 12437 10075 12495 10081
rect 8588 10044 8616 10072
rect 8938 10044 8944 10056
rect 8588 10016 8944 10044
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 12452 10044 12480 10075
rect 12618 10072 12624 10124
rect 12676 10121 12682 10124
rect 12676 10112 12684 10121
rect 12676 10084 12721 10112
rect 12676 10075 12684 10084
rect 12676 10072 12682 10075
rect 13354 10072 13360 10124
rect 13412 10112 13418 10124
rect 15028 10121 15056 10152
rect 15764 10152 17356 10180
rect 18785 10183 18843 10189
rect 15764 10121 15792 10152
rect 18785 10149 18797 10183
rect 18831 10180 18843 10183
rect 19122 10183 19180 10189
rect 19122 10180 19134 10183
rect 18831 10152 19134 10180
rect 18831 10149 18843 10152
rect 18785 10143 18843 10149
rect 19122 10149 19134 10152
rect 19168 10149 19180 10183
rect 19122 10143 19180 10149
rect 13725 10115 13783 10121
rect 13725 10112 13737 10115
rect 13412 10084 13737 10112
rect 13412 10072 13418 10084
rect 13725 10081 13737 10084
rect 13771 10081 13783 10115
rect 14553 10115 14611 10121
rect 14553 10112 14565 10115
rect 13725 10075 13783 10081
rect 13924 10084 14565 10112
rect 13446 10044 13452 10056
rect 12452 10016 13452 10044
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 13817 10047 13875 10053
rect 13817 10044 13829 10047
rect 13740 10016 13829 10044
rect 13740 9988 13768 10016
rect 13817 10013 13829 10016
rect 13863 10013 13875 10047
rect 13817 10007 13875 10013
rect 9030 9976 9036 9988
rect 8496 9948 9036 9976
rect 9030 9936 9036 9948
rect 9088 9936 9094 9988
rect 13722 9936 13728 9988
rect 13780 9936 13786 9988
rect 6454 9908 6460 9920
rect 6288 9880 6460 9908
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 7190 9868 7196 9920
rect 7248 9908 7254 9920
rect 8202 9908 8208 9920
rect 7248 9880 8208 9908
rect 7248 9868 7254 9880
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 10413 9911 10471 9917
rect 10413 9908 10425 9911
rect 8720 9880 10425 9908
rect 8720 9868 8726 9880
rect 10413 9877 10425 9880
rect 10459 9908 10471 9911
rect 13924 9908 13952 10084
rect 14553 10081 14565 10084
rect 14599 10112 14611 10115
rect 15013 10115 15071 10121
rect 14599 10084 14964 10112
rect 14599 10081 14611 10084
rect 14553 10075 14611 10081
rect 14001 10047 14059 10053
rect 14001 10013 14013 10047
rect 14047 10013 14059 10047
rect 14001 10007 14059 10013
rect 14016 9976 14044 10007
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10044 14795 10047
rect 14826 10044 14832 10056
rect 14783 10016 14832 10044
rect 14783 10013 14795 10016
rect 14737 10007 14795 10013
rect 14752 9976 14780 10007
rect 14826 10004 14832 10016
rect 14884 10004 14890 10056
rect 14936 10044 14964 10084
rect 15013 10081 15025 10115
rect 15059 10081 15071 10115
rect 15013 10075 15071 10081
rect 15749 10115 15807 10121
rect 15749 10081 15761 10115
rect 15795 10081 15807 10115
rect 15749 10075 15807 10081
rect 15933 10115 15991 10121
rect 15933 10081 15945 10115
rect 15979 10112 15991 10115
rect 16574 10112 16580 10124
rect 15979 10084 16580 10112
rect 15979 10081 15991 10084
rect 15933 10075 15991 10081
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 16666 10072 16672 10124
rect 16724 10072 16730 10124
rect 16850 10072 16856 10124
rect 16908 10112 16914 10124
rect 17037 10115 17095 10121
rect 17037 10112 17049 10115
rect 16908 10084 17049 10112
rect 16908 10072 16914 10084
rect 17037 10081 17049 10084
rect 17083 10081 17095 10115
rect 17037 10075 17095 10081
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10081 17187 10115
rect 17129 10075 17187 10081
rect 17313 10115 17371 10121
rect 17313 10081 17325 10115
rect 17359 10112 17371 10115
rect 17586 10112 17592 10124
rect 17359 10084 17592 10112
rect 17359 10081 17371 10084
rect 17313 10075 17371 10081
rect 15102 10044 15108 10056
rect 14936 10016 15108 10044
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 17144 10044 17172 10075
rect 17586 10072 17592 10084
rect 17644 10072 17650 10124
rect 18690 10072 18696 10124
rect 18748 10112 18754 10124
rect 18877 10115 18935 10121
rect 18877 10112 18889 10115
rect 18748 10084 18889 10112
rect 18748 10072 18754 10084
rect 18877 10081 18889 10084
rect 18923 10081 18935 10115
rect 20272 10112 20300 10208
rect 21545 10183 21603 10189
rect 21545 10149 21557 10183
rect 21591 10180 21603 10183
rect 22370 10180 22376 10192
rect 21591 10152 22376 10180
rect 21591 10149 21603 10152
rect 21545 10143 21603 10149
rect 22370 10140 22376 10152
rect 22428 10140 22434 10192
rect 22465 10183 22523 10189
rect 22465 10149 22477 10183
rect 22511 10180 22523 10183
rect 23308 10180 23336 10208
rect 24118 10180 24124 10192
rect 22511 10152 23336 10180
rect 22511 10149 22523 10152
rect 22465 10143 22523 10149
rect 24105 10140 24124 10180
rect 24176 10180 24182 10192
rect 24176 10152 24808 10180
rect 24176 10140 24182 10152
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20272 10084 20913 10112
rect 18877 10075 18935 10081
rect 20901 10081 20913 10084
rect 20947 10081 20959 10115
rect 20901 10075 20959 10081
rect 21453 10115 21511 10121
rect 21453 10081 21465 10115
rect 21499 10081 21511 10115
rect 21453 10075 21511 10081
rect 17770 10044 17776 10056
rect 17144 10016 17776 10044
rect 17770 10004 17776 10016
rect 17828 10044 17834 10056
rect 17957 10047 18015 10053
rect 17957 10044 17969 10047
rect 17828 10016 17969 10044
rect 17828 10004 17834 10016
rect 17957 10013 17969 10016
rect 18003 10013 18015 10047
rect 17957 10007 18015 10013
rect 18230 10004 18236 10056
rect 18288 10004 18294 10056
rect 20162 10004 20168 10056
rect 20220 10044 20226 10056
rect 21468 10044 21496 10075
rect 21726 10072 21732 10124
rect 21784 10072 21790 10124
rect 22002 10115 22008 10124
rect 21836 10087 22008 10115
rect 21836 10044 21864 10087
rect 22002 10072 22008 10087
rect 22060 10072 22066 10124
rect 22186 10072 22192 10124
rect 22244 10112 22250 10124
rect 22281 10115 22339 10121
rect 22281 10112 22293 10115
rect 22244 10084 22293 10112
rect 22244 10072 22250 10084
rect 22281 10081 22293 10084
rect 22327 10112 22339 10115
rect 23109 10115 23167 10121
rect 23109 10112 23121 10115
rect 22327 10084 23121 10112
rect 22327 10081 22339 10084
rect 22281 10075 22339 10081
rect 23109 10081 23121 10084
rect 23155 10081 23167 10115
rect 23109 10075 23167 10081
rect 20220 10016 21864 10044
rect 20220 10004 20226 10016
rect 14016 9948 14780 9976
rect 17313 9979 17371 9985
rect 17313 9945 17325 9979
rect 17359 9976 17371 9979
rect 17862 9976 17868 9988
rect 17359 9948 17868 9976
rect 17359 9945 17371 9948
rect 17313 9939 17371 9945
rect 17862 9936 17868 9948
rect 17920 9936 17926 9988
rect 20349 9979 20407 9985
rect 20349 9945 20361 9979
rect 20395 9945 20407 9979
rect 23124 9976 23152 10075
rect 23290 10072 23296 10124
rect 23348 10072 23354 10124
rect 23382 10072 23388 10124
rect 23440 10112 23446 10124
rect 23750 10112 23756 10124
rect 23440 10084 23756 10112
rect 23440 10072 23446 10084
rect 23750 10072 23756 10084
rect 23808 10072 23814 10124
rect 24105 10121 24133 10140
rect 24053 10115 24133 10121
rect 24053 10081 24065 10115
rect 24099 10084 24133 10115
rect 24213 10115 24271 10121
rect 24099 10081 24111 10084
rect 24053 10075 24111 10081
rect 24213 10081 24225 10115
rect 24259 10081 24271 10115
rect 24213 10075 24271 10081
rect 24228 10044 24256 10075
rect 24302 10072 24308 10124
rect 24360 10072 24366 10124
rect 24394 10072 24400 10124
rect 24452 10072 24458 10124
rect 24780 10121 24808 10152
rect 24765 10115 24823 10121
rect 24765 10081 24777 10115
rect 24811 10081 24823 10115
rect 24765 10075 24823 10081
rect 24949 10115 25007 10121
rect 24949 10081 24961 10115
rect 24995 10081 25007 10115
rect 24949 10075 25007 10081
rect 24854 10044 24860 10056
rect 24228 10016 24860 10044
rect 24854 10004 24860 10016
rect 24912 10004 24918 10056
rect 24964 10044 24992 10075
rect 25038 10072 25044 10124
rect 25096 10072 25102 10124
rect 25130 10072 25136 10124
rect 25188 10072 25194 10124
rect 25222 10072 25228 10124
rect 25280 10112 25286 10124
rect 25685 10115 25743 10121
rect 25685 10112 25697 10115
rect 25280 10084 25697 10112
rect 25280 10072 25286 10084
rect 25685 10081 25697 10084
rect 25731 10081 25743 10115
rect 25685 10075 25743 10081
rect 25866 10072 25872 10124
rect 25924 10072 25930 10124
rect 25961 10115 26019 10121
rect 25961 10081 25973 10115
rect 26007 10081 26019 10115
rect 25961 10075 26019 10081
rect 25501 10047 25559 10053
rect 25501 10044 25513 10047
rect 24964 10016 25513 10044
rect 25501 10013 25513 10016
rect 25547 10013 25559 10047
rect 25501 10007 25559 10013
rect 24486 9976 24492 9988
rect 23124 9948 24492 9976
rect 20349 9939 20407 9945
rect 10459 9880 13952 9908
rect 10459 9877 10471 9880
rect 10413 9871 10471 9877
rect 15470 9868 15476 9920
rect 15528 9908 15534 9920
rect 16117 9911 16175 9917
rect 16117 9908 16129 9911
rect 15528 9880 16129 9908
rect 15528 9868 15534 9880
rect 16117 9877 16129 9880
rect 16163 9877 16175 9911
rect 16117 9871 16175 9877
rect 17034 9868 17040 9920
rect 17092 9908 17098 9920
rect 17405 9911 17463 9917
rect 17405 9908 17417 9911
rect 17092 9880 17417 9908
rect 17092 9868 17098 9880
rect 17405 9877 17417 9880
rect 17451 9877 17463 9911
rect 17405 9871 17463 9877
rect 19518 9868 19524 9920
rect 19576 9908 19582 9920
rect 20364 9908 20392 9939
rect 24486 9936 24492 9948
rect 24544 9936 24550 9988
rect 24670 9936 24676 9988
rect 24728 9936 24734 9988
rect 24946 9936 24952 9988
rect 25004 9976 25010 9988
rect 25976 9976 26004 10075
rect 26418 10072 26424 10124
rect 26476 10112 26482 10124
rect 26973 10115 27031 10121
rect 26973 10112 26985 10115
rect 26476 10084 26985 10112
rect 26476 10072 26482 10084
rect 26973 10081 26985 10084
rect 27019 10081 27031 10115
rect 26973 10075 27031 10081
rect 25004 9948 26004 9976
rect 25004 9936 25010 9948
rect 26418 9936 26424 9988
rect 26476 9936 26482 9988
rect 19576 9880 20392 9908
rect 19576 9868 19582 9880
rect 24302 9868 24308 9920
rect 24360 9908 24366 9920
rect 25038 9908 25044 9920
rect 24360 9880 25044 9908
rect 24360 9868 24366 9880
rect 25038 9868 25044 9880
rect 25096 9868 25102 9920
rect 552 9818 27416 9840
rect 552 9766 3756 9818
rect 3808 9766 3820 9818
rect 3872 9766 3884 9818
rect 3936 9766 3948 9818
rect 4000 9766 4012 9818
rect 4064 9766 10472 9818
rect 10524 9766 10536 9818
rect 10588 9766 10600 9818
rect 10652 9766 10664 9818
rect 10716 9766 10728 9818
rect 10780 9766 17188 9818
rect 17240 9766 17252 9818
rect 17304 9766 17316 9818
rect 17368 9766 17380 9818
rect 17432 9766 17444 9818
rect 17496 9766 23904 9818
rect 23956 9766 23968 9818
rect 24020 9766 24032 9818
rect 24084 9766 24096 9818
rect 24148 9766 24160 9818
rect 24212 9766 27416 9818
rect 552 9744 27416 9766
rect 5629 9707 5687 9713
rect 5629 9673 5641 9707
rect 5675 9704 5687 9707
rect 6362 9704 6368 9716
rect 5675 9676 6368 9704
rect 5675 9673 5687 9676
rect 5629 9667 5687 9673
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 13446 9664 13452 9716
rect 13504 9704 13510 9716
rect 16022 9704 16028 9716
rect 13504 9676 16028 9704
rect 13504 9664 13510 9676
rect 16022 9664 16028 9676
rect 16080 9664 16086 9716
rect 16500 9676 17724 9704
rect 2777 9639 2835 9645
rect 2777 9605 2789 9639
rect 2823 9605 2835 9639
rect 2777 9599 2835 9605
rect 2792 9568 2820 9599
rect 2866 9596 2872 9648
rect 2924 9596 2930 9648
rect 3602 9596 3608 9648
rect 3660 9636 3666 9648
rect 3973 9639 4031 9645
rect 3973 9636 3985 9639
rect 3660 9608 3985 9636
rect 3660 9596 3666 9608
rect 3973 9605 3985 9608
rect 4019 9605 4031 9639
rect 3973 9599 4031 9605
rect 4080 9608 5304 9636
rect 3789 9571 3847 9577
rect 3789 9568 3801 9571
rect 2792 9540 3801 9568
rect 3620 9512 3648 9540
rect 3789 9537 3801 9540
rect 3835 9568 3847 9571
rect 4080 9568 4108 9608
rect 5276 9577 5304 9608
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 6089 9639 6147 9645
rect 6089 9636 6101 9639
rect 5592 9608 6101 9636
rect 5592 9596 5598 9608
rect 6089 9605 6101 9608
rect 6135 9605 6147 9639
rect 9306 9636 9312 9648
rect 6089 9599 6147 9605
rect 9140 9608 9312 9636
rect 4893 9571 4951 9577
rect 4893 9568 4905 9571
rect 3835 9540 4108 9568
rect 4172 9540 4905 9568
rect 3835 9537 3847 9540
rect 3789 9531 3847 9537
rect 4172 9512 4200 9540
rect 4893 9537 4905 9540
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 5626 9528 5632 9580
rect 5684 9568 5690 9580
rect 5721 9571 5779 9577
rect 5721 9568 5733 9571
rect 5684 9540 5733 9568
rect 5684 9528 5690 9540
rect 5721 9537 5733 9540
rect 5767 9537 5779 9571
rect 6822 9568 6828 9580
rect 5721 9531 5779 9537
rect 6196 9540 6828 9568
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 2406 9500 2412 9512
rect 1443 9472 2412 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 3050 9460 3056 9512
rect 3108 9460 3114 9512
rect 3602 9460 3608 9512
rect 3660 9460 3666 9512
rect 4154 9460 4160 9512
rect 4212 9460 4218 9512
rect 4430 9460 4436 9512
rect 4488 9460 4494 9512
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9469 4767 9503
rect 4709 9463 4767 9469
rect 1670 9441 1676 9444
rect 1664 9395 1676 9441
rect 1670 9392 1676 9395
rect 1728 9392 1734 9444
rect 3142 9392 3148 9444
rect 3200 9432 3206 9444
rect 4341 9435 4399 9441
rect 4341 9432 4353 9435
rect 3200 9404 4353 9432
rect 3200 9392 3206 9404
rect 4341 9401 4353 9404
rect 4387 9432 4399 9435
rect 4724 9432 4752 9463
rect 5442 9460 5448 9512
rect 5500 9460 5506 9512
rect 5905 9503 5963 9509
rect 5905 9469 5917 9503
rect 5951 9469 5963 9503
rect 5905 9463 5963 9469
rect 4982 9432 4988 9444
rect 4387 9404 4988 9432
rect 4387 9401 4399 9404
rect 4341 9395 4399 9401
rect 4982 9392 4988 9404
rect 5040 9392 5046 9444
rect 5460 9432 5488 9460
rect 5718 9432 5724 9444
rect 5460 9404 5724 9432
rect 5718 9392 5724 9404
rect 5776 9392 5782 9444
rect 5920 9432 5948 9463
rect 5994 9460 6000 9512
rect 6052 9460 6058 9512
rect 6196 9509 6224 9540
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9469 6239 9503
rect 6181 9463 6239 9469
rect 6270 9460 6276 9512
rect 6328 9500 6334 9512
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 6328 9472 6377 9500
rect 6328 9460 6334 9472
rect 6365 9469 6377 9472
rect 6411 9500 6423 9503
rect 6638 9500 6644 9512
rect 6411 9472 6644 9500
rect 6411 9469 6423 9472
rect 6365 9463 6423 9469
rect 6638 9460 6644 9472
rect 6696 9460 6702 9512
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9500 7711 9503
rect 8110 9500 8116 9512
rect 7699 9472 8116 9500
rect 7699 9469 7711 9472
rect 7653 9463 7711 9469
rect 8110 9460 8116 9472
rect 8168 9460 8174 9512
rect 8754 9460 8760 9512
rect 8812 9500 8818 9512
rect 9140 9509 9168 9608
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 14458 9596 14464 9648
rect 14516 9596 14522 9648
rect 15746 9596 15752 9648
rect 15804 9636 15810 9648
rect 16500 9636 16528 9676
rect 15804 9608 16528 9636
rect 15804 9596 15810 9608
rect 11514 9528 11520 9580
rect 11572 9568 11578 9580
rect 11609 9571 11667 9577
rect 11609 9568 11621 9571
rect 11572 9540 11621 9568
rect 11572 9528 11578 9540
rect 11609 9537 11621 9540
rect 11655 9537 11667 9571
rect 11609 9531 11667 9537
rect 15286 9528 15292 9580
rect 15344 9568 15350 9580
rect 15344 9540 16252 9568
rect 15344 9528 15350 9540
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 8812 9472 8953 9500
rect 8812 9460 8818 9472
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 6086 9432 6092 9444
rect 5920 9404 6092 9432
rect 6086 9392 6092 9404
rect 6144 9432 6150 9444
rect 6730 9432 6736 9444
rect 6144 9404 6736 9432
rect 6144 9392 6150 9404
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 8956 9432 8984 9463
rect 9214 9460 9220 9512
rect 9272 9460 9278 9512
rect 9309 9503 9367 9509
rect 9309 9469 9321 9503
rect 9355 9500 9367 9503
rect 9490 9500 9496 9512
rect 9355 9472 9496 9500
rect 9355 9469 9367 9472
rect 9309 9463 9367 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 9582 9460 9588 9512
rect 9640 9500 9646 9512
rect 9677 9503 9735 9509
rect 9677 9500 9689 9503
rect 9640 9472 9689 9500
rect 9640 9460 9646 9472
rect 9677 9469 9689 9472
rect 9723 9500 9735 9503
rect 11532 9500 11560 9528
rect 9723 9472 11560 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 12986 9460 12992 9512
rect 13044 9500 13050 9512
rect 13170 9500 13176 9512
rect 13044 9472 13176 9500
rect 13044 9460 13050 9472
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 16114 9460 16120 9512
rect 16172 9460 16178 9512
rect 16224 9509 16252 9540
rect 16500 9509 16528 9608
rect 16574 9596 16580 9648
rect 16632 9636 16638 9648
rect 16669 9639 16727 9645
rect 16669 9636 16681 9639
rect 16632 9608 16681 9636
rect 16632 9596 16638 9608
rect 16669 9605 16681 9608
rect 16715 9605 16727 9639
rect 17586 9636 17592 9648
rect 16669 9599 16727 9605
rect 17052 9608 17592 9636
rect 16942 9528 16948 9580
rect 17000 9528 17006 9580
rect 17052 9577 17080 9608
rect 17586 9596 17592 9608
rect 17644 9596 17650 9648
rect 17696 9636 17724 9676
rect 18230 9664 18236 9716
rect 18288 9704 18294 9716
rect 18969 9707 19027 9713
rect 18969 9704 18981 9707
rect 18288 9676 18981 9704
rect 18288 9664 18294 9676
rect 18969 9673 18981 9676
rect 19015 9673 19027 9707
rect 18969 9667 19027 9673
rect 22370 9664 22376 9716
rect 22428 9704 22434 9716
rect 22428 9676 23336 9704
rect 22428 9664 22434 9676
rect 18598 9636 18604 9648
rect 17696 9608 18604 9636
rect 18598 9596 18604 9608
rect 18656 9636 18662 9648
rect 18656 9608 19656 9636
rect 18656 9596 18662 9608
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 17218 9528 17224 9580
rect 17276 9568 17282 9580
rect 17313 9571 17371 9577
rect 17313 9568 17325 9571
rect 17276 9540 17325 9568
rect 17276 9528 17282 9540
rect 17313 9537 17325 9540
rect 17359 9537 17371 9571
rect 17313 9531 17371 9537
rect 17494 9528 17500 9580
rect 17552 9528 17558 9580
rect 19518 9568 19524 9580
rect 19260 9540 19524 9568
rect 16209 9503 16267 9509
rect 16209 9469 16221 9503
rect 16255 9469 16267 9503
rect 16209 9463 16267 9469
rect 16301 9503 16359 9509
rect 16301 9469 16313 9503
rect 16347 9469 16359 9503
rect 16301 9463 16359 9469
rect 16485 9503 16543 9509
rect 16485 9469 16497 9503
rect 16531 9469 16543 9503
rect 16485 9463 16543 9469
rect 9398 9432 9404 9444
rect 8956 9404 9404 9432
rect 9398 9392 9404 9404
rect 9456 9392 9462 9444
rect 11882 9441 11888 9444
rect 9922 9435 9980 9441
rect 9922 9432 9934 9435
rect 9600 9404 9934 9432
rect 2866 9324 2872 9376
rect 2924 9364 2930 9376
rect 3237 9367 3295 9373
rect 3237 9364 3249 9367
rect 2924 9336 3249 9364
rect 2924 9324 2930 9336
rect 3237 9333 3249 9336
rect 3283 9333 3295 9367
rect 3237 9327 3295 9333
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 4614 9364 4620 9376
rect 4571 9336 4620 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 8205 9367 8263 9373
rect 8205 9333 8217 9367
rect 8251 9364 8263 9367
rect 8386 9364 8392 9376
rect 8251 9336 8392 9364
rect 8251 9333 8263 9336
rect 8205 9327 8263 9333
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 9600 9373 9628 9404
rect 9922 9401 9934 9404
rect 9968 9401 9980 9435
rect 9922 9395 9980 9401
rect 11876 9395 11888 9441
rect 11882 9392 11888 9395
rect 11940 9392 11946 9444
rect 12342 9392 12348 9444
rect 12400 9432 12406 9444
rect 13262 9432 13268 9444
rect 12400 9404 13268 9432
rect 12400 9392 12406 9404
rect 13262 9392 13268 9404
rect 13320 9392 13326 9444
rect 15746 9392 15752 9444
rect 15804 9392 15810 9444
rect 15930 9392 15936 9444
rect 15988 9432 15994 9444
rect 16316 9432 16344 9463
rect 16850 9460 16856 9512
rect 16908 9460 16914 9512
rect 17126 9460 17132 9512
rect 17184 9460 17190 9512
rect 17589 9503 17647 9509
rect 17589 9469 17601 9503
rect 17635 9500 17647 9503
rect 17954 9500 17960 9512
rect 17635 9472 17960 9500
rect 17635 9469 17647 9472
rect 17589 9463 17647 9469
rect 17954 9460 17960 9472
rect 18012 9460 18018 9512
rect 19260 9509 19288 9540
rect 19518 9528 19524 9540
rect 19576 9528 19582 9580
rect 19628 9568 19656 9608
rect 20438 9596 20444 9648
rect 20496 9636 20502 9648
rect 20533 9639 20591 9645
rect 20533 9636 20545 9639
rect 20496 9608 20545 9636
rect 20496 9596 20502 9608
rect 20533 9605 20545 9608
rect 20579 9605 20591 9639
rect 20533 9599 20591 9605
rect 21358 9596 21364 9648
rect 21416 9636 21422 9648
rect 21634 9636 21640 9648
rect 21416 9608 21640 9636
rect 21416 9596 21422 9608
rect 21634 9596 21640 9608
rect 21692 9596 21698 9648
rect 20456 9568 20484 9596
rect 19628 9540 20484 9568
rect 19245 9503 19303 9509
rect 19245 9469 19257 9503
rect 19291 9469 19303 9503
rect 19245 9463 19303 9469
rect 19334 9460 19340 9512
rect 19392 9460 19398 9512
rect 19628 9509 19656 9540
rect 22738 9528 22744 9580
rect 22796 9528 22802 9580
rect 23308 9577 23336 9676
rect 24673 9639 24731 9645
rect 24673 9605 24685 9639
rect 24719 9636 24731 9639
rect 24762 9636 24768 9648
rect 24719 9608 24768 9636
rect 24719 9605 24731 9608
rect 24673 9599 24731 9605
rect 24762 9596 24768 9608
rect 24820 9596 24826 9648
rect 24854 9596 24860 9648
rect 24912 9596 24918 9648
rect 23201 9571 23259 9577
rect 23201 9568 23213 9571
rect 22940 9540 23213 9568
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9469 19487 9503
rect 19429 9463 19487 9469
rect 19613 9503 19671 9509
rect 19613 9469 19625 9503
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 15988 9404 16344 9432
rect 16868 9432 16896 9460
rect 17494 9432 17500 9444
rect 16868 9404 17500 9432
rect 15988 9392 15994 9404
rect 17494 9392 17500 9404
rect 17552 9392 17558 9444
rect 19444 9432 19472 9463
rect 19886 9460 19892 9512
rect 19944 9460 19950 9512
rect 20162 9500 20168 9512
rect 19996 9472 20168 9500
rect 19705 9435 19763 9441
rect 19705 9432 19717 9435
rect 19444 9404 19717 9432
rect 19705 9401 19717 9404
rect 19751 9401 19763 9435
rect 19705 9395 19763 9401
rect 9585 9367 9643 9373
rect 9585 9333 9597 9367
rect 9631 9333 9643 9367
rect 9585 9327 9643 9333
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 11057 9367 11115 9373
rect 11057 9364 11069 9367
rect 9732 9336 11069 9364
rect 9732 9324 9738 9336
rect 11057 9333 11069 9336
rect 11103 9364 11115 9367
rect 12434 9364 12440 9376
rect 11103 9336 12440 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 12989 9367 13047 9373
rect 12989 9333 13001 9367
rect 13035 9364 13047 9367
rect 13170 9364 13176 9376
rect 13035 9336 13176 9364
rect 13035 9333 13047 9336
rect 12989 9327 13047 9333
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 15841 9367 15899 9373
rect 15841 9333 15853 9367
rect 15887 9364 15899 9367
rect 16022 9364 16028 9376
rect 15887 9336 16028 9364
rect 15887 9333 15899 9336
rect 15841 9327 15899 9333
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 17313 9367 17371 9373
rect 17313 9364 17325 9367
rect 17092 9336 17325 9364
rect 17092 9324 17098 9336
rect 17313 9333 17325 9336
rect 17359 9333 17371 9367
rect 17313 9327 17371 9333
rect 18046 9324 18052 9376
rect 18104 9364 18110 9376
rect 19996 9364 20024 9472
rect 20162 9460 20168 9472
rect 20220 9460 20226 9512
rect 20349 9503 20407 9509
rect 20349 9469 20361 9503
rect 20395 9500 20407 9503
rect 21174 9500 21180 9512
rect 20395 9472 21180 9500
rect 20395 9469 20407 9472
rect 20349 9463 20407 9469
rect 21174 9460 21180 9472
rect 21232 9460 21238 9512
rect 22094 9460 22100 9512
rect 22152 9500 22158 9512
rect 22940 9500 22968 9540
rect 23201 9537 23213 9540
rect 23247 9537 23259 9571
rect 23201 9531 23259 9537
rect 23293 9571 23351 9577
rect 23293 9537 23305 9571
rect 23339 9537 23351 9571
rect 24946 9568 24952 9580
rect 23293 9531 23351 9537
rect 24228 9540 24952 9568
rect 22152 9472 22968 9500
rect 23017 9503 23075 9509
rect 22152 9460 22158 9472
rect 23017 9469 23029 9503
rect 23063 9469 23075 9503
rect 23017 9463 23075 9469
rect 23109 9503 23167 9509
rect 23109 9469 23121 9503
rect 23155 9500 23167 9503
rect 23382 9500 23388 9512
rect 23155 9472 23388 9500
rect 23155 9469 23167 9472
rect 23109 9463 23167 9469
rect 22186 9392 22192 9444
rect 22244 9432 22250 9444
rect 22474 9435 22532 9441
rect 22474 9432 22486 9435
rect 22244 9404 22486 9432
rect 22244 9392 22250 9404
rect 22474 9401 22486 9404
rect 22520 9401 22532 9435
rect 23032 9432 23060 9463
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 23750 9460 23756 9512
rect 23808 9500 23814 9512
rect 24228 9509 24256 9540
rect 24946 9528 24952 9540
rect 25004 9568 25010 9580
rect 25004 9540 25360 9568
rect 25004 9528 25010 9540
rect 24213 9503 24271 9509
rect 24213 9500 24225 9503
rect 23808 9472 24225 9500
rect 23808 9460 23814 9472
rect 24213 9469 24225 9472
rect 24259 9469 24271 9503
rect 24213 9463 24271 9469
rect 24486 9460 24492 9512
rect 24544 9500 24550 9512
rect 25041 9503 25099 9509
rect 25041 9500 25053 9503
rect 24544 9472 25053 9500
rect 24544 9460 24550 9472
rect 25041 9469 25053 9472
rect 25087 9500 25099 9503
rect 25222 9500 25228 9512
rect 25087 9472 25228 9500
rect 25087 9469 25099 9472
rect 25041 9463 25099 9469
rect 25222 9460 25228 9472
rect 25280 9460 25286 9512
rect 25332 9509 25360 9540
rect 25317 9503 25375 9509
rect 25317 9469 25329 9503
rect 25363 9469 25375 9503
rect 25317 9463 25375 9469
rect 23290 9432 23296 9444
rect 23032 9404 23296 9432
rect 22474 9395 22532 9401
rect 23290 9392 23296 9404
rect 23348 9392 23354 9444
rect 18104 9336 20024 9364
rect 20073 9367 20131 9373
rect 18104 9324 18110 9336
rect 20073 9333 20085 9367
rect 20119 9364 20131 9367
rect 20438 9364 20444 9376
rect 20119 9336 20444 9364
rect 20119 9333 20131 9336
rect 20073 9327 20131 9333
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 21174 9324 21180 9376
rect 21232 9364 21238 9376
rect 22278 9364 22284 9376
rect 21232 9336 22284 9364
rect 21232 9324 21238 9336
rect 22278 9324 22284 9336
rect 22336 9324 22342 9376
rect 22738 9324 22744 9376
rect 22796 9364 22802 9376
rect 22833 9367 22891 9373
rect 22833 9364 22845 9367
rect 22796 9336 22845 9364
rect 22796 9324 22802 9336
rect 22833 9333 22845 9336
rect 22879 9333 22891 9367
rect 22833 9327 22891 9333
rect 24305 9367 24363 9373
rect 24305 9333 24317 9367
rect 24351 9364 24363 9367
rect 24486 9364 24492 9376
rect 24351 9336 24492 9364
rect 24351 9333 24363 9336
rect 24305 9327 24363 9333
rect 24486 9324 24492 9336
rect 24544 9324 24550 9376
rect 24946 9324 24952 9376
rect 25004 9364 25010 9376
rect 25225 9367 25283 9373
rect 25225 9364 25237 9367
rect 25004 9336 25237 9364
rect 25004 9324 25010 9336
rect 25225 9333 25237 9336
rect 25271 9333 25283 9367
rect 25225 9327 25283 9333
rect 552 9274 27576 9296
rect 552 9222 7114 9274
rect 7166 9222 7178 9274
rect 7230 9222 7242 9274
rect 7294 9222 7306 9274
rect 7358 9222 7370 9274
rect 7422 9222 13830 9274
rect 13882 9222 13894 9274
rect 13946 9222 13958 9274
rect 14010 9222 14022 9274
rect 14074 9222 14086 9274
rect 14138 9222 20546 9274
rect 20598 9222 20610 9274
rect 20662 9222 20674 9274
rect 20726 9222 20738 9274
rect 20790 9222 20802 9274
rect 20854 9222 27262 9274
rect 27314 9222 27326 9274
rect 27378 9222 27390 9274
rect 27442 9222 27454 9274
rect 27506 9222 27518 9274
rect 27570 9222 27576 9274
rect 552 9200 27576 9222
rect 1670 9120 1676 9172
rect 1728 9169 1734 9172
rect 1728 9160 1737 9169
rect 1728 9132 1773 9160
rect 1728 9123 1737 9132
rect 1728 9120 1734 9123
rect 2038 9120 2044 9172
rect 2096 9160 2102 9172
rect 4433 9163 4491 9169
rect 4433 9160 4445 9163
rect 2096 9132 4445 9160
rect 2096 9120 2102 9132
rect 4433 9129 4445 9132
rect 4479 9129 4491 9163
rect 4433 9123 4491 9129
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 8110 9120 8116 9172
rect 8168 9120 8174 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8754 9160 8760 9172
rect 8352 9132 8760 9160
rect 8352 9120 8358 9132
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 8904 9132 9168 9160
rect 8904 9120 8910 9132
rect 1765 9095 1823 9101
rect 1765 9061 1777 9095
rect 1811 9092 1823 9095
rect 1811 9064 1992 9092
rect 1811 9061 1823 9064
rect 1765 9055 1823 9061
rect 1581 9027 1639 9033
rect 1581 8993 1593 9027
rect 1627 8993 1639 9027
rect 1581 8987 1639 8993
rect 1596 8956 1624 8987
rect 1854 8984 1860 9036
rect 1912 8984 1918 9036
rect 1964 9033 1992 9064
rect 5166 9052 5172 9104
rect 5224 9052 5230 9104
rect 8386 9052 8392 9104
rect 8444 9092 8450 9104
rect 9033 9095 9091 9101
rect 9033 9092 9045 9095
rect 8444 9064 9045 9092
rect 8444 9052 8450 9064
rect 9033 9061 9045 9064
rect 9079 9061 9091 9095
rect 9033 9055 9091 9061
rect 9140 9092 9168 9132
rect 9306 9120 9312 9172
rect 9364 9120 9370 9172
rect 11882 9120 11888 9172
rect 11940 9120 11946 9172
rect 12158 9120 12164 9172
rect 12216 9160 12222 9172
rect 12621 9163 12679 9169
rect 12621 9160 12633 9163
rect 12216 9132 12633 9160
rect 12216 9120 12222 9132
rect 12621 9129 12633 9132
rect 12667 9129 12679 9163
rect 12621 9123 12679 9129
rect 14274 9120 14280 9172
rect 14332 9160 14338 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 14332 9132 14381 9160
rect 14332 9120 14338 9132
rect 14369 9129 14381 9132
rect 14415 9129 14427 9163
rect 14369 9123 14427 9129
rect 17770 9120 17776 9172
rect 17828 9160 17834 9172
rect 17865 9163 17923 9169
rect 17865 9160 17877 9163
rect 17828 9132 17877 9160
rect 17828 9120 17834 9132
rect 17865 9129 17877 9132
rect 17911 9129 17923 9163
rect 17865 9123 17923 9129
rect 9766 9092 9772 9104
rect 9140 9064 9772 9092
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 9024 2007 9027
rect 2866 9024 2872 9036
rect 1995 8996 2872 9024
rect 1995 8993 2007 8996
rect 1949 8987 2007 8993
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 2961 9027 3019 9033
rect 2961 8993 2973 9027
rect 3007 9024 3019 9027
rect 3881 9027 3939 9033
rect 3881 9024 3893 9027
rect 3007 8996 3893 9024
rect 3007 8993 3019 8996
rect 2961 8987 3019 8993
rect 3881 8993 3893 8996
rect 3927 8993 3939 9027
rect 3881 8987 3939 8993
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 9024 4123 9027
rect 4111 8996 4568 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 2225 8959 2283 8965
rect 1596 8928 2176 8956
rect 2038 8848 2044 8900
rect 2096 8848 2102 8900
rect 2148 8897 2176 8928
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2314 8956 2320 8968
rect 2271 8928 2320 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 3142 8916 3148 8968
rect 3200 8916 3206 8968
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8956 3847 8959
rect 4341 8959 4399 8965
rect 4341 8956 4353 8959
rect 3835 8928 4353 8956
rect 3835 8925 3847 8928
rect 3789 8919 3847 8925
rect 4341 8925 4353 8928
rect 4387 8925 4399 8959
rect 4341 8919 4399 8925
rect 2133 8891 2191 8897
rect 2133 8857 2145 8891
rect 2179 8857 2191 8891
rect 4540 8888 4568 8996
rect 4614 8984 4620 9036
rect 4672 8984 4678 9036
rect 4893 9027 4951 9033
rect 4893 9024 4905 9027
rect 4816 8996 4905 9024
rect 4816 8968 4844 8996
rect 4893 8993 4905 8996
rect 4939 8993 4951 9027
rect 4893 8987 4951 8993
rect 5810 8984 5816 9036
rect 5868 9024 5874 9036
rect 7006 9033 7012 9036
rect 6733 9027 6791 9033
rect 6733 9024 6745 9027
rect 5868 8996 6745 9024
rect 5868 8984 5874 8996
rect 6733 8993 6745 8996
rect 6779 8993 6791 9027
rect 6733 8987 6791 8993
rect 7000 8987 7012 9033
rect 7006 8984 7012 8987
rect 7064 8984 7070 9036
rect 8573 9027 8631 9033
rect 8573 8993 8585 9027
rect 8619 8993 8631 9027
rect 8573 8987 8631 8993
rect 8665 9027 8723 9033
rect 8665 8993 8677 9027
rect 8711 8993 8723 9027
rect 8665 8987 8723 8993
rect 8758 9027 8816 9033
rect 8758 8993 8770 9027
rect 8804 9024 8816 9027
rect 8804 8996 8892 9024
rect 8804 8993 8816 8996
rect 8758 8987 8816 8993
rect 4798 8916 4804 8968
rect 4856 8916 4862 8968
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 8588 8956 8616 8987
rect 8260 8928 8616 8956
rect 8260 8916 8266 8928
rect 5169 8891 5227 8897
rect 5169 8888 5181 8891
rect 4540 8860 5181 8888
rect 2133 8851 2191 8857
rect 5169 8857 5181 8860
rect 5215 8857 5227 8891
rect 5169 8851 5227 8857
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 2317 8823 2375 8829
rect 2317 8820 2329 8823
rect 2280 8792 2329 8820
rect 2280 8780 2286 8792
rect 2317 8789 2329 8792
rect 2363 8789 2375 8823
rect 2317 8783 2375 8789
rect 4249 8823 4307 8829
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 4430 8820 4436 8832
rect 4295 8792 4436 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 4430 8780 4436 8792
rect 4488 8820 4494 8832
rect 4798 8820 4804 8832
rect 4488 8792 4804 8820
rect 4488 8780 4494 8792
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 7466 8780 7472 8832
rect 7524 8820 7530 8832
rect 8205 8823 8263 8829
rect 8205 8820 8217 8823
rect 7524 8792 8217 8820
rect 7524 8780 7530 8792
rect 8205 8789 8217 8792
rect 8251 8789 8263 8823
rect 8588 8820 8616 8928
rect 8680 8888 8708 8987
rect 8754 8888 8760 8900
rect 8680 8860 8760 8888
rect 8754 8848 8760 8860
rect 8812 8848 8818 8900
rect 8864 8888 8892 8996
rect 8938 8984 8944 9036
rect 8996 8984 9002 9036
rect 9140 9033 9168 9064
rect 9766 9052 9772 9064
rect 9824 9052 9830 9104
rect 10962 9052 10968 9104
rect 11020 9092 11026 9104
rect 11020 9064 13124 9092
rect 11020 9052 11026 9064
rect 9130 9027 9188 9033
rect 9130 8993 9142 9027
rect 9176 8993 9188 9027
rect 9130 8987 9188 8993
rect 9306 8984 9312 9036
rect 9364 9024 9370 9036
rect 11330 9024 11336 9036
rect 9364 8996 11336 9024
rect 9364 8984 9370 8996
rect 11330 8984 11336 8996
rect 11388 9024 11394 9036
rect 12342 9024 12348 9036
rect 11388 8996 12348 9024
rect 11388 8984 11394 8996
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 11882 8916 11888 8968
rect 11940 8956 11946 8968
rect 12437 8959 12495 8965
rect 12437 8956 12449 8959
rect 11940 8928 12449 8956
rect 11940 8916 11946 8928
rect 12437 8925 12449 8928
rect 12483 8925 12495 8959
rect 13096 8956 13124 9064
rect 13262 9052 13268 9104
rect 13320 9092 13326 9104
rect 13320 9064 14044 9092
rect 13320 9052 13326 9064
rect 13170 8984 13176 9036
rect 13228 8984 13234 9036
rect 13538 9033 13544 9036
rect 13536 9024 13544 9033
rect 13499 8996 13544 9024
rect 13536 8987 13544 8996
rect 13538 8984 13544 8987
rect 13596 8984 13602 9036
rect 13630 8984 13636 9036
rect 13688 8984 13694 9036
rect 14016 9033 14044 9064
rect 15470 9052 15476 9104
rect 15528 9101 15534 9104
rect 15528 9092 15540 9101
rect 15528 9064 15573 9092
rect 15528 9055 15540 9064
rect 15528 9052 15534 9055
rect 16758 9033 16764 9036
rect 13725 9027 13783 9033
rect 13725 8993 13737 9027
rect 13771 8993 13783 9027
rect 13725 8987 13783 8993
rect 13908 9027 13966 9033
rect 13908 8993 13920 9027
rect 13954 8993 13966 9027
rect 13908 8987 13966 8993
rect 14001 9027 14059 9033
rect 14001 8993 14013 9027
rect 14047 8993 14059 9027
rect 16752 9024 16764 9033
rect 16719 8996 16764 9024
rect 14001 8987 14059 8993
rect 16752 8987 16764 8996
rect 13446 8956 13452 8968
rect 13096 8928 13452 8956
rect 12437 8919 12495 8925
rect 13446 8916 13452 8928
rect 13504 8956 13510 8968
rect 13740 8956 13768 8987
rect 13504 8928 13768 8956
rect 13924 8956 13952 8987
rect 16758 8984 16764 8987
rect 16816 8984 16822 9036
rect 17880 9024 17908 9123
rect 18782 9120 18788 9172
rect 18840 9160 18846 9172
rect 19153 9163 19211 9169
rect 19153 9160 19165 9163
rect 18840 9132 19165 9160
rect 18840 9120 18846 9132
rect 19153 9129 19165 9132
rect 19199 9129 19211 9163
rect 19153 9123 19211 9129
rect 22370 9120 22376 9172
rect 22428 9160 22434 9172
rect 22649 9163 22707 9169
rect 22649 9160 22661 9163
rect 22428 9132 22661 9160
rect 22428 9120 22434 9132
rect 22649 9129 22661 9132
rect 22695 9160 22707 9163
rect 23937 9163 23995 9169
rect 22695 9132 23704 9160
rect 22695 9129 22707 9132
rect 22649 9123 22707 9129
rect 18046 9052 18052 9104
rect 18104 9092 18110 9104
rect 19886 9092 19892 9104
rect 18104 9064 18644 9092
rect 18104 9052 18110 9064
rect 18509 9027 18567 9033
rect 18509 9024 18521 9027
rect 17880 8996 18521 9024
rect 18509 8993 18521 8996
rect 18555 8993 18567 9027
rect 18616 9024 18644 9064
rect 18984 9064 19892 9092
rect 18693 9027 18751 9033
rect 18693 9024 18705 9027
rect 18616 8996 18705 9024
rect 18509 8987 18567 8993
rect 18693 8993 18705 8996
rect 18739 8993 18751 9027
rect 18693 8987 18751 8993
rect 18782 8984 18788 9036
rect 18840 8984 18846 9036
rect 18984 9033 19012 9064
rect 19886 9052 19892 9064
rect 19944 9052 19950 9104
rect 21726 9092 21732 9104
rect 21284 9064 21732 9092
rect 18969 9027 19027 9033
rect 18969 8993 18981 9027
rect 19015 8993 19027 9027
rect 18969 8987 19027 8993
rect 19797 9027 19855 9033
rect 19797 8993 19809 9027
rect 19843 9024 19855 9027
rect 20070 9024 20076 9036
rect 19843 8996 20076 9024
rect 19843 8993 19855 8996
rect 19797 8987 19855 8993
rect 20070 8984 20076 8996
rect 20128 8984 20134 9036
rect 20898 8984 20904 9036
rect 20956 9024 20962 9036
rect 21284 9033 21312 9064
rect 21726 9052 21732 9064
rect 21784 9092 21790 9104
rect 23676 9101 23704 9132
rect 23937 9129 23949 9163
rect 23983 9129 23995 9163
rect 23937 9123 23995 9129
rect 23017 9095 23075 9101
rect 23017 9092 23029 9095
rect 21784 9064 23029 9092
rect 21784 9052 21790 9064
rect 23017 9061 23029 9064
rect 23063 9061 23075 9095
rect 23661 9095 23719 9101
rect 23017 9055 23075 9061
rect 23216 9064 23428 9092
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 20956 8996 21281 9024
rect 20956 8984 20962 8996
rect 21269 8993 21281 8996
rect 21315 8993 21327 9027
rect 21269 8987 21327 8993
rect 21453 9027 21511 9033
rect 21453 8993 21465 9027
rect 21499 8993 21511 9027
rect 21453 8987 21511 8993
rect 14274 8956 14280 8968
rect 13924 8928 14280 8956
rect 13504 8916 13510 8928
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8956 15807 8959
rect 16298 8956 16304 8968
rect 15795 8928 16304 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 16298 8916 16304 8928
rect 16356 8956 16362 8968
rect 16485 8959 16543 8965
rect 16485 8956 16497 8959
rect 16356 8928 16497 8956
rect 16356 8916 16362 8928
rect 16485 8925 16497 8928
rect 16531 8925 16543 8959
rect 16485 8919 16543 8925
rect 9030 8888 9036 8900
rect 8864 8860 9036 8888
rect 9030 8848 9036 8860
rect 9088 8848 9094 8900
rect 9398 8848 9404 8900
rect 9456 8888 9462 8900
rect 10042 8888 10048 8900
rect 9456 8860 10048 8888
rect 9456 8848 9462 8860
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 12342 8848 12348 8900
rect 12400 8888 12406 8900
rect 13357 8891 13415 8897
rect 13357 8888 13369 8891
rect 12400 8860 13369 8888
rect 12400 8848 12406 8860
rect 13357 8857 13369 8860
rect 13403 8857 13415 8891
rect 21468 8888 21496 8987
rect 22094 8984 22100 9036
rect 22152 9024 22158 9036
rect 22741 9027 22799 9033
rect 22741 9024 22753 9027
rect 22152 8996 22753 9024
rect 22152 8984 22158 8996
rect 22741 8993 22753 8996
rect 22787 8993 22799 9027
rect 22741 8987 22799 8993
rect 22833 9027 22891 9033
rect 22833 8993 22845 9027
rect 22879 9024 22891 9027
rect 23216 9024 23244 9064
rect 23400 9036 23428 9064
rect 23661 9061 23673 9095
rect 23707 9061 23719 9095
rect 23952 9092 23980 9123
rect 25142 9095 25200 9101
rect 25142 9092 25154 9095
rect 23952 9064 25154 9092
rect 23661 9055 23719 9061
rect 25142 9061 25154 9064
rect 25188 9061 25200 9095
rect 25142 9055 25200 9061
rect 25685 9095 25743 9101
rect 25685 9061 25697 9095
rect 25731 9092 25743 9095
rect 26418 9092 26424 9104
rect 25731 9064 26424 9092
rect 25731 9061 25743 9064
rect 25685 9055 25743 9061
rect 22879 8996 23244 9024
rect 22879 8993 22891 8996
rect 22833 8987 22891 8993
rect 21634 8916 21640 8968
rect 21692 8956 21698 8968
rect 22373 8959 22431 8965
rect 22373 8956 22385 8959
rect 21692 8928 22385 8956
rect 21692 8916 21698 8928
rect 22373 8925 22385 8928
rect 22419 8956 22431 8959
rect 22465 8959 22523 8965
rect 22465 8956 22477 8959
rect 22419 8928 22477 8956
rect 22419 8925 22431 8928
rect 22373 8919 22431 8925
rect 22465 8925 22477 8928
rect 22511 8925 22523 8959
rect 22756 8956 22784 8987
rect 23290 8984 23296 9036
rect 23348 8984 23354 9036
rect 23382 8984 23388 9036
rect 23440 8984 23446 9036
rect 23477 9027 23535 9033
rect 23477 8993 23489 9027
rect 23523 8993 23535 9027
rect 23477 8987 23535 8993
rect 23198 8956 23204 8968
rect 22756 8928 23204 8956
rect 22465 8919 22523 8925
rect 23198 8916 23204 8928
rect 23256 8956 23262 8968
rect 23492 8956 23520 8987
rect 23256 8928 23520 8956
rect 23256 8916 23262 8928
rect 23290 8888 23296 8900
rect 21468 8860 23296 8888
rect 13357 8851 13415 8857
rect 23290 8848 23296 8860
rect 23348 8888 23354 8900
rect 23566 8888 23572 8900
rect 23348 8860 23572 8888
rect 23348 8848 23354 8860
rect 23566 8848 23572 8860
rect 23624 8848 23630 8900
rect 23676 8888 23704 9055
rect 26418 9052 26424 9064
rect 26476 9052 26482 9104
rect 23750 8984 23756 9036
rect 23808 8984 23814 9036
rect 24302 8984 24308 9036
rect 24360 9024 24366 9036
rect 25501 9027 25559 9033
rect 25501 9024 25513 9027
rect 24360 8996 25513 9024
rect 24360 8984 24366 8996
rect 25501 8993 25513 8996
rect 25547 8993 25559 9027
rect 25501 8987 25559 8993
rect 25774 8984 25780 9036
rect 25832 8984 25838 9036
rect 26145 9027 26203 9033
rect 26145 8993 26157 9027
rect 26191 8993 26203 9027
rect 26145 8987 26203 8993
rect 25406 8916 25412 8968
rect 25464 8916 25470 8968
rect 25682 8916 25688 8968
rect 25740 8956 25746 8968
rect 26160 8956 26188 8987
rect 25740 8928 26188 8956
rect 25740 8916 25746 8928
rect 24029 8891 24087 8897
rect 24029 8888 24041 8891
rect 23676 8860 24041 8888
rect 24029 8857 24041 8860
rect 24075 8857 24087 8891
rect 25590 8888 25596 8900
rect 24029 8851 24087 8857
rect 25424 8860 25596 8888
rect 12250 8820 12256 8832
rect 8588 8792 12256 8820
rect 8205 8783 8263 8789
rect 12250 8780 12256 8792
rect 12308 8780 12314 8832
rect 17954 8780 17960 8832
rect 18012 8780 18018 8832
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 19613 8823 19671 8829
rect 19613 8820 19625 8823
rect 19576 8792 19625 8820
rect 19576 8780 19582 8792
rect 19613 8789 19625 8792
rect 19659 8789 19671 8823
rect 19613 8783 19671 8789
rect 21361 8823 21419 8829
rect 21361 8789 21373 8823
rect 21407 8820 21419 8823
rect 21634 8820 21640 8832
rect 21407 8792 21640 8820
rect 21407 8789 21419 8792
rect 21361 8783 21419 8789
rect 21634 8780 21640 8792
rect 21692 8780 21698 8832
rect 21729 8823 21787 8829
rect 21729 8789 21741 8823
rect 21775 8820 21787 8823
rect 21910 8820 21916 8832
rect 21775 8792 21916 8820
rect 21775 8789 21787 8792
rect 21729 8783 21787 8789
rect 21910 8780 21916 8792
rect 21968 8780 21974 8832
rect 23106 8780 23112 8832
rect 23164 8780 23170 8832
rect 24394 8780 24400 8832
rect 24452 8820 24458 8832
rect 25424 8820 25452 8860
rect 25590 8848 25596 8860
rect 25648 8888 25654 8900
rect 25961 8891 26019 8897
rect 25961 8888 25973 8891
rect 25648 8860 25973 8888
rect 25648 8848 25654 8860
rect 25961 8857 25973 8860
rect 26007 8857 26019 8891
rect 25961 8851 26019 8857
rect 24452 8792 25452 8820
rect 24452 8780 24458 8792
rect 25498 8780 25504 8832
rect 25556 8780 25562 8832
rect 552 8730 27416 8752
rect 552 8678 3756 8730
rect 3808 8678 3820 8730
rect 3872 8678 3884 8730
rect 3936 8678 3948 8730
rect 4000 8678 4012 8730
rect 4064 8678 10472 8730
rect 10524 8678 10536 8730
rect 10588 8678 10600 8730
rect 10652 8678 10664 8730
rect 10716 8678 10728 8730
rect 10780 8678 17188 8730
rect 17240 8678 17252 8730
rect 17304 8678 17316 8730
rect 17368 8678 17380 8730
rect 17432 8678 17444 8730
rect 17496 8678 23904 8730
rect 23956 8678 23968 8730
rect 24020 8678 24032 8730
rect 24084 8678 24096 8730
rect 24148 8678 24160 8730
rect 24212 8678 27416 8730
rect 552 8656 27416 8678
rect 2961 8619 3019 8625
rect 2961 8585 2973 8619
rect 3007 8616 3019 8619
rect 3142 8616 3148 8628
rect 3007 8588 3148 8616
rect 3007 8585 3019 8588
rect 2961 8579 3019 8585
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 7006 8576 7012 8628
rect 7064 8576 7070 8628
rect 8662 8576 8668 8628
rect 8720 8616 8726 8628
rect 9030 8616 9036 8628
rect 8720 8588 9036 8616
rect 8720 8576 8726 8588
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 10962 8616 10968 8628
rect 9600 8588 10968 8616
rect 9600 8560 9628 8588
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 12618 8616 12624 8628
rect 11440 8588 12624 8616
rect 4338 8548 4344 8560
rect 3712 8520 4344 8548
rect 1486 8372 1492 8424
rect 1544 8412 1550 8424
rect 1581 8415 1639 8421
rect 1581 8412 1593 8415
rect 1544 8384 1593 8412
rect 1544 8372 1550 8384
rect 1581 8381 1593 8384
rect 1627 8412 1639 8415
rect 2682 8412 2688 8424
rect 1627 8384 2688 8412
rect 1627 8381 1639 8384
rect 1581 8375 1639 8381
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 3712 8421 3740 8520
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 8938 8508 8944 8560
rect 8996 8548 9002 8560
rect 9582 8548 9588 8560
rect 8996 8520 9588 8548
rect 8996 8508 9002 8520
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 9766 8508 9772 8560
rect 9824 8548 9830 8560
rect 11440 8548 11468 8588
rect 12618 8576 12624 8588
rect 12676 8616 12682 8628
rect 13538 8616 13544 8628
rect 12676 8588 13544 8616
rect 12676 8576 12682 8588
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 13630 8576 13636 8628
rect 13688 8616 13694 8628
rect 14921 8619 14979 8625
rect 14921 8616 14933 8619
rect 13688 8588 14933 8616
rect 13688 8576 13694 8588
rect 14921 8585 14933 8588
rect 14967 8585 14979 8619
rect 14921 8579 14979 8585
rect 9824 8520 11468 8548
rect 9824 8508 9830 8520
rect 3786 8440 3792 8492
rect 3844 8480 3850 8492
rect 4430 8480 4436 8492
rect 3844 8452 4436 8480
rect 3844 8440 3850 8452
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 10410 8480 10416 8492
rect 9272 8452 10416 8480
rect 9272 8440 9278 8452
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 11330 8480 11336 8492
rect 11164 8452 11336 8480
rect 3605 8415 3663 8421
rect 3605 8381 3617 8415
rect 3651 8381 3663 8415
rect 3605 8375 3663 8381
rect 3697 8415 3755 8421
rect 3697 8381 3709 8415
rect 3743 8381 3755 8415
rect 3697 8375 3755 8381
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8412 3939 8415
rect 4062 8412 4068 8424
rect 3927 8384 4068 8412
rect 3927 8381 3939 8384
rect 3881 8375 3939 8381
rect 1848 8347 1906 8353
rect 1848 8313 1860 8347
rect 1894 8344 1906 8347
rect 2222 8344 2228 8356
rect 1894 8316 2228 8344
rect 1894 8313 1906 8316
rect 1848 8307 1906 8313
rect 2222 8304 2228 8316
rect 2280 8304 2286 8356
rect 3620 8344 3648 8375
rect 4062 8372 4068 8384
rect 4120 8412 4126 8424
rect 4617 8415 4675 8421
rect 4617 8412 4629 8415
rect 4120 8384 4629 8412
rect 4120 8372 4126 8384
rect 4617 8381 4629 8384
rect 4663 8412 4675 8415
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 4663 8384 5549 8412
rect 4663 8381 4675 8384
rect 4617 8375 4675 8381
rect 5537 8381 5549 8384
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 5718 8372 5724 8424
rect 5776 8372 5782 8424
rect 7558 8372 7564 8424
rect 7616 8372 7622 8424
rect 7929 8415 7987 8421
rect 7929 8381 7941 8415
rect 7975 8412 7987 8415
rect 8478 8412 8484 8424
rect 7975 8384 8484 8412
rect 7975 8381 7987 8384
rect 7929 8375 7987 8381
rect 8478 8372 8484 8384
rect 8536 8372 8542 8424
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 9306 8412 9312 8424
rect 8812 8384 9312 8412
rect 8812 8372 8818 8384
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 9398 8372 9404 8424
rect 9456 8412 9462 8424
rect 9456 8384 9501 8412
rect 9456 8372 9462 8384
rect 9582 8372 9588 8424
rect 9640 8372 9646 8424
rect 9766 8372 9772 8424
rect 9824 8421 9830 8424
rect 11164 8421 11192 8452
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 9824 8412 9832 8421
rect 11149 8415 11207 8421
rect 9824 8384 9869 8412
rect 9824 8375 9832 8384
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 9824 8372 9830 8375
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 11440 8412 11468 8520
rect 11793 8551 11851 8557
rect 11793 8517 11805 8551
rect 11839 8548 11851 8551
rect 11839 8520 12434 8548
rect 11839 8517 11851 8520
rect 11793 8511 11851 8517
rect 11882 8440 11888 8492
rect 11940 8440 11946 8492
rect 12406 8480 12434 8520
rect 12526 8508 12532 8560
rect 12584 8548 12590 8560
rect 12584 8520 12940 8548
rect 12584 8508 12590 8520
rect 12406 8452 12848 8480
rect 11614 8415 11672 8421
rect 11614 8412 11626 8415
rect 11296 8384 11341 8412
rect 11440 8384 11626 8412
rect 11296 8372 11302 8384
rect 11614 8381 11626 8384
rect 11660 8381 11672 8415
rect 11614 8375 11672 8381
rect 12158 8372 12164 8424
rect 12216 8372 12222 8424
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8381 12311 8415
rect 12253 8375 12311 8381
rect 4249 8347 4307 8353
rect 4249 8344 4261 8347
rect 3620 8316 4261 8344
rect 4249 8313 4261 8316
rect 4295 8344 4307 8347
rect 4522 8344 4528 8356
rect 4295 8316 4528 8344
rect 4295 8313 4307 8316
rect 4249 8307 4307 8313
rect 4522 8304 4528 8316
rect 4580 8304 4586 8356
rect 5905 8347 5963 8353
rect 5905 8313 5917 8347
rect 5951 8344 5963 8347
rect 7006 8344 7012 8356
rect 5951 8316 7012 8344
rect 5951 8313 5963 8316
rect 5905 8307 5963 8313
rect 7006 8304 7012 8316
rect 7064 8304 7070 8356
rect 8113 8347 8171 8353
rect 8113 8313 8125 8347
rect 8159 8344 8171 8347
rect 8202 8344 8208 8356
rect 8159 8316 8208 8344
rect 8159 8313 8171 8316
rect 8113 8307 8171 8313
rect 8202 8304 8208 8316
rect 8260 8344 8266 8356
rect 8389 8347 8447 8353
rect 8389 8344 8401 8347
rect 8260 8316 8401 8344
rect 8260 8304 8266 8316
rect 8389 8313 8401 8316
rect 8435 8313 8447 8347
rect 8389 8307 8447 8313
rect 8570 8304 8576 8356
rect 8628 8344 8634 8356
rect 9677 8347 9735 8353
rect 8628 8316 9536 8344
rect 8628 8304 8634 8316
rect 3418 8236 3424 8288
rect 3476 8236 3482 8288
rect 3602 8236 3608 8288
rect 3660 8276 3666 8288
rect 4065 8279 4123 8285
rect 4065 8276 4077 8279
rect 3660 8248 4077 8276
rect 3660 8236 3666 8248
rect 4065 8245 4077 8248
rect 4111 8245 4123 8279
rect 4065 8239 4123 8245
rect 4338 8236 4344 8288
rect 4396 8236 4402 8288
rect 4430 8236 4436 8288
rect 4488 8236 4494 8288
rect 7742 8236 7748 8288
rect 7800 8236 7806 8288
rect 8757 8279 8815 8285
rect 8757 8245 8769 8279
rect 8803 8276 8815 8279
rect 8846 8276 8852 8288
rect 8803 8248 8852 8276
rect 8803 8245 8815 8248
rect 8757 8239 8815 8245
rect 8846 8236 8852 8248
rect 8904 8236 8910 8288
rect 9508 8276 9536 8316
rect 9677 8313 9689 8347
rect 9723 8313 9735 8347
rect 9677 8307 9735 8313
rect 9692 8276 9720 8307
rect 10962 8304 10968 8356
rect 11020 8344 11026 8356
rect 11425 8347 11483 8353
rect 11425 8344 11437 8347
rect 11020 8316 11437 8344
rect 11020 8304 11026 8316
rect 11425 8313 11437 8316
rect 11471 8313 11483 8347
rect 11425 8307 11483 8313
rect 11517 8347 11575 8353
rect 11517 8313 11529 8347
rect 11563 8344 11575 8347
rect 12066 8344 12072 8356
rect 11563 8316 12072 8344
rect 11563 8313 11575 8316
rect 11517 8307 11575 8313
rect 12066 8304 12072 8316
rect 12124 8304 12130 8356
rect 12268 8344 12296 8375
rect 12342 8372 12348 8424
rect 12400 8372 12406 8424
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 12820 8421 12848 8452
rect 12912 8421 12940 8520
rect 12621 8415 12679 8421
rect 12621 8412 12633 8415
rect 12584 8384 12633 8412
rect 12584 8372 12590 8384
rect 12621 8381 12633 8384
rect 12667 8381 12679 8415
rect 12621 8375 12679 8381
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 12434 8344 12440 8356
rect 12268 8316 12440 8344
rect 9508 8248 9720 8276
rect 9953 8279 10011 8285
rect 9953 8245 9965 8279
rect 9999 8276 10011 8279
rect 10318 8276 10324 8288
rect 9999 8248 10324 8276
rect 9999 8245 10011 8248
rect 9953 8239 10011 8245
rect 10318 8236 10324 8248
rect 10376 8236 10382 8288
rect 10410 8236 10416 8288
rect 10468 8276 10474 8288
rect 12268 8276 12296 8316
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 12636 8344 12664 8375
rect 12986 8372 12992 8424
rect 13044 8412 13050 8424
rect 14274 8412 14280 8424
rect 13044 8384 14280 8412
rect 13044 8372 13050 8384
rect 14274 8372 14280 8384
rect 14332 8372 14338 8424
rect 13078 8344 13084 8356
rect 12636 8316 13084 8344
rect 13078 8304 13084 8316
rect 13136 8304 13142 8356
rect 14936 8344 14964 8579
rect 16114 8576 16120 8628
rect 16172 8616 16178 8628
rect 16393 8619 16451 8625
rect 16393 8616 16405 8619
rect 16172 8588 16405 8616
rect 16172 8576 16178 8588
rect 16393 8585 16405 8588
rect 16439 8585 16451 8619
rect 16393 8579 16451 8585
rect 16758 8576 16764 8628
rect 16816 8616 16822 8628
rect 17129 8619 17187 8625
rect 17129 8616 17141 8619
rect 16816 8588 17141 8616
rect 16816 8576 16822 8588
rect 17129 8585 17141 8588
rect 17175 8585 17187 8619
rect 17129 8579 17187 8585
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 20625 8619 20683 8625
rect 20625 8616 20637 8619
rect 19484 8588 20637 8616
rect 19484 8576 19490 8588
rect 20625 8585 20637 8588
rect 20671 8585 20683 8619
rect 20625 8579 20683 8585
rect 17770 8508 17776 8560
rect 17828 8508 17834 8560
rect 20640 8548 20668 8579
rect 22186 8576 22192 8628
rect 22244 8576 22250 8628
rect 22278 8576 22284 8628
rect 22336 8616 22342 8628
rect 22741 8619 22799 8625
rect 22741 8616 22753 8619
rect 22336 8588 22753 8616
rect 22336 8576 22342 8588
rect 22741 8585 22753 8588
rect 22787 8585 22799 8619
rect 22741 8579 22799 8585
rect 22925 8619 22983 8625
rect 22925 8585 22937 8619
rect 22971 8616 22983 8619
rect 23750 8616 23756 8628
rect 22971 8588 23756 8616
rect 22971 8585 22983 8588
rect 22925 8579 22983 8585
rect 23750 8576 23756 8588
rect 23808 8576 23814 8628
rect 24121 8619 24179 8625
rect 24121 8585 24133 8619
rect 24167 8616 24179 8619
rect 24302 8616 24308 8628
rect 24167 8588 24308 8616
rect 24167 8585 24179 8588
rect 24121 8579 24179 8585
rect 24302 8576 24308 8588
rect 24360 8576 24366 8628
rect 25406 8616 25412 8628
rect 25148 8588 25412 8616
rect 22373 8551 22431 8557
rect 22373 8548 22385 8551
rect 20640 8520 21220 8548
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 19245 8483 19303 8489
rect 19245 8480 19257 8483
rect 16356 8452 19257 8480
rect 16356 8440 16362 8452
rect 19245 8449 19257 8452
rect 19291 8449 19303 8483
rect 19245 8443 19303 8449
rect 20898 8440 20904 8492
rect 20956 8440 20962 8492
rect 21192 8489 21220 8520
rect 22066 8520 22385 8548
rect 21177 8483 21235 8489
rect 21177 8449 21189 8483
rect 21223 8480 21235 8483
rect 21358 8480 21364 8492
rect 21223 8452 21364 8480
rect 21223 8449 21235 8452
rect 21177 8443 21235 8449
rect 21358 8440 21364 8452
rect 21416 8440 21422 8492
rect 22066 8480 22094 8520
rect 22373 8517 22385 8520
rect 22419 8548 22431 8551
rect 23106 8548 23112 8560
rect 22419 8520 23112 8548
rect 22419 8517 22431 8520
rect 22373 8511 22431 8517
rect 23106 8508 23112 8520
rect 23164 8508 23170 8560
rect 23566 8508 23572 8560
rect 23624 8548 23630 8560
rect 24029 8551 24087 8557
rect 24029 8548 24041 8551
rect 23624 8520 24041 8548
rect 23624 8508 23630 8520
rect 24029 8517 24041 8520
rect 24075 8517 24087 8551
rect 24029 8511 24087 8517
rect 21836 8452 22094 8480
rect 16022 8372 16028 8424
rect 16080 8421 16086 8424
rect 16080 8412 16092 8421
rect 16945 8415 17003 8421
rect 16080 8384 16125 8412
rect 16080 8375 16092 8384
rect 16945 8381 16957 8415
rect 16991 8381 17003 8415
rect 16945 8375 17003 8381
rect 16080 8372 16086 8375
rect 16960 8344 16988 8375
rect 17034 8372 17040 8424
rect 17092 8412 17098 8424
rect 17129 8415 17187 8421
rect 17129 8412 17141 8415
rect 17092 8384 17141 8412
rect 17092 8372 17098 8384
rect 17129 8381 17141 8384
rect 17175 8381 17187 8415
rect 17129 8375 17187 8381
rect 17402 8372 17408 8424
rect 17460 8372 17466 8424
rect 17586 8372 17592 8424
rect 17644 8412 17650 8424
rect 19334 8412 19340 8424
rect 17644 8384 19340 8412
rect 17644 8372 17650 8384
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 19518 8421 19524 8424
rect 19512 8412 19524 8421
rect 19479 8384 19524 8412
rect 19512 8375 19524 8384
rect 19518 8372 19524 8375
rect 19576 8372 19582 8424
rect 20990 8372 20996 8424
rect 21048 8372 21054 8424
rect 21085 8415 21143 8421
rect 21085 8381 21097 8415
rect 21131 8412 21143 8415
rect 21131 8384 21404 8412
rect 21131 8381 21143 8384
rect 21085 8375 21143 8381
rect 14936 8316 16988 8344
rect 17313 8347 17371 8353
rect 17313 8313 17325 8347
rect 17359 8344 17371 8347
rect 17954 8344 17960 8356
rect 17359 8316 17960 8344
rect 17359 8313 17371 8316
rect 17313 8307 17371 8313
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 18046 8304 18052 8356
rect 18104 8344 18110 8356
rect 21174 8344 21180 8356
rect 18104 8316 21180 8344
rect 18104 8304 18110 8316
rect 21174 8304 21180 8316
rect 21232 8304 21238 8356
rect 21376 8344 21404 8384
rect 21450 8372 21456 8424
rect 21508 8412 21514 8424
rect 21545 8415 21603 8421
rect 21545 8412 21557 8415
rect 21508 8384 21557 8412
rect 21508 8372 21514 8384
rect 21545 8381 21557 8384
rect 21591 8381 21603 8415
rect 21545 8375 21603 8381
rect 21634 8372 21640 8424
rect 21692 8412 21698 8424
rect 21836 8421 21864 8452
rect 23842 8440 23848 8492
rect 23900 8480 23906 8492
rect 24213 8483 24271 8489
rect 24213 8480 24225 8483
rect 23900 8452 24225 8480
rect 23900 8440 23906 8452
rect 24213 8449 24225 8452
rect 24259 8480 24271 8483
rect 24394 8480 24400 8492
rect 24259 8452 24400 8480
rect 24259 8449 24271 8452
rect 24213 8443 24271 8449
rect 24394 8440 24400 8452
rect 24452 8440 24458 8492
rect 24946 8440 24952 8492
rect 25004 8440 25010 8492
rect 25148 8489 25176 8588
rect 25406 8576 25412 8588
rect 25464 8576 25470 8628
rect 25133 8483 25191 8489
rect 25133 8449 25145 8483
rect 25179 8449 25191 8483
rect 25133 8443 25191 8449
rect 21729 8415 21787 8421
rect 21729 8412 21741 8415
rect 21692 8384 21741 8412
rect 21692 8372 21698 8384
rect 21729 8381 21741 8384
rect 21775 8381 21787 8415
rect 21729 8375 21787 8381
rect 21821 8415 21879 8421
rect 21821 8381 21833 8415
rect 21867 8381 21879 8415
rect 21821 8375 21879 8381
rect 21910 8372 21916 8424
rect 21968 8372 21974 8424
rect 23937 8415 23995 8421
rect 23937 8381 23949 8415
rect 23983 8381 23995 8415
rect 23937 8375 23995 8381
rect 21376 8316 21864 8344
rect 21836 8288 21864 8316
rect 22738 8304 22744 8356
rect 22796 8304 22802 8356
rect 22830 8304 22836 8356
rect 22888 8344 22894 8356
rect 23290 8344 23296 8356
rect 22888 8316 23296 8344
rect 22888 8304 22894 8316
rect 23290 8304 23296 8316
rect 23348 8344 23354 8356
rect 23952 8344 23980 8375
rect 24118 8372 24124 8424
rect 24176 8412 24182 8424
rect 24305 8415 24363 8421
rect 24305 8412 24317 8415
rect 24176 8384 24317 8412
rect 24176 8372 24182 8384
rect 24305 8381 24317 8384
rect 24351 8381 24363 8415
rect 24305 8375 24363 8381
rect 24964 8384 26556 8412
rect 24964 8344 24992 8384
rect 23348 8316 24992 8344
rect 25400 8347 25458 8353
rect 23348 8304 23354 8316
rect 25400 8313 25412 8347
rect 25446 8344 25458 8347
rect 25498 8344 25504 8356
rect 25446 8316 25504 8344
rect 25446 8313 25458 8316
rect 25400 8307 25458 8313
rect 25498 8304 25504 8316
rect 25556 8304 25562 8356
rect 26528 8288 26556 8384
rect 10468 8248 12296 8276
rect 10468 8236 10474 8248
rect 13262 8236 13268 8288
rect 13320 8236 13326 8288
rect 20717 8279 20775 8285
rect 20717 8245 20729 8279
rect 20763 8276 20775 8279
rect 20898 8276 20904 8288
rect 20763 8248 20904 8276
rect 20763 8245 20775 8248
rect 20717 8239 20775 8245
rect 20898 8236 20904 8248
rect 20956 8236 20962 8288
rect 21818 8236 21824 8288
rect 21876 8236 21882 8288
rect 23014 8236 23020 8288
rect 23072 8276 23078 8288
rect 25682 8276 25688 8288
rect 23072 8248 25688 8276
rect 23072 8236 23078 8248
rect 25682 8236 25688 8248
rect 25740 8236 25746 8288
rect 26510 8236 26516 8288
rect 26568 8236 26574 8288
rect 552 8186 27576 8208
rect 552 8134 7114 8186
rect 7166 8134 7178 8186
rect 7230 8134 7242 8186
rect 7294 8134 7306 8186
rect 7358 8134 7370 8186
rect 7422 8134 13830 8186
rect 13882 8134 13894 8186
rect 13946 8134 13958 8186
rect 14010 8134 14022 8186
rect 14074 8134 14086 8186
rect 14138 8134 20546 8186
rect 20598 8134 20610 8186
rect 20662 8134 20674 8186
rect 20726 8134 20738 8186
rect 20790 8134 20802 8186
rect 20854 8134 27262 8186
rect 27314 8134 27326 8186
rect 27378 8134 27390 8186
rect 27442 8134 27454 8186
rect 27506 8134 27518 8186
rect 27570 8134 27576 8186
rect 552 8112 27576 8134
rect 2593 8075 2651 8081
rect 2593 8041 2605 8075
rect 2639 8041 2651 8075
rect 2593 8035 2651 8041
rect 2608 8004 2636 8035
rect 4062 8032 4068 8084
rect 4120 8032 4126 8084
rect 6917 8075 6975 8081
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 7558 8072 7564 8084
rect 6963 8044 7564 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 7742 8032 7748 8084
rect 7800 8032 7806 8084
rect 8478 8032 8484 8084
rect 8536 8032 8542 8084
rect 8570 8032 8576 8084
rect 8628 8072 8634 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 8628 8044 9321 8072
rect 8628 8032 8634 8044
rect 9309 8041 9321 8044
rect 9355 8041 9367 8075
rect 12526 8072 12532 8084
rect 9309 8035 9367 8041
rect 12084 8044 12532 8072
rect 2930 8007 2988 8013
rect 2930 8004 2942 8007
rect 2608 7976 2942 8004
rect 2930 7973 2942 7976
rect 2976 7973 2988 8007
rect 7760 8004 7788 8032
rect 2930 7967 2988 7973
rect 6380 7976 7788 8004
rect 8496 8004 8524 8032
rect 9769 8007 9827 8013
rect 9769 8004 9781 8007
rect 8496 7976 9781 8004
rect 2406 7896 2412 7948
rect 2464 7896 2470 7948
rect 2682 7896 2688 7948
rect 2740 7896 2746 7948
rect 6380 7945 6408 7976
rect 9769 7973 9781 7976
rect 9815 7973 9827 8007
rect 9769 7967 9827 7973
rect 10042 7964 10048 8016
rect 10100 8004 10106 8016
rect 12084 8004 12112 8044
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 19889 8075 19947 8081
rect 19889 8041 19901 8075
rect 19935 8072 19947 8075
rect 20898 8072 20904 8084
rect 19935 8044 20904 8072
rect 19935 8041 19947 8044
rect 19889 8035 19947 8041
rect 20898 8032 20904 8044
rect 20956 8032 20962 8084
rect 20990 8032 20996 8084
rect 21048 8072 21054 8084
rect 21637 8075 21695 8081
rect 21637 8072 21649 8075
rect 21048 8044 21649 8072
rect 21048 8032 21054 8044
rect 21637 8041 21649 8044
rect 21683 8041 21695 8075
rect 21637 8035 21695 8041
rect 10100 7976 12112 8004
rect 10100 7964 10106 7976
rect 6181 7939 6239 7945
rect 6181 7905 6193 7939
rect 6227 7905 6239 7939
rect 6181 7899 6239 7905
rect 6365 7939 6423 7945
rect 6365 7905 6377 7939
rect 6411 7905 6423 7939
rect 6365 7899 6423 7905
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7936 6699 7939
rect 6730 7936 6736 7948
rect 6687 7908 6736 7936
rect 6687 7905 6699 7908
rect 6641 7899 6699 7905
rect 6196 7868 6224 7899
rect 6730 7896 6736 7908
rect 6788 7936 6794 7948
rect 7101 7939 7159 7945
rect 7101 7936 7113 7939
rect 6788 7908 7113 7936
rect 6788 7896 6794 7908
rect 7101 7905 7113 7908
rect 7147 7905 7159 7939
rect 7101 7899 7159 7905
rect 7282 7896 7288 7948
rect 7340 7896 7346 7948
rect 7374 7896 7380 7948
rect 7432 7896 7438 7948
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7936 7619 7939
rect 9030 7936 9036 7948
rect 7607 7908 9036 7936
rect 7607 7905 7619 7908
rect 7561 7899 7619 7905
rect 6270 7868 6276 7880
rect 6196 7840 6276 7868
rect 6270 7828 6276 7840
rect 6328 7868 6334 7880
rect 7576 7868 7604 7899
rect 9030 7896 9036 7908
rect 9088 7896 9094 7948
rect 9306 7896 9312 7948
rect 9364 7936 9370 7948
rect 9401 7939 9459 7945
rect 9401 7936 9413 7939
rect 9364 7908 9413 7936
rect 9364 7896 9370 7908
rect 9401 7905 9413 7908
rect 9447 7905 9459 7939
rect 9401 7899 9459 7905
rect 9490 7896 9496 7948
rect 9548 7936 9554 7948
rect 9548 7908 9593 7936
rect 9548 7896 9554 7908
rect 9674 7896 9680 7948
rect 9732 7896 9738 7948
rect 9858 7896 9864 7948
rect 9916 7945 9922 7948
rect 10152 7945 10180 7976
rect 9916 7936 9924 7945
rect 10137 7939 10195 7945
rect 9916 7908 9961 7936
rect 9916 7899 9924 7908
rect 10137 7905 10149 7939
rect 10183 7905 10195 7939
rect 10137 7899 10195 7905
rect 9916 7896 9922 7899
rect 10318 7896 10324 7948
rect 10376 7896 10382 7948
rect 10410 7896 10416 7948
rect 10468 7896 10474 7948
rect 12084 7945 12112 7976
rect 13072 8007 13130 8013
rect 13072 7973 13084 8007
rect 13118 8004 13130 8007
rect 13262 8004 13268 8016
rect 13118 7976 13268 8004
rect 13118 7973 13130 7976
rect 13072 7967 13130 7973
rect 13262 7964 13268 7976
rect 13320 7964 13326 8016
rect 21652 8004 21680 8035
rect 21726 8032 21732 8084
rect 21784 8032 21790 8084
rect 21818 8032 21824 8084
rect 21876 8072 21882 8084
rect 24673 8075 24731 8081
rect 24673 8072 24685 8075
rect 21876 8044 24685 8072
rect 21876 8032 21882 8044
rect 22370 8004 22376 8016
rect 21652 7976 22376 8004
rect 10505 7939 10563 7945
rect 10505 7905 10517 7939
rect 10551 7936 10563 7939
rect 11333 7939 11391 7945
rect 11333 7936 11345 7939
rect 10551 7908 11345 7936
rect 10551 7905 10563 7908
rect 10505 7899 10563 7905
rect 11333 7905 11345 7908
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 12069 7939 12127 7945
rect 12069 7905 12081 7939
rect 12115 7905 12127 7939
rect 12069 7899 12127 7905
rect 12253 7939 12311 7945
rect 12253 7905 12265 7939
rect 12299 7905 12311 7939
rect 12253 7899 12311 7905
rect 6328 7840 7604 7868
rect 6328 7828 6334 7840
rect 7926 7828 7932 7880
rect 7984 7828 7990 7880
rect 8754 7828 8760 7880
rect 8812 7828 8818 7880
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 11296 7840 11989 7868
rect 11296 7828 11302 7840
rect 11977 7837 11989 7840
rect 12023 7868 12035 7871
rect 12158 7868 12164 7880
rect 12023 7840 12164 7868
rect 12023 7837 12035 7840
rect 11977 7831 12035 7837
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 5902 7760 5908 7812
rect 5960 7800 5966 7812
rect 6457 7803 6515 7809
rect 6457 7800 6469 7803
rect 5960 7772 6469 7800
rect 5960 7760 5966 7772
rect 6457 7769 6469 7772
rect 6503 7769 6515 7803
rect 6457 7763 6515 7769
rect 6549 7803 6607 7809
rect 6549 7769 6561 7803
rect 6595 7800 6607 7803
rect 7193 7803 7251 7809
rect 6595 7772 7144 7800
rect 6595 7769 6607 7772
rect 6549 7763 6607 7769
rect 6822 7692 6828 7744
rect 6880 7692 6886 7744
rect 7116 7732 7144 7772
rect 7193 7769 7205 7803
rect 7239 7800 7251 7803
rect 7834 7800 7840 7812
rect 7239 7772 7840 7800
rect 7239 7769 7251 7772
rect 7193 7763 7251 7769
rect 7834 7760 7840 7772
rect 7892 7760 7898 7812
rect 8570 7760 8576 7812
rect 8628 7800 8634 7812
rect 9858 7800 9864 7812
rect 8628 7772 9864 7800
rect 8628 7760 8634 7772
rect 9858 7760 9864 7772
rect 9916 7760 9922 7812
rect 10045 7803 10103 7809
rect 10045 7769 10057 7803
rect 10091 7800 10103 7803
rect 12268 7800 12296 7899
rect 12342 7896 12348 7948
rect 12400 7936 12406 7948
rect 12483 7939 12541 7945
rect 12400 7908 12445 7936
rect 12400 7896 12406 7908
rect 12483 7905 12495 7939
rect 12529 7936 12541 7939
rect 12710 7936 12716 7948
rect 12529 7908 12716 7936
rect 12529 7905 12541 7908
rect 12483 7899 12541 7905
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 20717 7939 20775 7945
rect 20717 7905 20729 7939
rect 20763 7936 20775 7939
rect 21174 7936 21180 7948
rect 20763 7908 21180 7936
rect 20763 7905 20775 7908
rect 20717 7899 20775 7905
rect 21174 7896 21180 7908
rect 21232 7896 21238 7948
rect 21358 7896 21364 7948
rect 21416 7896 21422 7948
rect 21545 7939 21603 7945
rect 21545 7905 21557 7939
rect 21591 7936 21603 7939
rect 21818 7936 21824 7948
rect 21591 7908 21824 7936
rect 21591 7905 21603 7908
rect 21545 7899 21603 7905
rect 21818 7896 21824 7908
rect 21876 7896 21882 7948
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 10091 7772 12296 7800
rect 10091 7769 10103 7772
rect 10045 7763 10103 7769
rect 12342 7760 12348 7812
rect 12400 7800 12406 7812
rect 12820 7800 12848 7831
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 20993 7871 21051 7877
rect 20993 7868 21005 7871
rect 13872 7840 21005 7868
rect 13872 7828 13878 7840
rect 20993 7837 21005 7840
rect 21039 7868 21051 7871
rect 21450 7868 21456 7880
rect 21039 7840 21456 7868
rect 21039 7837 21051 7840
rect 20993 7831 21051 7837
rect 21450 7828 21456 7840
rect 21508 7828 21514 7880
rect 22296 7868 22324 7976
rect 22370 7964 22376 7976
rect 22428 7964 22434 8016
rect 22489 7877 22517 8044
rect 24673 8041 24685 8044
rect 24719 8072 24731 8075
rect 24946 8072 24952 8084
rect 24719 8044 24952 8072
rect 24719 8041 24731 8044
rect 24673 8035 24731 8041
rect 22646 7964 22652 8016
rect 22704 8004 22710 8016
rect 23750 8004 23756 8016
rect 22704 7976 23756 8004
rect 22704 7964 22710 7976
rect 23750 7964 23756 7976
rect 23808 8004 23814 8016
rect 23808 7976 24440 8004
rect 23808 7964 23814 7976
rect 22557 7939 22615 7945
rect 22557 7905 22569 7939
rect 22603 7936 22615 7939
rect 22830 7936 22836 7948
rect 22603 7908 22836 7936
rect 22603 7905 22615 7908
rect 22557 7899 22615 7905
rect 22830 7896 22836 7908
rect 22888 7896 22894 7948
rect 23014 7896 23020 7948
rect 23072 7896 23078 7948
rect 23198 7896 23204 7948
rect 23256 7896 23262 7948
rect 23290 7896 23296 7948
rect 23348 7896 23354 7948
rect 23474 7896 23480 7948
rect 23532 7896 23538 7948
rect 24044 7945 24072 7976
rect 24029 7939 24087 7945
rect 24029 7905 24041 7939
rect 24075 7905 24087 7939
rect 24029 7899 24087 7905
rect 24118 7896 24124 7948
rect 24176 7896 24182 7948
rect 24412 7945 24440 7976
rect 24397 7939 24455 7945
rect 24397 7905 24409 7939
rect 24443 7905 24455 7939
rect 24397 7899 24455 7905
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 22296 7840 22385 7868
rect 22373 7837 22385 7840
rect 22419 7837 22431 7871
rect 22373 7831 22431 7837
rect 22465 7871 22523 7877
rect 22465 7837 22477 7871
rect 22511 7837 22523 7871
rect 22465 7831 22523 7837
rect 22649 7871 22707 7877
rect 22649 7837 22661 7871
rect 22695 7868 22707 7871
rect 23216 7868 23244 7896
rect 22695 7840 23244 7868
rect 22695 7837 22707 7840
rect 22649 7831 22707 7837
rect 23566 7828 23572 7880
rect 23624 7868 23630 7880
rect 23842 7868 23848 7880
rect 23624 7840 23848 7868
rect 23624 7828 23630 7840
rect 23842 7828 23848 7840
rect 23900 7828 23906 7880
rect 24213 7871 24271 7877
rect 24213 7837 24225 7871
rect 24259 7868 24271 7871
rect 24688 7868 24716 8035
rect 24946 8032 24952 8044
rect 25004 8032 25010 8084
rect 26418 8032 26424 8084
rect 26476 8032 26482 8084
rect 25406 7964 25412 8016
rect 25464 8004 25470 8016
rect 25464 7976 26096 8004
rect 25464 7964 25470 7976
rect 25498 7896 25504 7948
rect 25556 7936 25562 7948
rect 26068 7945 26096 7976
rect 25786 7939 25844 7945
rect 25786 7936 25798 7939
rect 25556 7908 25798 7936
rect 25556 7896 25562 7908
rect 25786 7905 25798 7908
rect 25832 7905 25844 7939
rect 25786 7899 25844 7905
rect 26053 7939 26111 7945
rect 26053 7905 26065 7939
rect 26099 7905 26111 7939
rect 26053 7899 26111 7905
rect 26510 7896 26516 7948
rect 26568 7936 26574 7948
rect 26973 7939 27031 7945
rect 26973 7936 26985 7939
rect 26568 7908 26985 7936
rect 26568 7896 26574 7908
rect 26973 7905 26985 7908
rect 27019 7905 27031 7939
rect 26973 7899 27031 7905
rect 24259 7840 24716 7868
rect 24259 7837 24271 7840
rect 24213 7831 24271 7837
rect 12400 7772 12848 7800
rect 12400 7760 12406 7772
rect 17402 7760 17408 7812
rect 17460 7800 17466 7812
rect 19521 7803 19579 7809
rect 19521 7800 19533 7803
rect 17460 7772 19533 7800
rect 17460 7760 17466 7772
rect 19521 7769 19533 7772
rect 19567 7800 19579 7803
rect 19567 7772 20024 7800
rect 19567 7769 19579 7772
rect 19521 7763 19579 7769
rect 8938 7732 8944 7744
rect 7116 7704 8944 7732
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 10781 7735 10839 7741
rect 10781 7701 10793 7735
rect 10827 7732 10839 7735
rect 11330 7732 11336 7744
rect 10827 7704 11336 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 11330 7692 11336 7704
rect 11388 7692 11394 7744
rect 12713 7735 12771 7741
rect 12713 7701 12725 7735
rect 12759 7732 12771 7735
rect 13814 7732 13820 7744
rect 12759 7704 13820 7732
rect 12759 7701 12771 7704
rect 12713 7695 12771 7701
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 14185 7735 14243 7741
rect 14185 7701 14197 7735
rect 14231 7732 14243 7735
rect 14274 7732 14280 7744
rect 14231 7704 14280 7732
rect 14231 7701 14243 7704
rect 14185 7695 14243 7701
rect 14274 7692 14280 7704
rect 14332 7732 14338 7744
rect 15378 7732 15384 7744
rect 14332 7704 15384 7732
rect 14332 7692 14338 7704
rect 15378 7692 15384 7704
rect 15436 7692 15442 7744
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 19886 7732 19892 7744
rect 19392 7704 19892 7732
rect 19392 7692 19398 7704
rect 19886 7692 19892 7704
rect 19944 7692 19950 7744
rect 19996 7732 20024 7772
rect 20070 7760 20076 7812
rect 20128 7760 20134 7812
rect 22278 7760 22284 7812
rect 22336 7800 22342 7812
rect 23201 7803 23259 7809
rect 23201 7800 23213 7803
rect 22336 7772 23213 7800
rect 22336 7760 22342 7772
rect 23201 7769 23213 7772
rect 23247 7769 23259 7803
rect 23201 7763 23259 7769
rect 23937 7803 23995 7809
rect 23937 7769 23949 7803
rect 23983 7800 23995 7803
rect 23983 7772 25176 7800
rect 23983 7769 23995 7772
rect 23937 7763 23995 7769
rect 21913 7735 21971 7741
rect 21913 7732 21925 7735
rect 19996 7704 21925 7732
rect 21913 7701 21925 7704
rect 21959 7701 21971 7735
rect 21913 7695 21971 7701
rect 22186 7692 22192 7744
rect 22244 7692 22250 7744
rect 22370 7692 22376 7744
rect 22428 7732 22434 7744
rect 22925 7735 22983 7741
rect 22925 7732 22937 7735
rect 22428 7704 22937 7732
rect 22428 7692 22434 7704
rect 22925 7701 22937 7704
rect 22971 7701 22983 7735
rect 22925 7695 22983 7701
rect 24578 7692 24584 7744
rect 24636 7692 24642 7744
rect 25148 7732 25176 7772
rect 25314 7732 25320 7744
rect 25148 7704 25320 7732
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 552 7642 27416 7664
rect 552 7590 3756 7642
rect 3808 7590 3820 7642
rect 3872 7590 3884 7642
rect 3936 7590 3948 7642
rect 4000 7590 4012 7642
rect 4064 7590 10472 7642
rect 10524 7590 10536 7642
rect 10588 7590 10600 7642
rect 10652 7590 10664 7642
rect 10716 7590 10728 7642
rect 10780 7590 17188 7642
rect 17240 7590 17252 7642
rect 17304 7590 17316 7642
rect 17368 7590 17380 7642
rect 17432 7590 17444 7642
rect 17496 7590 23904 7642
rect 23956 7590 23968 7642
rect 24020 7590 24032 7642
rect 24084 7590 24096 7642
rect 24148 7590 24160 7642
rect 24212 7590 27416 7642
rect 552 7568 27416 7590
rect 2406 7488 2412 7540
rect 2464 7528 2470 7540
rect 3237 7531 3295 7537
rect 3237 7528 3249 7531
rect 2464 7500 3249 7528
rect 2464 7488 2470 7500
rect 3237 7497 3249 7500
rect 3283 7497 3295 7531
rect 3237 7491 3295 7497
rect 3421 7531 3479 7537
rect 3421 7497 3433 7531
rect 3467 7528 3479 7531
rect 3510 7528 3516 7540
rect 3467 7500 3516 7528
rect 3467 7497 3479 7500
rect 3421 7491 3479 7497
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 5902 7488 5908 7540
rect 5960 7488 5966 7540
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 6788 7500 7512 7528
rect 6788 7488 6794 7500
rect 3326 7420 3332 7472
rect 3384 7460 3390 7472
rect 4065 7463 4123 7469
rect 4065 7460 4077 7463
rect 3384 7432 4077 7460
rect 3384 7420 3390 7432
rect 4065 7429 4077 7432
rect 4111 7429 4123 7463
rect 7484 7460 7512 7500
rect 7926 7488 7932 7540
rect 7984 7488 7990 7540
rect 11238 7528 11244 7540
rect 8312 7500 11244 7528
rect 8312 7460 8340 7500
rect 11238 7488 11244 7500
rect 11296 7528 11302 7540
rect 11296 7500 14596 7528
rect 11296 7488 11302 7500
rect 7484 7432 8340 7460
rect 4065 7423 4123 7429
rect 3602 7352 3608 7404
rect 3660 7392 3666 7404
rect 3789 7395 3847 7401
rect 3789 7392 3801 7395
rect 3660 7364 3801 7392
rect 3660 7352 3666 7364
rect 3789 7361 3801 7364
rect 3835 7361 3847 7395
rect 3789 7355 3847 7361
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 3510 7284 3516 7336
rect 3568 7324 3574 7336
rect 3896 7324 3924 7355
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 5500 7364 6009 7392
rect 5500 7352 5506 7364
rect 5997 7361 6009 7364
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 3568 7296 3924 7324
rect 3568 7284 3574 7296
rect 4154 7284 4160 7336
rect 4212 7284 4218 7336
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7293 4307 7327
rect 4249 7287 4307 7293
rect 3418 7216 3424 7268
rect 3476 7216 3482 7268
rect 3881 7259 3939 7265
rect 3881 7225 3893 7259
rect 3927 7256 3939 7259
rect 4264 7256 4292 7287
rect 4430 7284 4436 7336
rect 4488 7284 4494 7336
rect 4522 7284 4528 7336
rect 4580 7284 4586 7336
rect 5350 7284 5356 7336
rect 5408 7324 5414 7336
rect 5537 7327 5595 7333
rect 5537 7324 5549 7327
rect 5408 7296 5549 7324
rect 5408 7284 5414 7296
rect 5537 7293 5549 7296
rect 5583 7293 5595 7327
rect 5537 7287 5595 7293
rect 5718 7284 5724 7336
rect 5776 7324 5782 7336
rect 6178 7324 6184 7336
rect 5776 7296 6184 7324
rect 5776 7284 5782 7296
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 6546 7284 6552 7336
rect 6604 7284 6610 7336
rect 6822 7333 6828 7336
rect 6816 7324 6828 7333
rect 6783 7296 6828 7324
rect 6816 7287 6828 7296
rect 6822 7284 6828 7287
rect 6880 7284 6886 7336
rect 8312 7324 8340 7432
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 8444 7364 8677 7392
rect 8444 7352 8450 7364
rect 8665 7361 8677 7364
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 8312 7296 8585 7324
rect 8573 7293 8585 7296
rect 8619 7293 8631 7327
rect 8573 7287 8631 7293
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7293 8815 7327
rect 8757 7287 8815 7293
rect 3927 7228 4292 7256
rect 6365 7259 6423 7265
rect 3927 7225 3939 7228
rect 3881 7219 3939 7225
rect 6365 7225 6377 7259
rect 6411 7256 6423 7259
rect 8772 7256 8800 7287
rect 8846 7284 8852 7336
rect 8904 7284 8910 7336
rect 9030 7284 9036 7336
rect 9088 7284 9094 7336
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7324 9643 7327
rect 10962 7324 10968 7336
rect 9631 7296 10968 7324
rect 9631 7293 9643 7296
rect 9585 7287 9643 7293
rect 10962 7284 10968 7296
rect 11020 7324 11026 7336
rect 11057 7327 11115 7333
rect 11057 7324 11069 7327
rect 11020 7296 11069 7324
rect 11020 7284 11026 7296
rect 11057 7293 11069 7296
rect 11103 7324 11115 7327
rect 12342 7324 12348 7336
rect 11103 7296 12348 7324
rect 11103 7293 11115 7296
rect 11057 7287 11115 7293
rect 12342 7284 12348 7296
rect 12400 7324 12406 7336
rect 13814 7333 13820 7336
rect 13541 7327 13599 7333
rect 13541 7324 13553 7327
rect 12400 7296 13553 7324
rect 12400 7284 12406 7296
rect 13541 7293 13553 7296
rect 13587 7293 13599 7327
rect 13808 7324 13820 7333
rect 13775 7296 13820 7324
rect 13541 7287 13599 7293
rect 13808 7287 13820 7296
rect 13814 7284 13820 7287
rect 13872 7284 13878 7336
rect 14568 7324 14596 7500
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 15381 7531 15439 7537
rect 15381 7528 15393 7531
rect 15252 7500 15393 7528
rect 15252 7488 15258 7500
rect 15381 7497 15393 7500
rect 15427 7497 15439 7531
rect 15381 7491 15439 7497
rect 15930 7488 15936 7540
rect 15988 7488 15994 7540
rect 18509 7531 18567 7537
rect 18509 7497 18521 7531
rect 18555 7528 18567 7531
rect 18782 7528 18788 7540
rect 18555 7500 18788 7528
rect 18555 7497 18567 7500
rect 18509 7491 18567 7497
rect 18782 7488 18788 7500
rect 18840 7528 18846 7540
rect 18840 7500 19104 7528
rect 18840 7488 18846 7500
rect 19076 7469 19104 7500
rect 19886 7488 19892 7540
rect 19944 7528 19950 7540
rect 23014 7528 23020 7540
rect 19944 7500 23020 7528
rect 19944 7488 19950 7500
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 23474 7488 23480 7540
rect 23532 7528 23538 7540
rect 25133 7531 25191 7537
rect 25133 7528 25145 7531
rect 23532 7500 25145 7528
rect 23532 7488 23538 7500
rect 25133 7497 25145 7500
rect 25179 7497 25191 7531
rect 25133 7491 25191 7497
rect 25317 7531 25375 7537
rect 25317 7497 25329 7531
rect 25363 7528 25375 7531
rect 25498 7528 25504 7540
rect 25363 7500 25504 7528
rect 25363 7497 25375 7500
rect 25317 7491 25375 7497
rect 19061 7463 19119 7469
rect 19061 7429 19073 7463
rect 19107 7429 19119 7463
rect 19061 7423 19119 7429
rect 16040 7364 16252 7392
rect 16040 7336 16068 7364
rect 15565 7327 15623 7333
rect 15565 7324 15577 7327
rect 14568 7296 15577 7324
rect 15565 7293 15577 7296
rect 15611 7293 15623 7327
rect 15565 7287 15623 7293
rect 15841 7327 15899 7333
rect 15841 7293 15853 7327
rect 15887 7324 15899 7327
rect 16022 7324 16028 7336
rect 15887 7296 16028 7324
rect 15887 7293 15899 7296
rect 15841 7287 15899 7293
rect 6411 7228 8800 7256
rect 9852 7259 9910 7265
rect 6411 7225 6423 7228
rect 6365 7219 6423 7225
rect 9852 7225 9864 7259
rect 9898 7256 9910 7259
rect 10870 7256 10876 7268
rect 9898 7228 10876 7256
rect 9898 7225 9910 7228
rect 9852 7219 9910 7225
rect 10870 7216 10876 7228
rect 10928 7216 10934 7268
rect 11330 7265 11336 7268
rect 11324 7256 11336 7265
rect 11291 7228 11336 7256
rect 11324 7219 11336 7228
rect 11330 7216 11336 7219
rect 11388 7216 11394 7268
rect 15580 7256 15608 7287
rect 16022 7284 16028 7296
rect 16080 7284 16086 7336
rect 16117 7327 16175 7333
rect 16117 7293 16129 7327
rect 16163 7293 16175 7327
rect 16224 7324 16252 7364
rect 16298 7352 16304 7404
rect 16356 7392 16362 7404
rect 17129 7395 17187 7401
rect 17129 7392 17141 7395
rect 16356 7364 17141 7392
rect 16356 7352 16362 7364
rect 17129 7361 17141 7364
rect 17175 7361 17187 7395
rect 20254 7392 20260 7404
rect 17129 7355 17187 7361
rect 18616 7364 20260 7392
rect 16393 7327 16451 7333
rect 16393 7324 16405 7327
rect 16224 7296 16405 7324
rect 16117 7287 16175 7293
rect 16393 7293 16405 7296
rect 16439 7293 16451 7327
rect 18616 7324 18644 7364
rect 20254 7352 20260 7364
rect 20312 7352 20318 7404
rect 25148 7392 25176 7491
rect 25498 7488 25504 7500
rect 25556 7488 25562 7540
rect 25774 7460 25780 7472
rect 25516 7432 25780 7460
rect 25516 7392 25544 7432
rect 25774 7420 25780 7432
rect 25832 7420 25838 7472
rect 25148 7364 25544 7392
rect 16393 7287 16451 7293
rect 17328 7296 18644 7324
rect 16132 7256 16160 7287
rect 17328 7256 17356 7296
rect 18690 7284 18696 7336
rect 18748 7324 18754 7336
rect 18748 7296 18828 7324
rect 18748 7284 18754 7296
rect 15580 7228 16160 7256
rect 16224 7228 17356 7256
rect 17396 7259 17454 7265
rect 4338 7148 4344 7200
rect 4396 7148 4402 7200
rect 4709 7191 4767 7197
rect 4709 7157 4721 7191
rect 4755 7188 4767 7191
rect 4798 7188 4804 7200
rect 4755 7160 4804 7188
rect 4755 7157 4767 7160
rect 4709 7151 4767 7157
rect 4798 7148 4804 7160
rect 4856 7188 4862 7200
rect 5258 7188 5264 7200
rect 4856 7160 5264 7188
rect 4856 7148 4862 7160
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8389 7191 8447 7197
rect 8389 7188 8401 7191
rect 8352 7160 8401 7188
rect 8352 7148 8358 7160
rect 8389 7157 8401 7160
rect 8435 7157 8447 7191
rect 8389 7151 8447 7157
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 11422 7188 11428 7200
rect 11011 7160 11428 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 12158 7148 12164 7200
rect 12216 7188 12222 7200
rect 12437 7191 12495 7197
rect 12437 7188 12449 7191
rect 12216 7160 12449 7188
rect 12216 7148 12222 7160
rect 12437 7157 12449 7160
rect 12483 7157 12495 7191
rect 12437 7151 12495 7157
rect 12802 7148 12808 7200
rect 12860 7188 12866 7200
rect 14921 7191 14979 7197
rect 14921 7188 14933 7191
rect 12860 7160 14933 7188
rect 12860 7148 12866 7160
rect 14921 7157 14933 7160
rect 14967 7157 14979 7191
rect 14921 7151 14979 7157
rect 15749 7191 15807 7197
rect 15749 7157 15761 7191
rect 15795 7188 15807 7191
rect 16224 7188 16252 7228
rect 17396 7225 17408 7259
rect 17442 7256 17454 7259
rect 18800 7256 18828 7296
rect 18874 7284 18880 7336
rect 18932 7284 18938 7336
rect 19334 7284 19340 7336
rect 19392 7324 19398 7336
rect 19429 7327 19487 7333
rect 19429 7324 19441 7327
rect 19392 7296 19441 7324
rect 19392 7284 19398 7296
rect 19429 7293 19441 7296
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 21450 7284 21456 7336
rect 21508 7284 21514 7336
rect 21726 7284 21732 7336
rect 21784 7284 21790 7336
rect 24578 7284 24584 7336
rect 24636 7324 24642 7336
rect 25041 7327 25099 7333
rect 25041 7324 25053 7327
rect 24636 7296 25053 7324
rect 24636 7284 24642 7296
rect 25041 7293 25053 7296
rect 25087 7293 25099 7327
rect 25041 7287 25099 7293
rect 25314 7284 25320 7336
rect 25372 7284 25378 7336
rect 25516 7333 25544 7364
rect 25501 7327 25559 7333
rect 25501 7293 25513 7327
rect 25547 7293 25559 7327
rect 25501 7287 25559 7293
rect 25593 7327 25651 7333
rect 25593 7293 25605 7327
rect 25639 7293 25651 7327
rect 25593 7287 25651 7293
rect 19245 7259 19303 7265
rect 19245 7256 19257 7259
rect 17442 7228 18736 7256
rect 18800 7228 19257 7256
rect 17442 7225 17454 7228
rect 17396 7219 17454 7225
rect 15795 7160 16252 7188
rect 16301 7191 16359 7197
rect 15795 7157 15807 7160
rect 15749 7151 15807 7157
rect 16301 7157 16313 7191
rect 16347 7188 16359 7191
rect 18598 7188 18604 7200
rect 16347 7160 18604 7188
rect 16347 7157 16359 7160
rect 16301 7151 16359 7157
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 18708 7197 18736 7228
rect 19245 7225 19257 7228
rect 19291 7225 19303 7259
rect 19245 7219 19303 7225
rect 23382 7216 23388 7268
rect 23440 7216 23446 7268
rect 23750 7216 23756 7268
rect 23808 7256 23814 7268
rect 25608 7256 25636 7287
rect 25774 7284 25780 7336
rect 25832 7284 25838 7336
rect 23808 7228 25636 7256
rect 23808 7216 23814 7228
rect 18693 7191 18751 7197
rect 18693 7157 18705 7191
rect 18739 7157 18751 7191
rect 18693 7151 18751 7157
rect 19337 7191 19395 7197
rect 19337 7157 19349 7191
rect 19383 7188 19395 7191
rect 19518 7188 19524 7200
rect 19383 7160 19524 7188
rect 19383 7157 19395 7160
rect 19337 7151 19395 7157
rect 19518 7148 19524 7160
rect 19576 7148 19582 7200
rect 19613 7191 19671 7197
rect 19613 7157 19625 7191
rect 19659 7188 19671 7191
rect 19702 7188 19708 7200
rect 19659 7160 19708 7188
rect 19659 7157 19671 7160
rect 19613 7151 19671 7157
rect 19702 7148 19708 7160
rect 19760 7148 19766 7200
rect 21637 7191 21695 7197
rect 21637 7157 21649 7191
rect 21683 7188 21695 7191
rect 22094 7188 22100 7200
rect 21683 7160 22100 7188
rect 21683 7157 21695 7160
rect 21637 7151 21695 7157
rect 22094 7148 22100 7160
rect 22152 7148 22158 7200
rect 25682 7148 25688 7200
rect 25740 7148 25746 7200
rect 552 7098 27576 7120
rect 552 7046 7114 7098
rect 7166 7046 7178 7098
rect 7230 7046 7242 7098
rect 7294 7046 7306 7098
rect 7358 7046 7370 7098
rect 7422 7046 13830 7098
rect 13882 7046 13894 7098
rect 13946 7046 13958 7098
rect 14010 7046 14022 7098
rect 14074 7046 14086 7098
rect 14138 7046 20546 7098
rect 20598 7046 20610 7098
rect 20662 7046 20674 7098
rect 20726 7046 20738 7098
rect 20790 7046 20802 7098
rect 20854 7046 27262 7098
rect 27314 7046 27326 7098
rect 27378 7046 27390 7098
rect 27442 7046 27454 7098
rect 27506 7046 27518 7098
rect 27570 7046 27576 7098
rect 552 7024 27576 7046
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 4081 6987 4139 6993
rect 4081 6984 4093 6987
rect 3660 6956 4093 6984
rect 3660 6944 3666 6956
rect 4081 6953 4093 6956
rect 4127 6984 4139 6987
rect 4127 6956 4200 6984
rect 4127 6953 4139 6956
rect 4081 6947 4139 6953
rect 3881 6919 3939 6925
rect 3881 6885 3893 6919
rect 3927 6916 3939 6919
rect 4172 6916 4200 6956
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 4341 6987 4399 6993
rect 4341 6984 4353 6987
rect 4304 6956 4353 6984
rect 4304 6944 4310 6956
rect 4341 6953 4353 6956
rect 4387 6953 4399 6987
rect 5261 6987 5319 6993
rect 5261 6984 5273 6987
rect 4341 6947 4399 6953
rect 4448 6956 5273 6984
rect 4448 6916 4476 6956
rect 5261 6953 5273 6956
rect 5307 6953 5319 6987
rect 5261 6947 5319 6953
rect 5350 6944 5356 6996
rect 5408 6944 5414 6996
rect 5442 6944 5448 6996
rect 5500 6944 5506 6996
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 8849 6987 8907 6993
rect 8849 6984 8861 6987
rect 8812 6956 8861 6984
rect 8812 6944 8818 6956
rect 8849 6953 8861 6956
rect 8895 6953 8907 6987
rect 13909 6987 13967 6993
rect 13909 6984 13921 6987
rect 8849 6947 8907 6953
rect 13464 6956 13921 6984
rect 5460 6916 5488 6944
rect 3927 6888 4016 6916
rect 4172 6888 4476 6916
rect 5000 6888 5488 6916
rect 3927 6885 3939 6888
rect 3881 6879 3939 6885
rect 1486 6808 1492 6860
rect 1544 6808 1550 6860
rect 1756 6851 1814 6857
rect 1756 6817 1768 6851
rect 1802 6848 1814 6851
rect 2038 6848 2044 6860
rect 1802 6820 2044 6848
rect 1802 6817 1814 6820
rect 1756 6811 1814 6817
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 2314 6808 2320 6860
rect 2372 6848 2378 6860
rect 3510 6848 3516 6860
rect 2372 6820 3516 6848
rect 2372 6808 2378 6820
rect 3510 6808 3516 6820
rect 3568 6808 3574 6860
rect 3988 6848 4016 6888
rect 4798 6848 4804 6860
rect 3988 6820 4804 6848
rect 4798 6808 4804 6820
rect 4856 6848 4862 6860
rect 5000 6857 5028 6888
rect 8110 6876 8116 6928
rect 8168 6916 8174 6928
rect 9490 6916 9496 6928
rect 8168 6888 9496 6916
rect 8168 6876 8174 6888
rect 9490 6876 9496 6888
rect 9548 6876 9554 6928
rect 13464 6916 13492 6956
rect 13909 6953 13921 6956
rect 13955 6984 13967 6987
rect 18325 6987 18383 6993
rect 13955 6956 14964 6984
rect 13955 6953 13967 6956
rect 13909 6947 13967 6953
rect 11992 6888 12480 6916
rect 4985 6851 5043 6857
rect 4985 6848 4997 6851
rect 4856 6820 4997 6848
rect 4856 6808 4862 6820
rect 4985 6817 4997 6820
rect 5031 6817 5043 6851
rect 4985 6811 5043 6817
rect 7736 6851 7794 6857
rect 7736 6817 7748 6851
rect 7782 6848 7794 6851
rect 8294 6848 8300 6860
rect 7782 6820 8300 6848
rect 7782 6817 7794 6820
rect 7736 6811 7794 6817
rect 8294 6808 8300 6820
rect 8352 6808 8358 6860
rect 9125 6851 9183 6857
rect 9125 6817 9137 6851
rect 9171 6848 9183 6851
rect 9171 6820 11100 6848
rect 9171 6817 9183 6820
rect 9125 6811 9183 6817
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6749 3663 6783
rect 3605 6743 3663 6749
rect 2590 6672 2596 6724
rect 2648 6712 2654 6724
rect 2961 6715 3019 6721
rect 2961 6712 2973 6715
rect 2648 6684 2973 6712
rect 2648 6672 2654 6684
rect 2961 6681 2973 6684
rect 3007 6681 3019 6715
rect 2961 6675 3019 6681
rect 3620 6712 3648 6743
rect 6546 6740 6552 6792
rect 6604 6780 6610 6792
rect 7466 6780 7472 6792
rect 6604 6752 7472 6780
rect 6604 6740 6610 6752
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 8478 6740 8484 6792
rect 8536 6780 8542 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8536 6752 8953 6780
rect 8536 6740 8542 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 5350 6712 5356 6724
rect 3620 6684 5356 6712
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3050 6644 3056 6656
rect 2915 6616 3056 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3050 6604 3056 6616
rect 3108 6644 3114 6656
rect 3620 6644 3648 6684
rect 4080 6653 4108 6684
rect 5350 6672 5356 6684
rect 5408 6672 5414 6724
rect 5629 6715 5687 6721
rect 5629 6681 5641 6715
rect 5675 6712 5687 6715
rect 6270 6712 6276 6724
rect 5675 6684 6276 6712
rect 5675 6681 5687 6684
rect 5629 6675 5687 6681
rect 6270 6672 6276 6684
rect 6328 6672 6334 6724
rect 3108 6616 3648 6644
rect 4065 6647 4123 6653
rect 3108 6604 3114 6616
rect 4065 6613 4077 6647
rect 4111 6613 4123 6647
rect 4065 6607 4123 6613
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 4430 6644 4436 6656
rect 4304 6616 4436 6644
rect 4304 6604 4310 6616
rect 4430 6604 4436 6616
rect 4488 6604 4494 6656
rect 5077 6647 5135 6653
rect 5077 6613 5089 6647
rect 5123 6644 5135 6647
rect 5718 6644 5724 6656
rect 5123 6616 5724 6644
rect 5123 6613 5135 6616
rect 5077 6607 5135 6613
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 6178 6604 6184 6656
rect 6236 6644 6242 6656
rect 9140 6644 9168 6811
rect 11072 6792 11100 6820
rect 11422 6808 11428 6860
rect 11480 6808 11486 6860
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 11992 6780 12020 6888
rect 12066 6808 12072 6860
rect 12124 6808 12130 6860
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12250 6848 12256 6860
rect 12207 6820 12256 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12250 6808 12256 6820
rect 12308 6808 12314 6860
rect 12345 6851 12403 6857
rect 12345 6817 12357 6851
rect 12391 6817 12403 6851
rect 12452 6848 12480 6888
rect 13372 6888 13492 6916
rect 13556 6888 14228 6916
rect 13372 6848 13400 6888
rect 12452 6820 13400 6848
rect 13449 6851 13507 6857
rect 12345 6811 12403 6817
rect 13449 6817 13461 6851
rect 13495 6848 13507 6851
rect 13556 6848 13584 6888
rect 13495 6820 13584 6848
rect 13633 6851 13691 6857
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 13633 6817 13645 6851
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 13817 6851 13875 6857
rect 13817 6817 13829 6851
rect 13863 6848 13875 6851
rect 14090 6848 14096 6860
rect 13863 6820 14096 6848
rect 13863 6817 13875 6820
rect 13817 6811 13875 6817
rect 11112 6752 12020 6780
rect 12084 6780 12112 6808
rect 12360 6780 12388 6811
rect 13648 6780 13676 6811
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 14200 6848 14228 6888
rect 14369 6851 14427 6857
rect 14369 6848 14381 6851
rect 14200 6820 14381 6848
rect 14369 6817 14381 6820
rect 14415 6848 14427 6851
rect 14550 6848 14556 6860
rect 14415 6820 14556 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 14550 6808 14556 6820
rect 14608 6808 14614 6860
rect 14734 6808 14740 6860
rect 14792 6848 14798 6860
rect 14829 6851 14887 6857
rect 14829 6848 14841 6851
rect 14792 6820 14841 6848
rect 14792 6808 14798 6820
rect 14829 6817 14841 6820
rect 14875 6817 14887 6851
rect 14936 6848 14964 6956
rect 18325 6953 18337 6987
rect 18371 6984 18383 6987
rect 18874 6984 18880 6996
rect 18371 6956 18880 6984
rect 18371 6953 18383 6956
rect 18325 6947 18383 6953
rect 18874 6944 18880 6956
rect 18932 6944 18938 6996
rect 23198 6944 23204 6996
rect 23256 6944 23262 6996
rect 23750 6944 23756 6996
rect 23808 6984 23814 6996
rect 23937 6987 23995 6993
rect 23937 6984 23949 6987
rect 23808 6956 23949 6984
rect 23808 6944 23814 6956
rect 23937 6953 23949 6956
rect 23983 6953 23995 6987
rect 24305 6987 24363 6993
rect 24305 6984 24317 6987
rect 23937 6947 23995 6953
rect 24044 6956 24317 6984
rect 18141 6919 18199 6925
rect 18141 6885 18153 6919
rect 18187 6885 18199 6919
rect 18141 6879 18199 6885
rect 15562 6848 15568 6860
rect 14936 6820 15568 6848
rect 14829 6811 14887 6817
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 14252 6783 14310 6789
rect 14252 6780 14264 6783
rect 12084 6752 12388 6780
rect 13464 6752 14264 6780
rect 11112 6740 11118 6752
rect 10226 6672 10232 6724
rect 10284 6712 10290 6724
rect 13464 6712 13492 6752
rect 14252 6749 14264 6752
rect 14298 6749 14310 6783
rect 14252 6743 14310 6749
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 15105 6783 15163 6789
rect 15105 6780 15117 6783
rect 14516 6752 15117 6780
rect 14516 6740 14522 6752
rect 15105 6749 15117 6752
rect 15151 6749 15163 6783
rect 18156 6780 18184 6879
rect 18782 6876 18788 6928
rect 18840 6876 18846 6928
rect 20714 6876 20720 6928
rect 20772 6916 20778 6928
rect 21726 6916 21732 6928
rect 20772 6888 21732 6916
rect 20772 6876 20778 6888
rect 21726 6876 21732 6888
rect 21784 6876 21790 6928
rect 22094 6925 22100 6928
rect 22088 6879 22100 6925
rect 22094 6876 22100 6879
rect 22152 6876 22158 6928
rect 23658 6876 23664 6928
rect 23716 6916 23722 6928
rect 24044 6916 24072 6956
rect 24305 6953 24317 6956
rect 24351 6984 24363 6987
rect 24394 6984 24400 6996
rect 24351 6956 24400 6984
rect 24351 6953 24363 6956
rect 24305 6947 24363 6953
rect 24394 6944 24400 6956
rect 24452 6944 24458 6996
rect 25774 6944 25780 6996
rect 25832 6944 25838 6996
rect 23716 6888 24072 6916
rect 24121 6919 24179 6925
rect 23716 6876 23722 6888
rect 24121 6885 24133 6919
rect 24167 6916 24179 6919
rect 24167 6888 24808 6916
rect 24167 6885 24179 6888
rect 24121 6879 24179 6885
rect 18506 6808 18512 6860
rect 18564 6848 18570 6860
rect 18693 6851 18751 6857
rect 18693 6848 18705 6851
rect 18564 6820 18705 6848
rect 18564 6808 18570 6820
rect 18693 6817 18705 6820
rect 18739 6817 18751 6851
rect 18800 6848 18828 6876
rect 24780 6860 24808 6888
rect 25222 6876 25228 6928
rect 25280 6916 25286 6928
rect 25280 6888 25452 6916
rect 25280 6876 25286 6888
rect 18877 6851 18935 6857
rect 18877 6848 18889 6851
rect 18800 6820 18889 6848
rect 18693 6811 18751 6817
rect 18877 6817 18889 6820
rect 18923 6817 18935 6851
rect 18877 6811 18935 6817
rect 20254 6808 20260 6860
rect 20312 6848 20318 6860
rect 20349 6851 20407 6857
rect 20349 6848 20361 6851
rect 20312 6820 20361 6848
rect 20312 6808 20318 6820
rect 20349 6817 20361 6820
rect 20395 6817 20407 6851
rect 20349 6811 20407 6817
rect 18417 6783 18475 6789
rect 18417 6780 18429 6783
rect 18156 6752 18429 6780
rect 15105 6743 15163 6749
rect 18417 6749 18429 6752
rect 18463 6749 18475 6783
rect 18417 6743 18475 6749
rect 18598 6740 18604 6792
rect 18656 6740 18662 6792
rect 18782 6740 18788 6792
rect 18840 6740 18846 6792
rect 19426 6740 19432 6792
rect 19484 6740 19490 6792
rect 20364 6780 20392 6811
rect 20438 6808 20444 6860
rect 20496 6808 20502 6860
rect 20530 6808 20536 6860
rect 20588 6848 20594 6860
rect 20625 6851 20683 6857
rect 20625 6848 20637 6851
rect 20588 6820 20637 6848
rect 20588 6808 20594 6820
rect 20625 6817 20637 6820
rect 20671 6817 20683 6851
rect 20625 6811 20683 6817
rect 20809 6851 20867 6857
rect 20809 6817 20821 6851
rect 20855 6817 20867 6851
rect 20809 6811 20867 6817
rect 20714 6780 20720 6792
rect 20364 6752 20720 6780
rect 20714 6740 20720 6752
rect 20772 6780 20778 6792
rect 20824 6780 20852 6811
rect 23014 6808 23020 6860
rect 23072 6848 23078 6860
rect 24213 6851 24271 6857
rect 24213 6848 24225 6851
rect 23072 6820 24225 6848
rect 23072 6808 23078 6820
rect 24213 6817 24225 6820
rect 24259 6817 24271 6851
rect 24213 6811 24271 6817
rect 20772 6752 20852 6780
rect 21821 6783 21879 6789
rect 20772 6740 20778 6752
rect 21821 6749 21833 6783
rect 21867 6749 21879 6783
rect 24228 6780 24256 6811
rect 24486 6808 24492 6860
rect 24544 6848 24550 6860
rect 24581 6851 24639 6857
rect 24581 6848 24593 6851
rect 24544 6820 24593 6848
rect 24544 6808 24550 6820
rect 24581 6817 24593 6820
rect 24627 6817 24639 6851
rect 24581 6811 24639 6817
rect 24762 6808 24768 6860
rect 24820 6848 24826 6860
rect 25317 6851 25375 6857
rect 25317 6848 25329 6851
rect 24820 6820 25329 6848
rect 24820 6808 24826 6820
rect 25317 6817 25329 6820
rect 25363 6817 25375 6851
rect 25424 6848 25452 6888
rect 25501 6851 25559 6857
rect 25501 6848 25513 6851
rect 25424 6820 25513 6848
rect 25317 6811 25375 6817
rect 25501 6817 25513 6820
rect 25547 6817 25559 6851
rect 25501 6811 25559 6817
rect 25590 6808 25596 6860
rect 25648 6848 25654 6860
rect 26053 6851 26111 6857
rect 25648 6820 25820 6848
rect 25648 6808 25654 6820
rect 24670 6780 24676 6792
rect 24228 6752 24676 6780
rect 21821 6743 21879 6749
rect 10284 6684 13492 6712
rect 13541 6715 13599 6721
rect 10284 6672 10290 6684
rect 13541 6681 13553 6715
rect 13587 6712 13599 6715
rect 14921 6715 14979 6721
rect 14921 6712 14933 6715
rect 13587 6684 14933 6712
rect 13587 6681 13599 6684
rect 13541 6675 13599 6681
rect 14921 6681 14933 6684
rect 14967 6681 14979 6715
rect 14921 6675 14979 6681
rect 17773 6715 17831 6721
rect 17773 6681 17785 6715
rect 17819 6712 17831 6715
rect 18616 6712 18644 6740
rect 19334 6712 19340 6724
rect 17819 6684 18552 6712
rect 18616 6684 19340 6712
rect 17819 6681 17831 6684
rect 17773 6675 17831 6681
rect 6236 6616 9168 6644
rect 9309 6647 9367 6653
rect 6236 6604 6242 6616
rect 9309 6613 9321 6647
rect 9355 6644 9367 6647
rect 11330 6644 11336 6656
rect 9355 6616 11336 6644
rect 9355 6613 9367 6616
rect 9309 6607 9367 6613
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 11422 6604 11428 6656
rect 11480 6644 11486 6656
rect 12529 6647 12587 6653
rect 12529 6644 12541 6647
rect 11480 6616 12541 6644
rect 11480 6604 11486 6616
rect 12529 6613 12541 6616
rect 12575 6613 12587 6647
rect 12529 6607 12587 6613
rect 14093 6647 14151 6653
rect 14093 6613 14105 6647
rect 14139 6644 14151 6647
rect 14274 6644 14280 6656
rect 14139 6616 14280 6644
rect 14139 6613 14151 6616
rect 14093 6607 14151 6613
rect 14274 6604 14280 6616
rect 14332 6604 14338 6656
rect 15289 6647 15347 6653
rect 15289 6613 15301 6647
rect 15335 6644 15347 6647
rect 15562 6644 15568 6656
rect 15335 6616 15568 6644
rect 15335 6613 15347 6616
rect 15289 6607 15347 6613
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 15841 6647 15899 6653
rect 15841 6613 15853 6647
rect 15887 6644 15899 6647
rect 16022 6644 16028 6656
rect 15887 6616 16028 6644
rect 15887 6613 15899 6616
rect 15841 6607 15899 6613
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 18141 6647 18199 6653
rect 18141 6644 18153 6647
rect 18012 6616 18153 6644
rect 18012 6604 18018 6616
rect 18141 6613 18153 6616
rect 18187 6613 18199 6647
rect 18524 6644 18552 6684
rect 19334 6672 19340 6684
rect 19392 6712 19398 6724
rect 20165 6715 20223 6721
rect 20165 6712 20177 6715
rect 19392 6684 20177 6712
rect 19392 6672 19398 6684
rect 20165 6681 20177 6684
rect 20211 6681 20223 6715
rect 20165 6675 20223 6681
rect 19702 6644 19708 6656
rect 18524 6616 19708 6644
rect 18141 6607 18199 6613
rect 19702 6604 19708 6616
rect 19760 6604 19766 6656
rect 20070 6604 20076 6656
rect 20128 6604 20134 6656
rect 20438 6604 20444 6656
rect 20496 6644 20502 6656
rect 20717 6647 20775 6653
rect 20717 6644 20729 6647
rect 20496 6616 20729 6644
rect 20496 6604 20502 6616
rect 20717 6613 20729 6616
rect 20763 6613 20775 6647
rect 21836 6644 21864 6743
rect 24670 6740 24676 6752
rect 24728 6740 24734 6792
rect 25130 6740 25136 6792
rect 25188 6780 25194 6792
rect 25792 6789 25820 6820
rect 26053 6817 26065 6851
rect 26099 6848 26111 6851
rect 26421 6851 26479 6857
rect 26421 6848 26433 6851
rect 26099 6820 26433 6848
rect 26099 6817 26111 6820
rect 26053 6811 26111 6817
rect 26421 6817 26433 6820
rect 26467 6817 26479 6851
rect 26421 6811 26479 6817
rect 25685 6783 25743 6789
rect 25685 6780 25697 6783
rect 25188 6752 25697 6780
rect 25188 6740 25194 6752
rect 25685 6749 25697 6752
rect 25731 6749 25743 6783
rect 25685 6743 25743 6749
rect 25777 6783 25835 6789
rect 25777 6749 25789 6783
rect 25823 6749 25835 6783
rect 25777 6743 25835 6749
rect 25866 6740 25872 6792
rect 25924 6780 25930 6792
rect 26973 6783 27031 6789
rect 26973 6780 26985 6783
rect 25924 6752 26985 6780
rect 25924 6740 25930 6752
rect 26973 6749 26985 6752
rect 27019 6749 27031 6783
rect 26973 6743 27031 6749
rect 23382 6712 23388 6724
rect 23124 6684 23388 6712
rect 23124 6644 23152 6684
rect 23382 6672 23388 6684
rect 23440 6672 23446 6724
rect 24489 6715 24547 6721
rect 24489 6681 24501 6715
rect 24535 6712 24547 6715
rect 25884 6712 25912 6740
rect 24535 6684 25912 6712
rect 24535 6681 24547 6684
rect 24489 6675 24547 6681
rect 21836 6616 23152 6644
rect 20717 6607 20775 6613
rect 24946 6604 24952 6656
rect 25004 6644 25010 6656
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 25004 6616 25973 6644
rect 25004 6604 25010 6616
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 25961 6607 26019 6613
rect 552 6554 27416 6576
rect 552 6502 3756 6554
rect 3808 6502 3820 6554
rect 3872 6502 3884 6554
rect 3936 6502 3948 6554
rect 4000 6502 4012 6554
rect 4064 6502 10472 6554
rect 10524 6502 10536 6554
rect 10588 6502 10600 6554
rect 10652 6502 10664 6554
rect 10716 6502 10728 6554
rect 10780 6502 17188 6554
rect 17240 6502 17252 6554
rect 17304 6502 17316 6554
rect 17368 6502 17380 6554
rect 17432 6502 17444 6554
rect 17496 6502 23904 6554
rect 23956 6502 23968 6554
rect 24020 6502 24032 6554
rect 24084 6502 24096 6554
rect 24148 6502 24160 6554
rect 24212 6502 27416 6554
rect 552 6480 27416 6502
rect 2038 6400 2044 6452
rect 2096 6400 2102 6452
rect 2501 6443 2559 6449
rect 2501 6409 2513 6443
rect 2547 6440 2559 6443
rect 2866 6440 2872 6452
rect 2547 6412 2872 6440
rect 2547 6409 2559 6412
rect 2501 6403 2559 6409
rect 2866 6400 2872 6412
rect 2924 6440 2930 6452
rect 3602 6440 3608 6452
rect 2924 6412 3608 6440
rect 2924 6400 2930 6412
rect 3602 6400 3608 6412
rect 3660 6400 3666 6452
rect 4798 6400 4804 6452
rect 4856 6400 4862 6452
rect 6270 6400 6276 6452
rect 6328 6400 6334 6452
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 9088 6412 11560 6440
rect 9088 6400 9094 6412
rect 9769 6375 9827 6381
rect 9769 6341 9781 6375
rect 9815 6372 9827 6375
rect 10226 6372 10232 6384
rect 9815 6344 10232 6372
rect 9815 6341 9827 6344
rect 9769 6335 9827 6341
rect 10226 6332 10232 6344
rect 10284 6332 10290 6384
rect 11330 6332 11336 6384
rect 11388 6332 11394 6384
rect 11532 6372 11560 6412
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11664 6412 11805 6440
rect 11664 6400 11670 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 14369 6443 14427 6449
rect 14369 6409 14381 6443
rect 14415 6440 14427 6443
rect 14458 6440 14464 6452
rect 14415 6412 14464 6440
rect 14415 6409 14427 6412
rect 14369 6403 14427 6409
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 18509 6443 18567 6449
rect 18509 6409 18521 6443
rect 18555 6440 18567 6443
rect 18690 6440 18696 6452
rect 18555 6412 18696 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 18690 6400 18696 6412
rect 18748 6400 18754 6452
rect 21450 6400 21456 6452
rect 21508 6440 21514 6452
rect 22005 6443 22063 6449
rect 22005 6440 22017 6443
rect 21508 6412 22017 6440
rect 21508 6400 21514 6412
rect 22005 6409 22017 6412
rect 22051 6409 22063 6443
rect 22005 6403 22063 6409
rect 22186 6400 22192 6452
rect 22244 6400 22250 6452
rect 24670 6400 24676 6452
rect 24728 6440 24734 6452
rect 24765 6443 24823 6449
rect 24765 6440 24777 6443
rect 24728 6412 24777 6440
rect 24728 6400 24734 6412
rect 24765 6409 24777 6412
rect 24811 6409 24823 6443
rect 24765 6403 24823 6409
rect 24946 6400 24952 6452
rect 25004 6400 25010 6452
rect 25406 6440 25412 6452
rect 25148 6412 25412 6440
rect 13078 6372 13084 6384
rect 11532 6344 11744 6372
rect 2314 6264 2320 6316
rect 2372 6264 2378 6316
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 2740 6276 3464 6304
rect 2740 6264 2746 6276
rect 2041 6239 2099 6245
rect 2041 6205 2053 6239
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6236 2283 6239
rect 2271 6208 2544 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 2056 6168 2084 6199
rect 2317 6171 2375 6177
rect 2317 6168 2329 6171
rect 2056 6140 2329 6168
rect 2317 6137 2329 6140
rect 2363 6137 2375 6171
rect 2516 6168 2544 6208
rect 2590 6196 2596 6248
rect 2648 6196 2654 6248
rect 2866 6196 2872 6248
rect 2924 6196 2930 6248
rect 3050 6196 3056 6248
rect 3108 6196 3114 6248
rect 3436 6245 3464 6276
rect 10870 6264 10876 6316
rect 10928 6304 10934 6316
rect 10965 6307 11023 6313
rect 10965 6304 10977 6307
rect 10928 6276 10977 6304
rect 10928 6264 10934 6276
rect 10965 6273 10977 6276
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 11054 6264 11060 6316
rect 11112 6264 11118 6316
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6236 3479 6239
rect 4893 6239 4951 6245
rect 4893 6236 4905 6239
rect 3467 6208 4905 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 4893 6205 4905 6208
rect 4939 6236 4951 6239
rect 5534 6236 5540 6248
rect 4939 6208 5540 6236
rect 4939 6205 4951 6208
rect 4893 6199 4951 6205
rect 5534 6196 5540 6208
rect 5592 6236 5598 6248
rect 6546 6236 6552 6248
rect 5592 6208 6552 6236
rect 5592 6196 5598 6208
rect 6546 6196 6552 6208
rect 6604 6196 6610 6248
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 7524 6208 8125 6236
rect 7524 6196 7530 6208
rect 8113 6205 8125 6208
rect 8159 6236 8171 6239
rect 8389 6239 8447 6245
rect 8389 6236 8401 6239
rect 8159 6208 8401 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 8389 6205 8401 6208
rect 8435 6205 8447 6239
rect 8389 6199 8447 6205
rect 10226 6196 10232 6248
rect 10284 6196 10290 6248
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6205 10379 6239
rect 10321 6199 10379 6205
rect 2685 6171 2743 6177
rect 2685 6168 2697 6171
rect 2516 6140 2697 6168
rect 2317 6131 2375 6137
rect 2685 6137 2697 6140
rect 2731 6168 2743 6171
rect 3326 6168 3332 6180
rect 2731 6140 3332 6168
rect 2731 6137 2743 6140
rect 2685 6131 2743 6137
rect 3326 6128 3332 6140
rect 3384 6128 3390 6180
rect 3688 6171 3746 6177
rect 3688 6137 3700 6171
rect 3734 6168 3746 6171
rect 4338 6168 4344 6180
rect 3734 6140 4344 6168
rect 3734 6137 3746 6140
rect 3688 6131 3746 6137
rect 4338 6128 4344 6140
rect 4396 6128 4402 6180
rect 5166 6177 5172 6180
rect 5160 6131 5172 6177
rect 5166 6128 5172 6131
rect 5224 6128 5230 6180
rect 6362 6128 6368 6180
rect 6420 6128 6426 6180
rect 8662 6177 8668 6180
rect 8656 6131 8668 6177
rect 8662 6128 8668 6131
rect 8720 6128 8726 6180
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 9030 6100 9036 6112
rect 4580 6072 9036 6100
rect 4580 6060 4586 6072
rect 9030 6060 9036 6072
rect 9088 6060 9094 6112
rect 9122 6060 9128 6112
rect 9180 6100 9186 6112
rect 10045 6103 10103 6109
rect 10045 6100 10057 6103
rect 9180 6072 10057 6100
rect 9180 6060 9186 6072
rect 10045 6069 10057 6072
rect 10091 6100 10103 6103
rect 10226 6100 10232 6112
rect 10091 6072 10232 6100
rect 10091 6069 10103 6072
rect 10045 6063 10103 6069
rect 10226 6060 10232 6072
rect 10284 6100 10290 6112
rect 10336 6100 10364 6199
rect 10410 6196 10416 6248
rect 10468 6196 10474 6248
rect 10594 6196 10600 6248
rect 10652 6196 10658 6248
rect 10689 6239 10747 6245
rect 10689 6205 10701 6239
rect 10735 6236 10747 6239
rect 11072 6236 11100 6264
rect 11621 6249 11679 6255
rect 10735 6208 11100 6236
rect 11149 6239 11207 6245
rect 10735 6205 10747 6208
rect 10689 6199 10747 6205
rect 11149 6205 11161 6239
rect 11195 6205 11207 6239
rect 11149 6199 11207 6205
rect 11241 6239 11299 6245
rect 11241 6205 11253 6239
rect 11287 6205 11299 6239
rect 11241 6199 11299 6205
rect 10870 6128 10876 6180
rect 10928 6128 10934 6180
rect 10284 6072 10364 6100
rect 11164 6100 11192 6199
rect 11257 6168 11285 6199
rect 11422 6196 11428 6248
rect 11480 6236 11486 6248
rect 11480 6208 11524 6236
rect 11621 6215 11633 6249
rect 11667 6246 11679 6249
rect 11716 6246 11744 6344
rect 12452 6344 13084 6372
rect 12452 6313 12480 6344
rect 13078 6332 13084 6344
rect 13136 6372 13142 6384
rect 13633 6375 13691 6381
rect 13633 6372 13645 6375
rect 13136 6344 13645 6372
rect 13136 6332 13142 6344
rect 13633 6341 13645 6344
rect 13679 6341 13691 6375
rect 13633 6335 13691 6341
rect 15838 6332 15844 6384
rect 15896 6332 15902 6384
rect 19518 6372 19524 6384
rect 18524 6344 19524 6372
rect 18524 6316 18552 6344
rect 19518 6332 19524 6344
rect 19576 6332 19582 6384
rect 19702 6332 19708 6384
rect 19760 6372 19766 6384
rect 23014 6372 23020 6384
rect 19760 6344 23020 6372
rect 19760 6332 19766 6344
rect 23014 6332 23020 6344
rect 23072 6332 23078 6384
rect 23382 6332 23388 6384
rect 23440 6372 23446 6384
rect 25148 6372 25176 6412
rect 25406 6400 25412 6412
rect 25464 6400 25470 6452
rect 25866 6400 25872 6452
rect 25924 6440 25930 6452
rect 26513 6443 26571 6449
rect 26513 6440 26525 6443
rect 25924 6412 26525 6440
rect 25924 6400 25930 6412
rect 26513 6409 26525 6412
rect 26559 6409 26571 6443
rect 26513 6403 26571 6409
rect 23440 6344 25176 6372
rect 23440 6332 23446 6344
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6304 15807 6307
rect 16298 6304 16304 6316
rect 15795 6276 16304 6304
rect 15795 6273 15807 6276
rect 15749 6267 15807 6273
rect 16298 6264 16304 6276
rect 16356 6304 16362 6316
rect 17129 6307 17187 6313
rect 17129 6304 17141 6307
rect 16356 6276 17141 6304
rect 16356 6264 16362 6276
rect 17129 6273 17141 6276
rect 17175 6273 17187 6307
rect 17129 6267 17187 6273
rect 11667 6218 11744 6246
rect 11667 6215 11679 6218
rect 11621 6209 11679 6215
rect 11480 6196 11486 6208
rect 11882 6196 11888 6248
rect 11940 6236 11946 6248
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 11940 6208 12173 6236
rect 11940 6196 11946 6208
rect 12161 6205 12173 6208
rect 12207 6236 12219 6239
rect 12986 6236 12992 6248
rect 12207 6208 12992 6236
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 12986 6196 12992 6208
rect 13044 6196 13050 6248
rect 13817 6239 13875 6245
rect 13817 6205 13829 6239
rect 13863 6236 13875 6239
rect 14090 6236 14096 6248
rect 13863 6208 14096 6236
rect 13863 6205 13875 6208
rect 13817 6199 13875 6205
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 16117 6239 16175 6245
rect 16117 6205 16129 6239
rect 16163 6236 16175 6239
rect 16390 6236 16396 6248
rect 16163 6208 16396 6236
rect 16163 6205 16175 6208
rect 16117 6199 16175 6205
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 16853 6239 16911 6245
rect 16853 6205 16865 6239
rect 16899 6205 16911 6239
rect 16853 6199 16911 6205
rect 11257 6140 11376 6168
rect 11238 6100 11244 6112
rect 11164 6072 11244 6100
rect 10284 6060 10290 6072
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 11348 6100 11376 6140
rect 14918 6128 14924 6180
rect 14976 6168 14982 6180
rect 15482 6171 15540 6177
rect 15482 6168 15494 6171
rect 14976 6140 15494 6168
rect 14976 6128 14982 6140
rect 15482 6137 15494 6140
rect 15528 6137 15540 6171
rect 15482 6131 15540 6137
rect 15841 6171 15899 6177
rect 15841 6137 15853 6171
rect 15887 6137 15899 6171
rect 15841 6131 15899 6137
rect 11974 6100 11980 6112
rect 11348 6072 11980 6100
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12253 6103 12311 6109
rect 12253 6069 12265 6103
rect 12299 6100 12311 6103
rect 13538 6100 13544 6112
rect 12299 6072 13544 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 13538 6060 13544 6072
rect 13596 6060 13602 6112
rect 15286 6060 15292 6112
rect 15344 6100 15350 6112
rect 15856 6100 15884 6131
rect 15344 6072 15884 6100
rect 15344 6060 15350 6072
rect 16022 6060 16028 6112
rect 16080 6100 16086 6112
rect 16482 6100 16488 6112
rect 16080 6072 16488 6100
rect 16080 6060 16086 6072
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 16868 6100 16896 6199
rect 17034 6196 17040 6248
rect 17092 6196 17098 6248
rect 17144 6236 17172 6267
rect 18506 6264 18512 6316
rect 18564 6264 18570 6316
rect 19334 6264 19340 6316
rect 19392 6304 19398 6316
rect 21821 6307 21879 6313
rect 21821 6304 21833 6307
rect 19392 6276 21833 6304
rect 19392 6264 19398 6276
rect 21821 6273 21833 6276
rect 21867 6273 21879 6307
rect 22833 6307 22891 6313
rect 22833 6304 22845 6307
rect 21821 6267 21879 6273
rect 22066 6276 22845 6304
rect 17954 6236 17960 6248
rect 17144 6208 17960 6236
rect 17954 6196 17960 6208
rect 18012 6236 18018 6248
rect 18693 6239 18751 6245
rect 18693 6236 18705 6239
rect 18012 6208 18705 6236
rect 18012 6196 18018 6208
rect 18693 6205 18705 6208
rect 18739 6236 18751 6239
rect 19242 6236 19248 6248
rect 18739 6208 19248 6236
rect 18739 6205 18751 6208
rect 18693 6199 18751 6205
rect 19242 6196 19248 6208
rect 19300 6196 19306 6248
rect 20441 6239 20499 6245
rect 20441 6205 20453 6239
rect 20487 6236 20499 6239
rect 20622 6236 20628 6248
rect 20487 6208 20628 6236
rect 20487 6205 20499 6208
rect 20441 6199 20499 6205
rect 20622 6196 20628 6208
rect 20680 6196 20686 6248
rect 20714 6196 20720 6248
rect 20772 6196 20778 6248
rect 20993 6239 21051 6245
rect 20993 6236 21005 6239
rect 20824 6208 21005 6236
rect 16945 6171 17003 6177
rect 16945 6137 16957 6171
rect 16991 6168 17003 6171
rect 17374 6171 17432 6177
rect 17374 6168 17386 6171
rect 16991 6140 17386 6168
rect 16991 6137 17003 6140
rect 16945 6131 17003 6137
rect 17374 6137 17386 6140
rect 17420 6137 17432 6171
rect 17374 6131 17432 6137
rect 18874 6128 18880 6180
rect 18932 6168 18938 6180
rect 20530 6168 20536 6180
rect 18932 6140 20536 6168
rect 18932 6128 18938 6140
rect 20530 6128 20536 6140
rect 20588 6128 20594 6180
rect 18046 6100 18052 6112
rect 16868 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 20346 6060 20352 6112
rect 20404 6100 20410 6112
rect 20824 6100 20852 6208
rect 20993 6205 21005 6208
rect 21039 6205 21051 6239
rect 20993 6199 21051 6205
rect 21637 6239 21695 6245
rect 21637 6205 21649 6239
rect 21683 6236 21695 6239
rect 21729 6239 21787 6245
rect 21729 6236 21741 6239
rect 21683 6208 21741 6236
rect 21683 6205 21695 6208
rect 21637 6199 21695 6205
rect 21729 6205 21741 6208
rect 21775 6205 21787 6239
rect 21729 6199 21787 6205
rect 21082 6128 21088 6180
rect 21140 6168 21146 6180
rect 22066 6168 22094 6276
rect 22833 6273 22845 6276
rect 22879 6304 22891 6307
rect 23566 6304 23572 6316
rect 22879 6276 23572 6304
rect 22879 6273 22891 6276
rect 22833 6267 22891 6273
rect 23566 6264 23572 6276
rect 23624 6264 23630 6316
rect 24394 6264 24400 6316
rect 24452 6304 24458 6316
rect 25148 6313 25176 6344
rect 25133 6307 25191 6313
rect 24452 6276 24624 6304
rect 24452 6264 24458 6276
rect 23109 6239 23167 6245
rect 23109 6205 23121 6239
rect 23155 6236 23167 6239
rect 23845 6239 23903 6245
rect 23845 6236 23857 6239
rect 23155 6208 23857 6236
rect 23155 6205 23167 6208
rect 23109 6199 23167 6205
rect 23845 6205 23857 6208
rect 23891 6205 23903 6239
rect 23845 6199 23903 6205
rect 21140 6140 22094 6168
rect 22173 6171 22231 6177
rect 21140 6128 21146 6140
rect 22173 6137 22185 6171
rect 22219 6168 22231 6171
rect 22278 6168 22284 6180
rect 22219 6140 22284 6168
rect 22219 6137 22231 6140
rect 22173 6131 22231 6137
rect 22278 6128 22284 6140
rect 22336 6128 22342 6180
rect 22370 6128 22376 6180
rect 22428 6128 22434 6180
rect 24596 6177 24624 6276
rect 25133 6273 25145 6307
rect 25179 6273 25191 6307
rect 25133 6267 25191 6273
rect 25400 6239 25458 6245
rect 25400 6205 25412 6239
rect 25446 6236 25458 6239
rect 25682 6236 25688 6248
rect 25446 6208 25688 6236
rect 25446 6205 25458 6208
rect 25400 6199 25458 6205
rect 25682 6196 25688 6208
rect 25740 6196 25746 6248
rect 24581 6171 24639 6177
rect 24581 6137 24593 6171
rect 24627 6137 24639 6171
rect 24581 6131 24639 6137
rect 24762 6128 24768 6180
rect 24820 6177 24826 6180
rect 24820 6171 24839 6177
rect 24827 6137 24839 6171
rect 24820 6131 24839 6137
rect 24820 6128 24826 6131
rect 20404 6072 20852 6100
rect 20901 6103 20959 6109
rect 20404 6060 20410 6072
rect 20901 6069 20913 6103
rect 20947 6100 20959 6103
rect 21450 6100 21456 6112
rect 20947 6072 21456 6100
rect 20947 6069 20959 6072
rect 20901 6063 20959 6069
rect 21450 6060 21456 6072
rect 21508 6060 21514 6112
rect 22554 6060 22560 6112
rect 22612 6100 22618 6112
rect 22833 6103 22891 6109
rect 22833 6100 22845 6103
rect 22612 6072 22845 6100
rect 22612 6060 22618 6072
rect 22833 6069 22845 6072
rect 22879 6069 22891 6103
rect 22833 6063 22891 6069
rect 552 6010 27576 6032
rect 552 5958 7114 6010
rect 7166 5958 7178 6010
rect 7230 5958 7242 6010
rect 7294 5958 7306 6010
rect 7358 5958 7370 6010
rect 7422 5958 13830 6010
rect 13882 5958 13894 6010
rect 13946 5958 13958 6010
rect 14010 5958 14022 6010
rect 14074 5958 14086 6010
rect 14138 5958 20546 6010
rect 20598 5958 20610 6010
rect 20662 5958 20674 6010
rect 20726 5958 20738 6010
rect 20790 5958 20802 6010
rect 20854 5958 27262 6010
rect 27314 5958 27326 6010
rect 27378 5958 27390 6010
rect 27442 5958 27454 6010
rect 27506 5958 27518 6010
rect 27570 5958 27576 6010
rect 552 5936 27576 5958
rect 6457 5899 6515 5905
rect 6457 5896 6469 5899
rect 5460 5868 6469 5896
rect 4985 5831 5043 5837
rect 4985 5797 4997 5831
rect 5031 5828 5043 5831
rect 5031 5800 5396 5828
rect 5031 5797 5043 5800
rect 4985 5791 5043 5797
rect 4246 5720 4252 5772
rect 4304 5760 4310 5772
rect 5368 5769 5396 5800
rect 5169 5763 5227 5769
rect 5169 5760 5181 5763
rect 4304 5732 5181 5760
rect 4304 5720 4310 5732
rect 5169 5729 5181 5732
rect 5215 5729 5227 5763
rect 5169 5723 5227 5729
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5729 5319 5763
rect 5261 5723 5319 5729
rect 5353 5763 5411 5769
rect 5353 5729 5365 5763
rect 5399 5729 5411 5763
rect 5353 5723 5411 5729
rect 3510 5652 3516 5704
rect 3568 5692 3574 5704
rect 4985 5695 5043 5701
rect 4985 5692 4997 5695
rect 3568 5664 4997 5692
rect 3568 5652 3574 5664
rect 4985 5661 4997 5664
rect 5031 5661 5043 5695
rect 5276 5692 5304 5723
rect 5460 5692 5488 5868
rect 6457 5865 6469 5868
rect 6503 5896 6515 5899
rect 8478 5896 8484 5908
rect 6503 5868 8484 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 8662 5856 8668 5908
rect 8720 5856 8726 5908
rect 10410 5856 10416 5908
rect 10468 5896 10474 5908
rect 10468 5868 13216 5896
rect 10468 5856 10474 5868
rect 5718 5828 5724 5840
rect 5552 5800 5724 5828
rect 5552 5769 5580 5800
rect 5718 5788 5724 5800
rect 5776 5828 5782 5840
rect 13188 5837 13216 5868
rect 13998 5856 14004 5908
rect 14056 5896 14062 5908
rect 14458 5896 14464 5908
rect 14056 5868 14464 5896
rect 14056 5856 14062 5868
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 14918 5856 14924 5908
rect 14976 5856 14982 5908
rect 17034 5856 17040 5908
rect 17092 5896 17098 5908
rect 17313 5899 17371 5905
rect 17313 5896 17325 5899
rect 17092 5868 17325 5896
rect 17092 5856 17098 5868
rect 17313 5865 17325 5868
rect 17359 5865 17371 5899
rect 17313 5859 17371 5865
rect 17681 5899 17739 5905
rect 17681 5865 17693 5899
rect 17727 5896 17739 5899
rect 18046 5896 18052 5908
rect 17727 5868 18052 5896
rect 17727 5865 17739 5868
rect 17681 5859 17739 5865
rect 18046 5856 18052 5868
rect 18104 5896 18110 5908
rect 18874 5896 18880 5908
rect 18104 5868 18880 5896
rect 18104 5856 18110 5868
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 20346 5856 20352 5908
rect 20404 5896 20410 5908
rect 20809 5899 20867 5905
rect 20809 5896 20821 5899
rect 20404 5868 20821 5896
rect 20404 5856 20410 5868
rect 20809 5865 20821 5868
rect 20855 5865 20867 5899
rect 22094 5896 22100 5908
rect 20809 5859 20867 5865
rect 21652 5868 22100 5896
rect 13173 5831 13231 5837
rect 5776 5800 13124 5828
rect 5776 5788 5782 5800
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5729 5595 5763
rect 5537 5723 5595 5729
rect 5905 5763 5963 5769
rect 5905 5729 5917 5763
rect 5951 5760 5963 5763
rect 6270 5760 6276 5772
rect 5951 5732 6276 5760
rect 5951 5729 5963 5732
rect 5905 5723 5963 5729
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 8481 5763 8539 5769
rect 8481 5729 8493 5763
rect 8527 5760 8539 5763
rect 8570 5760 8576 5772
rect 8527 5732 8576 5760
rect 8527 5729 8539 5732
rect 8481 5723 8539 5729
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 8846 5720 8852 5772
rect 8904 5760 8910 5772
rect 8941 5763 8999 5769
rect 8941 5760 8953 5763
rect 8904 5732 8953 5760
rect 8904 5720 8910 5732
rect 8941 5729 8953 5732
rect 8987 5729 8999 5763
rect 8941 5723 8999 5729
rect 9122 5720 9128 5772
rect 9180 5720 9186 5772
rect 10962 5720 10968 5772
rect 11020 5720 11026 5772
rect 11054 5720 11060 5772
rect 11112 5720 11118 5772
rect 11232 5763 11290 5769
rect 11232 5729 11244 5763
rect 11278 5760 11290 5763
rect 11606 5760 11612 5772
rect 11278 5732 11612 5760
rect 11278 5729 11290 5732
rect 11232 5723 11290 5729
rect 11606 5720 11612 5732
rect 11664 5720 11670 5772
rect 5276 5664 5488 5692
rect 4985 5655 5043 5661
rect 5000 5624 5028 5655
rect 8202 5652 8208 5704
rect 8260 5652 8266 5704
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 11072 5692 11100 5720
rect 12526 5692 12532 5704
rect 10928 5664 11100 5692
rect 12360 5664 12532 5692
rect 10928 5652 10934 5664
rect 10778 5624 10784 5636
rect 5000 5596 10784 5624
rect 10778 5584 10784 5596
rect 10836 5584 10842 5636
rect 12360 5633 12388 5664
rect 12526 5652 12532 5664
rect 12584 5692 12590 5704
rect 12989 5695 13047 5701
rect 12989 5692 13001 5695
rect 12584 5664 13001 5692
rect 12584 5652 12590 5664
rect 12989 5661 13001 5664
rect 13035 5661 13047 5695
rect 13096 5692 13124 5800
rect 13173 5797 13185 5831
rect 13219 5797 13231 5831
rect 14550 5828 14556 5840
rect 13173 5791 13231 5797
rect 13648 5800 14556 5828
rect 13648 5769 13676 5800
rect 14550 5788 14556 5800
rect 14608 5788 14614 5840
rect 16574 5828 16580 5840
rect 14844 5800 16580 5828
rect 13633 5763 13691 5769
rect 13633 5729 13645 5763
rect 13679 5729 13691 5763
rect 13633 5723 13691 5729
rect 13998 5720 14004 5772
rect 14056 5720 14062 5772
rect 14182 5720 14188 5772
rect 14240 5720 14246 5772
rect 14274 5720 14280 5772
rect 14332 5760 14338 5772
rect 14458 5760 14464 5772
rect 14332 5732 14464 5760
rect 14332 5720 14338 5732
rect 14458 5720 14464 5732
rect 14516 5760 14522 5772
rect 14844 5769 14872 5800
rect 16574 5788 16580 5800
rect 16632 5828 16638 5840
rect 17494 5828 17500 5840
rect 16632 5800 17500 5828
rect 16632 5788 16638 5800
rect 17494 5788 17500 5800
rect 17552 5788 17558 5840
rect 18141 5831 18199 5837
rect 18141 5828 18153 5831
rect 17604 5800 18153 5828
rect 14737 5763 14795 5769
rect 14737 5760 14749 5763
rect 14516 5732 14749 5760
rect 14516 5720 14522 5732
rect 14737 5729 14749 5732
rect 14783 5729 14795 5763
rect 14737 5723 14795 5729
rect 14829 5763 14887 5769
rect 14829 5729 14841 5763
rect 14875 5729 14887 5763
rect 14829 5723 14887 5729
rect 15013 5763 15071 5769
rect 15013 5729 15025 5763
rect 15059 5760 15071 5763
rect 15838 5760 15844 5772
rect 15059 5732 15844 5760
rect 15059 5729 15071 5732
rect 15013 5723 15071 5729
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 17604 5769 17632 5800
rect 18141 5797 18153 5800
rect 18187 5797 18199 5831
rect 18141 5791 18199 5797
rect 19696 5831 19754 5837
rect 19696 5797 19708 5831
rect 19742 5828 19754 5831
rect 20070 5828 20076 5840
rect 19742 5800 20076 5828
rect 19742 5797 19754 5800
rect 19696 5791 19754 5797
rect 20070 5788 20076 5800
rect 20128 5788 20134 5840
rect 20622 5788 20628 5840
rect 20680 5828 20686 5840
rect 21652 5837 21680 5868
rect 22094 5856 22100 5868
rect 22152 5896 22158 5908
rect 22370 5896 22376 5908
rect 22152 5868 22376 5896
rect 22152 5856 22158 5868
rect 22370 5856 22376 5868
rect 22428 5896 22434 5908
rect 23290 5896 23296 5908
rect 22428 5868 23296 5896
rect 22428 5856 22434 5868
rect 23290 5856 23296 5868
rect 23348 5856 23354 5908
rect 23658 5856 23664 5908
rect 23716 5896 23722 5908
rect 24029 5899 24087 5905
rect 24029 5896 24041 5899
rect 23716 5868 24041 5896
rect 23716 5856 23722 5868
rect 24029 5865 24041 5868
rect 24075 5896 24087 5899
rect 24394 5896 24400 5908
rect 24075 5868 24400 5896
rect 24075 5865 24087 5868
rect 24029 5859 24087 5865
rect 24394 5856 24400 5868
rect 24452 5856 24458 5908
rect 24581 5899 24639 5905
rect 24581 5865 24593 5899
rect 24627 5896 24639 5899
rect 25130 5896 25136 5908
rect 24627 5868 25136 5896
rect 24627 5865 24639 5868
rect 24581 5859 24639 5865
rect 25130 5856 25136 5868
rect 25188 5856 25194 5908
rect 21421 5831 21479 5837
rect 21421 5828 21433 5831
rect 20680 5800 21433 5828
rect 20680 5788 20686 5800
rect 21421 5797 21433 5800
rect 21467 5797 21479 5831
rect 21421 5791 21479 5797
rect 21637 5831 21695 5837
rect 21637 5797 21649 5831
rect 21683 5797 21695 5831
rect 23382 5828 23388 5840
rect 21637 5791 21695 5797
rect 22664 5800 23388 5828
rect 22664 5772 22692 5800
rect 23382 5788 23388 5800
rect 23440 5788 23446 5840
rect 25406 5788 25412 5840
rect 25464 5828 25470 5840
rect 25464 5800 26004 5828
rect 25464 5788 25470 5800
rect 17589 5763 17647 5769
rect 17589 5729 17601 5763
rect 17635 5729 17647 5763
rect 17589 5723 17647 5729
rect 17865 5763 17923 5769
rect 17865 5729 17877 5763
rect 17911 5729 17923 5763
rect 17865 5723 17923 5729
rect 18049 5763 18107 5769
rect 18049 5729 18061 5763
rect 18095 5760 18107 5763
rect 18690 5760 18696 5772
rect 18095 5732 18696 5760
rect 18095 5729 18107 5732
rect 18049 5723 18107 5729
rect 13096 5664 16620 5692
rect 12989 5655 13047 5661
rect 12345 5627 12403 5633
rect 12345 5593 12357 5627
rect 12391 5593 12403 5627
rect 12345 5587 12403 5593
rect 12434 5584 12440 5636
rect 12492 5584 12498 5636
rect 16592 5624 16620 5664
rect 17310 5652 17316 5704
rect 17368 5652 17374 5704
rect 17880 5692 17908 5723
rect 18690 5720 18696 5732
rect 18748 5720 18754 5772
rect 19242 5720 19248 5772
rect 19300 5760 19306 5772
rect 19429 5763 19487 5769
rect 19429 5760 19441 5763
rect 19300 5732 19441 5760
rect 19300 5720 19306 5732
rect 19429 5729 19441 5732
rect 19475 5729 19487 5763
rect 19429 5723 19487 5729
rect 21085 5763 21143 5769
rect 21085 5729 21097 5763
rect 21131 5760 21143 5763
rect 21131 5732 21312 5760
rect 21131 5729 21143 5732
rect 21085 5723 21143 5729
rect 18506 5692 18512 5704
rect 17512 5664 18512 5692
rect 17512 5633 17540 5664
rect 18506 5652 18512 5664
rect 18564 5652 18570 5704
rect 17497 5627 17555 5633
rect 17497 5624 17509 5627
rect 16592 5596 17509 5624
rect 17497 5593 17509 5596
rect 17543 5593 17555 5627
rect 17497 5587 17555 5593
rect 17586 5584 17592 5636
rect 17644 5624 17650 5636
rect 18782 5624 18788 5636
rect 17644 5596 18788 5624
rect 17644 5584 17650 5596
rect 18782 5584 18788 5596
rect 18840 5584 18846 5636
rect 21082 5624 21088 5636
rect 20824 5596 21088 5624
rect 5166 5516 5172 5568
rect 5224 5556 5230 5568
rect 5353 5559 5411 5565
rect 5353 5556 5365 5559
rect 5224 5528 5365 5556
rect 5224 5516 5230 5528
rect 5353 5525 5365 5528
rect 5399 5525 5411 5559
rect 5353 5519 5411 5525
rect 8297 5559 8355 5565
rect 8297 5525 8309 5559
rect 8343 5556 8355 5559
rect 8757 5559 8815 5565
rect 8757 5556 8769 5559
rect 8343 5528 8769 5556
rect 8343 5525 8355 5528
rect 8297 5519 8355 5525
rect 8757 5525 8769 5528
rect 8803 5525 8815 5559
rect 8757 5519 8815 5525
rect 9030 5516 9036 5568
rect 9088 5556 9094 5568
rect 14458 5556 14464 5568
rect 9088 5528 14464 5556
rect 9088 5516 9094 5528
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 14553 5559 14611 5565
rect 14553 5525 14565 5559
rect 14599 5556 14611 5559
rect 15930 5556 15936 5568
rect 14599 5528 15936 5556
rect 14599 5525 14611 5528
rect 14553 5519 14611 5525
rect 15930 5516 15936 5528
rect 15988 5516 15994 5568
rect 17310 5516 17316 5568
rect 17368 5556 17374 5568
rect 20824 5556 20852 5596
rect 21082 5584 21088 5596
rect 21140 5584 21146 5636
rect 21284 5633 21312 5732
rect 22370 5720 22376 5772
rect 22428 5720 22434 5772
rect 22554 5720 22560 5772
rect 22612 5720 22618 5772
rect 22646 5720 22652 5772
rect 22704 5720 22710 5772
rect 22905 5763 22963 5769
rect 22905 5760 22917 5763
rect 22756 5732 22917 5760
rect 22465 5695 22523 5701
rect 22465 5661 22477 5695
rect 22511 5692 22523 5695
rect 22756 5692 22784 5732
rect 22905 5729 22917 5732
rect 22951 5729 22963 5763
rect 22905 5723 22963 5729
rect 24486 5720 24492 5772
rect 24544 5720 24550 5772
rect 25682 5720 25688 5772
rect 25740 5769 25746 5772
rect 25976 5769 26004 5800
rect 25740 5723 25752 5769
rect 25961 5763 26019 5769
rect 25961 5729 25973 5763
rect 26007 5729 26019 5763
rect 25961 5723 26019 5729
rect 25740 5720 25746 5723
rect 22511 5664 22784 5692
rect 22511 5661 22523 5664
rect 22465 5655 22523 5661
rect 21269 5627 21327 5633
rect 21269 5593 21281 5627
rect 21315 5593 21327 5627
rect 21269 5587 21327 5593
rect 17368 5528 20852 5556
rect 20901 5559 20959 5565
rect 17368 5516 17374 5528
rect 20901 5525 20913 5559
rect 20947 5556 20959 5559
rect 20990 5556 20996 5568
rect 20947 5528 20996 5556
rect 20947 5525 20959 5528
rect 20901 5519 20959 5525
rect 20990 5516 20996 5528
rect 21048 5516 21054 5568
rect 21450 5516 21456 5568
rect 21508 5516 21514 5568
rect 24302 5516 24308 5568
rect 24360 5556 24366 5568
rect 24397 5559 24455 5565
rect 24397 5556 24409 5559
rect 24360 5528 24409 5556
rect 24360 5516 24366 5528
rect 24397 5525 24409 5528
rect 24443 5525 24455 5559
rect 24397 5519 24455 5525
rect 552 5466 27416 5488
rect 552 5414 3756 5466
rect 3808 5414 3820 5466
rect 3872 5414 3884 5466
rect 3936 5414 3948 5466
rect 4000 5414 4012 5466
rect 4064 5414 10472 5466
rect 10524 5414 10536 5466
rect 10588 5414 10600 5466
rect 10652 5414 10664 5466
rect 10716 5414 10728 5466
rect 10780 5414 17188 5466
rect 17240 5414 17252 5466
rect 17304 5414 17316 5466
rect 17368 5414 17380 5466
rect 17432 5414 17444 5466
rect 17496 5414 23904 5466
rect 23956 5414 23968 5466
rect 24020 5414 24032 5466
rect 24084 5414 24096 5466
rect 24148 5414 24160 5466
rect 24212 5414 27416 5466
rect 552 5392 27416 5414
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 5626 5352 5632 5364
rect 4120 5324 5632 5352
rect 4120 5312 4126 5324
rect 5626 5312 5632 5324
rect 5684 5352 5690 5364
rect 7190 5352 7196 5364
rect 5684 5324 7196 5352
rect 5684 5312 5690 5324
rect 7190 5312 7196 5324
rect 7248 5352 7254 5364
rect 7466 5352 7472 5364
rect 7248 5324 7472 5352
rect 7248 5312 7254 5324
rect 7466 5312 7472 5324
rect 7524 5352 7530 5364
rect 9950 5352 9956 5364
rect 7524 5324 9956 5352
rect 7524 5312 7530 5324
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 10137 5355 10195 5361
rect 10137 5321 10149 5355
rect 10183 5352 10195 5355
rect 10962 5352 10968 5364
rect 10183 5324 10968 5352
rect 10183 5321 10195 5324
rect 10137 5315 10195 5321
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11701 5355 11759 5361
rect 11701 5321 11713 5355
rect 11747 5352 11759 5355
rect 11790 5352 11796 5364
rect 11747 5324 11796 5352
rect 11747 5321 11759 5324
rect 11701 5315 11759 5321
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 13538 5312 13544 5364
rect 13596 5312 13602 5364
rect 14369 5355 14427 5361
rect 14369 5321 14381 5355
rect 14415 5352 14427 5355
rect 14642 5352 14648 5364
rect 14415 5324 14648 5352
rect 14415 5321 14427 5324
rect 14369 5315 14427 5321
rect 14642 5312 14648 5324
rect 14700 5312 14706 5364
rect 15102 5312 15108 5364
rect 15160 5352 15166 5364
rect 19889 5355 19947 5361
rect 15160 5324 16436 5352
rect 15160 5312 15166 5324
rect 7650 5244 7656 5296
rect 7708 5284 7714 5296
rect 9968 5284 9996 5312
rect 10870 5284 10876 5296
rect 7708 5256 9720 5284
rect 9968 5256 10876 5284
rect 7708 5244 7714 5256
rect 5350 5176 5356 5228
rect 5408 5216 5414 5228
rect 9033 5219 9091 5225
rect 9033 5216 9045 5219
rect 5408 5188 9045 5216
rect 5408 5176 5414 5188
rect 9033 5185 9045 5188
rect 9079 5185 9091 5219
rect 9033 5179 9091 5185
rect 9122 5176 9128 5228
rect 9180 5216 9186 5228
rect 9180 5188 9628 5216
rect 9180 5176 9186 5188
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5148 4307 5151
rect 5534 5148 5540 5160
rect 4295 5120 5540 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 5902 5108 5908 5160
rect 5960 5108 5966 5160
rect 6457 5151 6515 5157
rect 6457 5117 6469 5151
rect 6503 5148 6515 5151
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6503 5120 6837 5148
rect 6503 5117 6515 5120
rect 6457 5111 6515 5117
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 6914 5108 6920 5160
rect 6972 5108 6978 5160
rect 7009 5151 7067 5157
rect 7009 5117 7021 5151
rect 7055 5117 7067 5151
rect 7009 5111 7067 5117
rect 4516 5083 4574 5089
rect 4516 5049 4528 5083
rect 4562 5080 4574 5083
rect 6549 5083 6607 5089
rect 6549 5080 6561 5083
rect 4562 5052 6561 5080
rect 4562 5049 4574 5052
rect 4516 5043 4574 5049
rect 6549 5049 6561 5052
rect 6595 5049 6607 5083
rect 7024 5080 7052 5111
rect 7190 5108 7196 5160
rect 7248 5108 7254 5160
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 8018 5148 8024 5160
rect 7975 5120 8024 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 8113 5151 8171 5157
rect 8113 5117 8125 5151
rect 8159 5148 8171 5151
rect 8294 5148 8300 5160
rect 8159 5120 8300 5148
rect 8159 5117 8171 5120
rect 8113 5111 8171 5117
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 8573 5151 8631 5157
rect 8573 5117 8585 5151
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 8665 5151 8723 5157
rect 8665 5117 8677 5151
rect 8711 5148 8723 5151
rect 8754 5148 8760 5160
rect 8711 5120 8760 5148
rect 8711 5117 8723 5120
rect 8665 5111 8723 5117
rect 8389 5083 8447 5089
rect 8389 5080 8401 5083
rect 7024 5052 8401 5080
rect 6549 5043 6607 5049
rect 8389 5049 8401 5052
rect 8435 5049 8447 5083
rect 8588 5080 8616 5111
rect 8754 5108 8760 5120
rect 8812 5108 8818 5160
rect 8846 5108 8852 5160
rect 8904 5108 8910 5160
rect 8941 5151 8999 5157
rect 8941 5117 8953 5151
rect 8987 5148 8999 5151
rect 9140 5148 9168 5176
rect 8987 5120 9168 5148
rect 9217 5151 9275 5157
rect 8987 5117 8999 5120
rect 8941 5111 8999 5117
rect 9217 5117 9229 5151
rect 9263 5117 9275 5151
rect 9217 5111 9275 5117
rect 9030 5080 9036 5092
rect 8588 5052 9036 5080
rect 8389 5043 8447 5049
rect 9030 5040 9036 5052
rect 9088 5080 9094 5092
rect 9232 5080 9260 5111
rect 9306 5108 9312 5160
rect 9364 5108 9370 5160
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 9600 5157 9628 5188
rect 9493 5151 9551 5157
rect 9493 5148 9505 5151
rect 9456 5120 9505 5148
rect 9456 5108 9462 5120
rect 9493 5117 9505 5120
rect 9539 5117 9551 5151
rect 9493 5111 9551 5117
rect 9585 5151 9643 5157
rect 9585 5117 9597 5151
rect 9631 5117 9643 5151
rect 9692 5148 9720 5256
rect 10870 5244 10876 5256
rect 10928 5244 10934 5296
rect 11146 5244 11152 5296
rect 11204 5284 11210 5296
rect 12529 5287 12587 5293
rect 12529 5284 12541 5287
rect 11204 5256 12541 5284
rect 11204 5244 11210 5256
rect 12529 5253 12541 5256
rect 12575 5253 12587 5287
rect 12529 5247 12587 5253
rect 15378 5244 15384 5296
rect 15436 5244 15442 5296
rect 15562 5244 15568 5296
rect 15620 5284 15626 5296
rect 15620 5256 15700 5284
rect 15620 5244 15626 5256
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 12345 5219 12403 5225
rect 12345 5216 12357 5219
rect 10652 5188 12357 5216
rect 10652 5176 10658 5188
rect 12345 5185 12357 5188
rect 12391 5216 12403 5219
rect 13078 5216 13084 5228
rect 12391 5188 13084 5216
rect 12391 5185 12403 5188
rect 12345 5179 12403 5185
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 14185 5219 14243 5225
rect 14185 5185 14197 5219
rect 14231 5216 14243 5219
rect 14642 5216 14648 5228
rect 14231 5188 14648 5216
rect 14231 5185 14243 5188
rect 14185 5179 14243 5185
rect 14642 5176 14648 5188
rect 14700 5216 14706 5228
rect 14921 5219 14979 5225
rect 14921 5216 14933 5219
rect 14700 5188 14933 5216
rect 14700 5176 14706 5188
rect 14921 5185 14933 5188
rect 14967 5185 14979 5219
rect 15396 5216 15424 5244
rect 15672 5216 15700 5256
rect 15396 5188 15608 5216
rect 14921 5179 14979 5185
rect 9692 5120 10732 5148
rect 9585 5111 9643 5117
rect 9674 5080 9680 5092
rect 9088 5052 9680 5080
rect 9088 5040 9094 5052
rect 9674 5040 9680 5052
rect 9732 5040 9738 5092
rect 10704 5080 10732 5120
rect 11422 5108 11428 5160
rect 11480 5108 11486 5160
rect 11514 5108 11520 5160
rect 11572 5148 11578 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11572 5120 12081 5148
rect 11572 5108 11578 5120
rect 12069 5117 12081 5120
rect 12115 5148 12127 5151
rect 12158 5148 12164 5160
rect 12115 5120 12164 5148
rect 12115 5117 12127 5120
rect 12069 5111 12127 5117
rect 12158 5108 12164 5120
rect 12216 5108 12222 5160
rect 12802 5108 12808 5160
rect 12860 5148 12866 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12860 5120 12909 5148
rect 12860 5108 12866 5120
rect 12897 5117 12909 5120
rect 12943 5148 12955 5151
rect 15378 5148 15384 5160
rect 12943 5120 15384 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 15378 5108 15384 5120
rect 15436 5108 15442 5160
rect 15470 5108 15476 5160
rect 15528 5108 15534 5160
rect 14737 5083 14795 5089
rect 14737 5080 14749 5083
rect 10704 5052 14749 5080
rect 14737 5049 14749 5052
rect 14783 5049 14795 5083
rect 14737 5043 14795 5049
rect 14826 5040 14832 5092
rect 14884 5040 14890 5092
rect 15488 5080 15516 5108
rect 14936 5052 15516 5080
rect 15580 5080 15608 5188
rect 15672 5188 16252 5216
rect 15672 5157 15700 5188
rect 15657 5151 15715 5157
rect 15657 5117 15669 5151
rect 15703 5117 15715 5151
rect 15657 5111 15715 5117
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5148 15899 5151
rect 15930 5148 15936 5160
rect 15887 5120 15936 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 15930 5108 15936 5120
rect 15988 5108 15994 5160
rect 16114 5108 16120 5160
rect 16172 5108 16178 5160
rect 16224 5148 16252 5188
rect 16408 5157 16436 5324
rect 19889 5321 19901 5355
rect 19935 5352 19947 5355
rect 20254 5352 20260 5364
rect 19935 5324 20260 5352
rect 19935 5321 19947 5324
rect 19889 5315 19947 5321
rect 20254 5312 20260 5324
rect 20312 5312 20318 5364
rect 22462 5352 22468 5364
rect 20364 5324 22468 5352
rect 16669 5287 16727 5293
rect 16669 5253 16681 5287
rect 16715 5253 16727 5287
rect 16669 5247 16727 5253
rect 16684 5216 16712 5247
rect 16850 5244 16856 5296
rect 16908 5284 16914 5296
rect 16908 5256 17264 5284
rect 16908 5244 16914 5256
rect 17236 5225 17264 5256
rect 18782 5244 18788 5296
rect 18840 5284 18846 5296
rect 20364 5284 20392 5324
rect 22462 5312 22468 5324
rect 22520 5312 22526 5364
rect 22741 5355 22799 5361
rect 22741 5321 22753 5355
rect 22787 5352 22799 5355
rect 23477 5355 23535 5361
rect 23477 5352 23489 5355
rect 22787 5324 23489 5352
rect 22787 5321 22799 5324
rect 22741 5315 22799 5321
rect 23477 5321 23489 5324
rect 23523 5321 23535 5355
rect 23477 5315 23535 5321
rect 24397 5355 24455 5361
rect 24397 5321 24409 5355
rect 24443 5352 24455 5355
rect 24946 5352 24952 5364
rect 24443 5324 24952 5352
rect 24443 5321 24455 5324
rect 24397 5315 24455 5321
rect 24946 5312 24952 5324
rect 25004 5312 25010 5364
rect 25682 5312 25688 5364
rect 25740 5352 25746 5364
rect 25777 5355 25835 5361
rect 25777 5352 25789 5355
rect 25740 5324 25789 5352
rect 25740 5312 25746 5324
rect 25777 5321 25789 5324
rect 25823 5321 25835 5355
rect 25777 5315 25835 5321
rect 18840 5256 20392 5284
rect 23124 5256 24072 5284
rect 18840 5244 18846 5256
rect 17221 5219 17279 5225
rect 16684 5188 16988 5216
rect 16301 5151 16359 5157
rect 16301 5148 16313 5151
rect 16224 5120 16313 5148
rect 16301 5117 16313 5120
rect 16347 5117 16359 5151
rect 16301 5111 16359 5117
rect 16389 5151 16447 5157
rect 16389 5117 16401 5151
rect 16435 5117 16447 5151
rect 16389 5111 16447 5117
rect 16485 5151 16543 5157
rect 16485 5117 16497 5151
rect 16531 5117 16543 5151
rect 16485 5111 16543 5117
rect 15749 5083 15807 5089
rect 15749 5080 15761 5083
rect 15580 5052 15761 5080
rect 5629 5015 5687 5021
rect 5629 4981 5641 5015
rect 5675 5012 5687 5015
rect 5902 5012 5908 5024
rect 5675 4984 5908 5012
rect 5675 4981 5687 4984
rect 5629 4975 5687 4981
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7929 5015 7987 5021
rect 7929 5012 7941 5015
rect 6972 4984 7941 5012
rect 6972 4972 6978 4984
rect 7929 4981 7941 4984
rect 7975 5012 7987 5015
rect 8202 5012 8208 5024
rect 7975 4984 8208 5012
rect 7975 4981 7987 4984
rect 7929 4975 7987 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 9398 4972 9404 5024
rect 9456 5012 9462 5024
rect 10318 5012 10324 5024
rect 9456 4984 10324 5012
rect 9456 4972 9462 4984
rect 10318 4972 10324 4984
rect 10376 4972 10382 5024
rect 12161 5015 12219 5021
rect 12161 4981 12173 5015
rect 12207 5012 12219 5015
rect 12618 5012 12624 5024
rect 12207 4984 12624 5012
rect 12207 4981 12219 4984
rect 12161 4975 12219 4981
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 12986 4972 12992 5024
rect 13044 4972 13050 5024
rect 13078 4972 13084 5024
rect 13136 5012 13142 5024
rect 13909 5015 13967 5021
rect 13909 5012 13921 5015
rect 13136 4984 13921 5012
rect 13136 4972 13142 4984
rect 13909 4981 13921 4984
rect 13955 4981 13967 5015
rect 13909 4975 13967 4981
rect 14001 5015 14059 5021
rect 14001 4981 14013 5015
rect 14047 5012 14059 5015
rect 14936 5012 14964 5052
rect 15749 5049 15761 5052
rect 15795 5049 15807 5083
rect 15948 5080 15976 5108
rect 16500 5080 16528 5111
rect 16850 5108 16856 5160
rect 16908 5108 16914 5160
rect 16960 5157 16988 5188
rect 17221 5185 17233 5219
rect 17267 5185 17279 5219
rect 17221 5179 17279 5185
rect 19337 5219 19395 5225
rect 19337 5185 19349 5219
rect 19383 5216 19395 5219
rect 19426 5216 19432 5228
rect 19383 5188 19432 5216
rect 19383 5185 19395 5188
rect 19337 5179 19395 5185
rect 19426 5176 19432 5188
rect 19484 5176 19490 5228
rect 21269 5219 21327 5225
rect 21269 5185 21281 5219
rect 21315 5216 21327 5219
rect 22646 5216 22652 5228
rect 21315 5188 22652 5216
rect 21315 5185 21327 5188
rect 21269 5179 21327 5185
rect 22646 5176 22652 5188
rect 22704 5176 22710 5228
rect 16945 5151 17003 5157
rect 16945 5117 16957 5151
rect 16991 5117 17003 5151
rect 16945 5111 17003 5117
rect 17405 5151 17463 5157
rect 17405 5117 17417 5151
rect 17451 5117 17463 5151
rect 17405 5111 17463 5117
rect 17589 5151 17647 5157
rect 17589 5117 17601 5151
rect 17635 5148 17647 5151
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 17635 5120 18061 5148
rect 17635 5117 17647 5120
rect 17589 5111 17647 5117
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 17420 5080 17448 5111
rect 18782 5108 18788 5160
rect 18840 5108 18846 5160
rect 18874 5108 18880 5160
rect 18932 5108 18938 5160
rect 19245 5151 19303 5157
rect 19245 5117 19257 5151
rect 19291 5148 19303 5151
rect 20622 5148 20628 5160
rect 19291 5120 20628 5148
rect 19291 5117 19303 5120
rect 19245 5111 19303 5117
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 20990 5108 20996 5160
rect 21048 5157 21054 5160
rect 21048 5148 21060 5157
rect 21048 5120 21093 5148
rect 21048 5111 21060 5120
rect 21048 5108 21054 5111
rect 22370 5108 22376 5160
rect 22428 5108 22434 5160
rect 23014 5108 23020 5160
rect 23072 5108 23078 5160
rect 15948 5052 16528 5080
rect 17052 5052 17448 5080
rect 15749 5043 15807 5049
rect 14047 4984 14964 5012
rect 16025 5015 16083 5021
rect 14047 4981 14059 4984
rect 14001 4975 14059 4981
rect 16025 4981 16037 5015
rect 16071 5012 16083 5015
rect 17052 5012 17080 5052
rect 18598 5040 18604 5092
rect 18656 5080 18662 5092
rect 19061 5083 19119 5089
rect 19061 5080 19073 5083
rect 18656 5052 19073 5080
rect 18656 5040 18662 5052
rect 19061 5049 19073 5052
rect 19107 5049 19119 5083
rect 19061 5043 19119 5049
rect 19153 5083 19211 5089
rect 19153 5049 19165 5083
rect 19199 5080 19211 5083
rect 19334 5080 19340 5092
rect 19199 5052 19340 5080
rect 19199 5049 19211 5052
rect 19153 5043 19211 5049
rect 19334 5040 19340 5052
rect 19392 5040 19398 5092
rect 16071 4984 17080 5012
rect 16071 4981 16083 4984
rect 16025 4975 16083 4981
rect 17126 4972 17132 5024
rect 17184 4972 17190 5024
rect 18230 4972 18236 5024
rect 18288 4972 18294 5024
rect 22388 5012 22416 5108
rect 22557 5083 22615 5089
rect 22557 5049 22569 5083
rect 22603 5080 22615 5083
rect 23124 5080 23152 5256
rect 23382 5176 23388 5228
rect 23440 5216 23446 5228
rect 24044 5216 24072 5256
rect 25222 5216 25228 5228
rect 23440 5188 23888 5216
rect 23440 5176 23446 5188
rect 23201 5151 23259 5157
rect 23201 5117 23213 5151
rect 23247 5148 23259 5151
rect 23658 5148 23664 5160
rect 23247 5120 23664 5148
rect 23247 5117 23259 5120
rect 23201 5111 23259 5117
rect 23658 5108 23664 5120
rect 23716 5108 23722 5160
rect 23860 5157 23888 5188
rect 24044 5188 25228 5216
rect 24044 5160 24072 5188
rect 25222 5176 25228 5188
rect 25280 5176 25286 5228
rect 23845 5151 23903 5157
rect 23845 5117 23857 5151
rect 23891 5117 23903 5151
rect 23845 5111 23903 5117
rect 24026 5108 24032 5160
rect 24084 5108 24090 5160
rect 24302 5108 24308 5160
rect 24360 5108 24366 5160
rect 24486 5108 24492 5160
rect 24544 5108 24550 5160
rect 24581 5151 24639 5157
rect 24581 5117 24593 5151
rect 24627 5148 24639 5151
rect 25133 5151 25191 5157
rect 25133 5148 25145 5151
rect 24627 5120 25145 5148
rect 24627 5117 24639 5120
rect 24581 5111 24639 5117
rect 25133 5117 25145 5120
rect 25179 5117 25191 5151
rect 25133 5111 25191 5117
rect 22603 5052 23152 5080
rect 22603 5049 22615 5052
rect 22557 5043 22615 5049
rect 23290 5040 23296 5092
rect 23348 5040 23354 5092
rect 23509 5083 23567 5089
rect 23509 5049 23521 5083
rect 23555 5080 23567 5083
rect 23937 5083 23995 5089
rect 23937 5080 23949 5083
rect 23555 5052 23949 5080
rect 23555 5049 23567 5052
rect 23509 5043 23567 5049
rect 23937 5049 23949 5052
rect 23983 5080 23995 5083
rect 24121 5083 24179 5089
rect 24121 5080 24133 5083
rect 23983 5052 24133 5080
rect 23983 5049 23995 5052
rect 23937 5043 23995 5049
rect 24121 5049 24133 5052
rect 24167 5049 24179 5083
rect 24121 5043 24179 5049
rect 22833 5015 22891 5021
rect 22833 5012 22845 5015
rect 22388 4984 22845 5012
rect 22833 4981 22845 4984
rect 22879 5012 22891 5015
rect 23382 5012 23388 5024
rect 22879 4984 23388 5012
rect 22879 4981 22891 4984
rect 22833 4975 22891 4981
rect 23382 4972 23388 4984
rect 23440 4972 23446 5024
rect 23658 4972 23664 5024
rect 23716 4972 23722 5024
rect 552 4922 27576 4944
rect 552 4870 7114 4922
rect 7166 4870 7178 4922
rect 7230 4870 7242 4922
rect 7294 4870 7306 4922
rect 7358 4870 7370 4922
rect 7422 4870 13830 4922
rect 13882 4870 13894 4922
rect 13946 4870 13958 4922
rect 14010 4870 14022 4922
rect 14074 4870 14086 4922
rect 14138 4870 20546 4922
rect 20598 4870 20610 4922
rect 20662 4870 20674 4922
rect 20726 4870 20738 4922
rect 20790 4870 20802 4922
rect 20854 4870 27262 4922
rect 27314 4870 27326 4922
rect 27378 4870 27390 4922
rect 27442 4870 27454 4922
rect 27506 4870 27518 4922
rect 27570 4870 27576 4922
rect 552 4848 27576 4870
rect 6914 4808 6920 4820
rect 5092 4780 6920 4808
rect 5092 4740 5120 4780
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 8294 4808 8300 4820
rect 7760 4780 8300 4808
rect 5813 4743 5871 4749
rect 5813 4740 5825 4743
rect 3804 4712 5120 4740
rect 3804 4681 3832 4712
rect 3697 4675 3755 4681
rect 3697 4641 3709 4675
rect 3743 4641 3755 4675
rect 3697 4635 3755 4641
rect 3789 4675 3847 4681
rect 3789 4641 3801 4675
rect 3835 4641 3847 4675
rect 3789 4635 3847 4641
rect 3881 4675 3939 4681
rect 3881 4641 3893 4675
rect 3927 4672 3939 4675
rect 3927 4644 4016 4672
rect 3927 4641 3939 4644
rect 3881 4635 3939 4641
rect 3712 4604 3740 4635
rect 3712 4576 3832 4604
rect 3418 4428 3424 4480
rect 3476 4428 3482 4480
rect 3804 4468 3832 4576
rect 3988 4536 4016 4644
rect 4062 4632 4068 4684
rect 4120 4632 4126 4684
rect 4798 4564 4804 4616
rect 4856 4564 4862 4616
rect 5092 4604 5120 4712
rect 5184 4712 5825 4740
rect 5184 4681 5212 4712
rect 5813 4709 5825 4712
rect 5859 4709 5871 4743
rect 5813 4703 5871 4709
rect 5902 4700 5908 4752
rect 5960 4740 5966 4752
rect 6825 4743 6883 4749
rect 6825 4740 6837 4743
rect 5960 4712 6837 4740
rect 5960 4700 5966 4712
rect 6825 4709 6837 4712
rect 6871 4709 6883 4743
rect 7650 4740 7656 4752
rect 6825 4703 6883 4709
rect 7116 4712 7656 4740
rect 7116 4684 7144 4712
rect 7650 4700 7656 4712
rect 7708 4700 7714 4752
rect 5169 4675 5227 4681
rect 5169 4641 5181 4675
rect 5215 4641 5227 4675
rect 5169 4635 5227 4641
rect 5261 4675 5319 4681
rect 5261 4641 5273 4675
rect 5307 4641 5319 4675
rect 5261 4635 5319 4641
rect 5276 4604 5304 4635
rect 5350 4632 5356 4684
rect 5408 4632 5414 4684
rect 5537 4675 5595 4681
rect 5537 4641 5549 4675
rect 5583 4672 5595 4675
rect 5626 4672 5632 4684
rect 5583 4644 5632 4672
rect 5583 4641 5595 4644
rect 5537 4635 5595 4641
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 6733 4675 6791 4681
rect 6733 4672 6745 4675
rect 5736 4644 6745 4672
rect 5092 4576 5304 4604
rect 5442 4564 5448 4616
rect 5500 4604 5506 4616
rect 5736 4604 5764 4644
rect 6733 4641 6745 4644
rect 6779 4641 6791 4675
rect 6733 4635 6791 4641
rect 6914 4632 6920 4684
rect 6972 4632 6978 4684
rect 7098 4632 7104 4684
rect 7156 4632 7162 4684
rect 7469 4675 7527 4681
rect 7469 4641 7481 4675
rect 7515 4641 7527 4675
rect 7469 4635 7527 4641
rect 5500 4576 5764 4604
rect 5500 4564 5506 4576
rect 6362 4564 6368 4616
rect 6420 4564 6426 4616
rect 7484 4604 7512 4635
rect 7558 4632 7564 4684
rect 7616 4632 7622 4684
rect 7760 4681 7788 4780
rect 8294 4768 8300 4780
rect 8352 4808 8358 4820
rect 8754 4808 8760 4820
rect 8352 4780 8760 4808
rect 8352 4768 8358 4780
rect 8018 4700 8024 4752
rect 8076 4740 8082 4752
rect 8076 4712 8524 4740
rect 8076 4700 8082 4712
rect 7745 4675 7803 4681
rect 7745 4641 7757 4675
rect 7791 4641 7803 4675
rect 7745 4635 7803 4641
rect 7837 4675 7895 4681
rect 7837 4641 7849 4675
rect 7883 4672 7895 4675
rect 8036 4672 8064 4700
rect 7883 4644 8064 4672
rect 8113 4675 8171 4681
rect 7883 4641 7895 4644
rect 7837 4635 7895 4641
rect 8113 4641 8125 4675
rect 8159 4641 8171 4675
rect 8113 4635 8171 4641
rect 8128 4604 8156 4635
rect 8202 4632 8208 4684
rect 8260 4632 8266 4684
rect 8294 4632 8300 4684
rect 8352 4672 8358 4684
rect 8496 4681 8524 4712
rect 8389 4675 8447 4681
rect 8389 4672 8401 4675
rect 8352 4644 8401 4672
rect 8352 4632 8358 4644
rect 8389 4641 8401 4644
rect 8435 4641 8447 4675
rect 8389 4635 8447 4641
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4672 8539 4675
rect 8570 4672 8576 4684
rect 8527 4644 8576 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 8680 4681 8708 4780
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 9214 4808 9220 4820
rect 8864 4780 9220 4808
rect 8864 4681 8892 4780
rect 9214 4768 9220 4780
rect 9272 4768 9278 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 10134 4808 10140 4820
rect 9640 4780 10140 4808
rect 9640 4768 9646 4780
rect 10134 4768 10140 4780
rect 10192 4808 10198 4820
rect 10778 4808 10784 4820
rect 10192 4780 10784 4808
rect 10192 4768 10198 4780
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 11514 4808 11520 4820
rect 10980 4780 11520 4808
rect 10980 4740 11008 4780
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 11606 4768 11612 4820
rect 11664 4768 11670 4820
rect 12434 4808 12440 4820
rect 12406 4768 12440 4808
rect 12492 4768 12498 4820
rect 15286 4768 15292 4820
rect 15344 4768 15350 4820
rect 15470 4768 15476 4820
rect 15528 4808 15534 4820
rect 19794 4808 19800 4820
rect 15528 4780 19800 4808
rect 15528 4768 15534 4780
rect 19794 4768 19800 4780
rect 19852 4768 19858 4820
rect 23937 4811 23995 4817
rect 23937 4777 23949 4811
rect 23983 4808 23995 4811
rect 24026 4808 24032 4820
rect 23983 4780 24032 4808
rect 23983 4777 23995 4780
rect 23937 4771 23995 4777
rect 24026 4768 24032 4780
rect 24084 4768 24090 4820
rect 12406 4740 12434 4768
rect 10520 4712 11008 4740
rect 11348 4712 12434 4740
rect 8665 4675 8723 4681
rect 8665 4641 8677 4675
rect 8711 4641 8723 4675
rect 8665 4635 8723 4641
rect 8849 4675 8907 4681
rect 8849 4641 8861 4675
rect 8895 4641 8907 4675
rect 8849 4635 8907 4641
rect 8941 4675 8999 4681
rect 8941 4641 8953 4675
rect 8987 4672 8999 4675
rect 9030 4672 9036 4684
rect 8987 4644 9036 4672
rect 8987 4641 8999 4644
rect 8941 4635 8999 4641
rect 8956 4604 8984 4635
rect 9030 4632 9036 4644
rect 9088 4632 9094 4684
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 9217 4675 9275 4681
rect 9217 4672 9229 4675
rect 9180 4644 9229 4672
rect 9180 4632 9186 4644
rect 9217 4641 9229 4644
rect 9263 4641 9275 4675
rect 9217 4635 9275 4641
rect 9306 4632 9312 4684
rect 9364 4632 9370 4684
rect 9447 4675 9505 4681
rect 9447 4641 9459 4675
rect 9493 4641 9505 4675
rect 9447 4635 9505 4641
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4641 9643 4675
rect 9585 4635 9643 4641
rect 7484 4576 8984 4604
rect 7285 4539 7343 4545
rect 7285 4536 7297 4539
rect 3988 4508 7297 4536
rect 7285 4505 7297 4508
rect 7331 4505 7343 4539
rect 7285 4499 7343 4505
rect 8570 4496 8576 4548
rect 8628 4536 8634 4548
rect 9140 4536 9168 4632
rect 8628 4508 9168 4536
rect 9468 4508 9496 4635
rect 9600 4604 9628 4635
rect 10226 4632 10232 4684
rect 10284 4632 10290 4684
rect 10318 4632 10324 4684
rect 10376 4632 10382 4684
rect 10520 4681 10548 4712
rect 10505 4675 10563 4681
rect 10505 4641 10517 4675
rect 10551 4641 10563 4675
rect 10505 4635 10563 4641
rect 10594 4632 10600 4684
rect 10652 4632 10658 4684
rect 10870 4632 10876 4684
rect 10928 4672 10934 4684
rect 10965 4675 11023 4681
rect 10965 4672 10977 4675
rect 10928 4644 10977 4672
rect 10928 4632 10934 4644
rect 10965 4641 10977 4644
rect 11011 4641 11023 4675
rect 10965 4635 11023 4641
rect 11054 4632 11060 4684
rect 11112 4672 11118 4684
rect 11149 4675 11207 4681
rect 11149 4672 11161 4675
rect 11112 4644 11161 4672
rect 11112 4632 11118 4644
rect 11149 4641 11161 4644
rect 11195 4641 11207 4675
rect 11149 4635 11207 4641
rect 11238 4632 11244 4684
rect 11296 4632 11302 4684
rect 11348 4681 11376 4712
rect 14642 4700 14648 4752
rect 14700 4740 14706 4752
rect 16666 4740 16672 4752
rect 14700 4712 16672 4740
rect 14700 4700 14706 4712
rect 16666 4700 16672 4712
rect 16724 4740 16730 4752
rect 17310 4740 17316 4752
rect 16724 4712 17316 4740
rect 16724 4700 16730 4712
rect 17310 4700 17316 4712
rect 17368 4700 17374 4752
rect 17954 4740 17960 4752
rect 17420 4712 17960 4740
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4641 11391 4675
rect 11333 4635 11391 4641
rect 12161 4675 12219 4681
rect 12161 4641 12173 4675
rect 12207 4641 12219 4675
rect 12161 4635 12219 4641
rect 9674 4604 9680 4616
rect 9600 4576 9680 4604
rect 9674 4564 9680 4576
rect 9732 4604 9738 4616
rect 10612 4604 10640 4632
rect 9732 4576 10640 4604
rect 12176 4604 12204 4635
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 12308 4644 12357 4672
rect 12308 4632 12314 4644
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 12434 4632 12440 4684
rect 12492 4632 12498 4684
rect 12529 4675 12587 4681
rect 12529 4641 12541 4675
rect 12575 4672 12587 4675
rect 12802 4672 12808 4684
rect 12575 4644 12808 4672
rect 12575 4641 12587 4644
rect 12529 4635 12587 4641
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 15105 4675 15163 4681
rect 15105 4641 15117 4675
rect 15151 4672 15163 4675
rect 15194 4672 15200 4684
rect 15151 4644 15200 4672
rect 15151 4641 15163 4644
rect 15105 4635 15163 4641
rect 15194 4632 15200 4644
rect 15252 4672 15258 4684
rect 15562 4672 15568 4684
rect 15252 4644 15568 4672
rect 15252 4632 15258 4644
rect 15562 4632 15568 4644
rect 15620 4672 15626 4684
rect 15838 4672 15844 4684
rect 15620 4644 15844 4672
rect 15620 4632 15626 4644
rect 15838 4632 15844 4644
rect 15896 4632 15902 4684
rect 17126 4632 17132 4684
rect 17184 4632 17190 4684
rect 17420 4681 17448 4712
rect 17954 4700 17960 4712
rect 18012 4700 18018 4752
rect 18230 4700 18236 4752
rect 18288 4740 18294 4752
rect 19122 4743 19180 4749
rect 19122 4740 19134 4743
rect 18288 4712 19134 4740
rect 18288 4700 18294 4712
rect 19122 4709 19134 4712
rect 19168 4709 19180 4743
rect 19122 4703 19180 4709
rect 22462 4700 22468 4752
rect 22520 4740 22526 4752
rect 24486 4740 24492 4752
rect 22520 4712 24492 4740
rect 22520 4700 22526 4712
rect 24486 4700 24492 4712
rect 24544 4700 24550 4752
rect 17405 4675 17463 4681
rect 17405 4641 17417 4675
rect 17451 4641 17463 4675
rect 17661 4675 17719 4681
rect 17661 4672 17673 4675
rect 17405 4635 17463 4641
rect 17512 4644 17673 4672
rect 13078 4604 13084 4616
rect 12176 4576 13084 4604
rect 9732 4564 9738 4576
rect 13078 4564 13084 4576
rect 13136 4564 13142 4616
rect 14918 4564 14924 4616
rect 14976 4604 14982 4616
rect 16390 4604 16396 4616
rect 14976 4576 16396 4604
rect 14976 4564 14982 4576
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 17512 4604 17540 4644
rect 17661 4641 17673 4644
rect 17707 4641 17719 4675
rect 17972 4672 18000 4700
rect 18877 4675 18935 4681
rect 18877 4672 18889 4675
rect 17972 4644 18889 4672
rect 17661 4635 17719 4641
rect 18877 4641 18889 4644
rect 18923 4672 18935 4675
rect 18966 4672 18972 4684
rect 18923 4644 18972 4672
rect 18923 4641 18935 4644
rect 18877 4635 18935 4641
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 22557 4675 22615 4681
rect 22557 4641 22569 4675
rect 22603 4672 22615 4675
rect 22646 4672 22652 4684
rect 22603 4644 22652 4672
rect 22603 4641 22615 4644
rect 22557 4635 22615 4641
rect 22646 4632 22652 4644
rect 22704 4632 22710 4684
rect 22830 4681 22836 4684
rect 22824 4635 22836 4681
rect 22830 4632 22836 4635
rect 22888 4632 22894 4684
rect 17328 4576 17540 4604
rect 8628 4496 8634 4508
rect 9490 4496 9496 4508
rect 9548 4496 9554 4548
rect 15286 4536 15292 4548
rect 12636 4508 15292 4536
rect 4157 4471 4215 4477
rect 4157 4468 4169 4471
rect 3804 4440 4169 4468
rect 4157 4437 4169 4440
rect 4203 4437 4215 4471
rect 4157 4431 4215 4437
rect 4890 4428 4896 4480
rect 4948 4428 4954 4480
rect 4982 4428 4988 4480
rect 5040 4468 5046 4480
rect 6549 4471 6607 4477
rect 6549 4468 6561 4471
rect 5040 4440 6561 4468
rect 5040 4428 5046 4440
rect 6549 4437 6561 4440
rect 6595 4437 6607 4471
rect 6549 4431 6607 4437
rect 7374 4428 7380 4480
rect 7432 4468 7438 4480
rect 7929 4471 7987 4477
rect 7929 4468 7941 4471
rect 7432 4440 7941 4468
rect 7432 4428 7438 4440
rect 7929 4437 7941 4440
rect 7975 4437 7987 4471
rect 7929 4431 7987 4437
rect 9030 4428 9036 4480
rect 9088 4468 9094 4480
rect 9125 4471 9183 4477
rect 9125 4468 9137 4471
rect 9088 4440 9137 4468
rect 9088 4428 9094 4440
rect 9125 4437 9137 4440
rect 9171 4437 9183 4471
rect 9125 4431 9183 4437
rect 9766 4428 9772 4480
rect 9824 4428 9830 4480
rect 10781 4471 10839 4477
rect 10781 4437 10793 4471
rect 10827 4468 10839 4471
rect 11146 4468 11152 4480
rect 10827 4440 11152 4468
rect 10827 4437 10839 4440
rect 10781 4431 10839 4437
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 12250 4428 12256 4480
rect 12308 4468 12314 4480
rect 12636 4468 12664 4508
rect 15286 4496 15292 4508
rect 15344 4496 15350 4548
rect 17328 4545 17356 4576
rect 17313 4539 17371 4545
rect 17313 4505 17325 4539
rect 17359 4505 17371 4539
rect 17313 4499 17371 4505
rect 12308 4440 12664 4468
rect 12308 4428 12314 4440
rect 12710 4428 12716 4480
rect 12768 4428 12774 4480
rect 14826 4428 14832 4480
rect 14884 4468 14890 4480
rect 16114 4468 16120 4480
rect 14884 4440 16120 4468
rect 14884 4428 14890 4440
rect 16114 4428 16120 4440
rect 16172 4468 16178 4480
rect 18785 4471 18843 4477
rect 18785 4468 18797 4471
rect 16172 4440 18797 4468
rect 16172 4428 16178 4440
rect 18785 4437 18797 4440
rect 18831 4468 18843 4471
rect 19242 4468 19248 4480
rect 18831 4440 19248 4468
rect 18831 4437 18843 4440
rect 18785 4431 18843 4437
rect 19242 4428 19248 4440
rect 19300 4428 19306 4480
rect 19794 4428 19800 4480
rect 19852 4468 19858 4480
rect 20257 4471 20315 4477
rect 20257 4468 20269 4471
rect 19852 4440 20269 4468
rect 19852 4428 19858 4440
rect 20257 4437 20269 4440
rect 20303 4437 20315 4471
rect 20257 4431 20315 4437
rect 552 4378 27416 4400
rect 552 4326 3756 4378
rect 3808 4326 3820 4378
rect 3872 4326 3884 4378
rect 3936 4326 3948 4378
rect 4000 4326 4012 4378
rect 4064 4326 10472 4378
rect 10524 4326 10536 4378
rect 10588 4326 10600 4378
rect 10652 4326 10664 4378
rect 10716 4326 10728 4378
rect 10780 4326 17188 4378
rect 17240 4326 17252 4378
rect 17304 4326 17316 4378
rect 17368 4326 17380 4378
rect 17432 4326 17444 4378
rect 17496 4326 23904 4378
rect 23956 4326 23968 4378
rect 24020 4326 24032 4378
rect 24084 4326 24096 4378
rect 24148 4326 24160 4378
rect 24212 4326 27416 4378
rect 552 4304 27416 4326
rect 5445 4267 5503 4273
rect 5445 4233 5457 4267
rect 5491 4264 5503 4267
rect 5626 4264 5632 4276
rect 5491 4236 5632 4264
rect 5491 4233 5503 4236
rect 5445 4227 5503 4233
rect 5626 4224 5632 4236
rect 5684 4264 5690 4276
rect 6362 4264 6368 4276
rect 5684 4236 6368 4264
rect 5684 4224 5690 4236
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 12618 4224 12624 4276
rect 12676 4224 12682 4276
rect 12986 4224 12992 4276
rect 13044 4264 13050 4276
rect 13541 4267 13599 4273
rect 13541 4264 13553 4267
rect 13044 4236 13553 4264
rect 13044 4224 13050 4236
rect 13541 4233 13553 4236
rect 13587 4233 13599 4267
rect 13541 4227 13599 4233
rect 14826 4224 14832 4276
rect 14884 4264 14890 4276
rect 15286 4264 15292 4276
rect 14884 4236 15292 4264
rect 14884 4224 14890 4236
rect 15286 4224 15292 4236
rect 15344 4224 15350 4276
rect 15930 4264 15936 4276
rect 15580 4236 15936 4264
rect 7098 4196 7104 4208
rect 6932 4168 7104 4196
rect 6178 4088 6184 4140
rect 6236 4128 6242 4140
rect 6932 4128 6960 4168
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 9950 4196 9956 4208
rect 9692 4168 9956 4196
rect 6236 4100 6960 4128
rect 6236 4088 6242 4100
rect 7006 4088 7012 4140
rect 7064 4128 7070 4140
rect 7064 4100 8984 4128
rect 7064 4088 7070 4100
rect 3789 4063 3847 4069
rect 3789 4029 3801 4063
rect 3835 4029 3847 4063
rect 3789 4023 3847 4029
rect 3605 3927 3663 3933
rect 3605 3893 3617 3927
rect 3651 3924 3663 3927
rect 3694 3924 3700 3936
rect 3651 3896 3700 3924
rect 3651 3893 3663 3896
rect 3605 3887 3663 3893
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 3804 3924 3832 4023
rect 3970 4020 3976 4072
rect 4028 4020 4034 4072
rect 4065 4063 4123 4069
rect 4065 4029 4077 4063
rect 4111 4060 4123 4063
rect 5534 4060 5540 4072
rect 4111 4032 5540 4060
rect 4111 4029 4123 4032
rect 4065 4023 4123 4029
rect 3878 3952 3884 4004
rect 3936 3992 3942 4004
rect 4080 3992 4108 4023
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 7208 4069 7236 4100
rect 7101 4063 7159 4069
rect 7101 4029 7113 4063
rect 7147 4029 7159 4063
rect 7101 4023 7159 4029
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4029 7251 4063
rect 7193 4023 7251 4029
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4060 7343 4063
rect 7374 4060 7380 4072
rect 7331 4032 7380 4060
rect 7331 4029 7343 4032
rect 7285 4023 7343 4029
rect 3936 3964 4108 3992
rect 4332 3995 4390 4001
rect 3936 3952 3942 3964
rect 4332 3961 4344 3995
rect 4378 3992 4390 3995
rect 4890 3992 4896 4004
rect 4378 3964 4896 3992
rect 4378 3961 4390 3964
rect 4332 3955 4390 3961
rect 4890 3952 4896 3964
rect 4948 3952 4954 4004
rect 7116 3992 7144 4023
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 7466 4020 7472 4072
rect 7524 4020 7530 4072
rect 7834 4020 7840 4072
rect 7892 4060 7898 4072
rect 8113 4063 8171 4069
rect 8113 4060 8125 4063
rect 7892 4032 8125 4060
rect 7892 4020 7898 4032
rect 8113 4029 8125 4032
rect 8159 4029 8171 4063
rect 8113 4023 8171 4029
rect 7561 3995 7619 4001
rect 7561 3992 7573 3995
rect 7116 3964 7573 3992
rect 7561 3961 7573 3964
rect 7607 3961 7619 3995
rect 7561 3955 7619 3961
rect 4982 3924 4988 3936
rect 3804 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 6822 3884 6828 3936
rect 6880 3884 6886 3936
rect 8570 3884 8576 3936
rect 8628 3884 8634 3936
rect 8772 3924 8800 4100
rect 8956 4069 8984 4100
rect 8849 4063 8907 4069
rect 8849 4029 8861 4063
rect 8895 4029 8907 4063
rect 8849 4023 8907 4029
rect 8941 4063 8999 4069
rect 8941 4029 8953 4063
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 8864 3992 8892 4023
rect 9030 4020 9036 4072
rect 9088 4020 9094 4072
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4060 9275 4063
rect 9692 4060 9720 4168
rect 9950 4156 9956 4168
rect 10008 4196 10014 4208
rect 14642 4196 14648 4208
rect 10008 4168 10640 4196
rect 10008 4156 10014 4168
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 9824 4100 10548 4128
rect 9824 4088 9830 4100
rect 9263 4032 9720 4060
rect 9263 4029 9275 4032
rect 9217 4023 9275 4029
rect 9858 4020 9864 4072
rect 9916 4020 9922 4072
rect 10318 4020 10324 4072
rect 10376 4020 10382 4072
rect 10520 4069 10548 4100
rect 10413 4063 10471 4069
rect 10413 4029 10425 4063
rect 10459 4029 10471 4063
rect 10413 4023 10471 4029
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4029 10563 4063
rect 10612 4060 10640 4168
rect 13280 4168 14648 4196
rect 13280 4137 13308 4168
rect 14200 4137 14228 4168
rect 14642 4156 14648 4168
rect 14700 4156 14706 4208
rect 15010 4156 15016 4208
rect 15068 4196 15074 4208
rect 15580 4196 15608 4236
rect 15930 4224 15936 4236
rect 15988 4264 15994 4276
rect 16298 4264 16304 4276
rect 15988 4236 16304 4264
rect 15988 4224 15994 4236
rect 16298 4224 16304 4236
rect 16356 4224 16362 4276
rect 22094 4264 22100 4276
rect 19306 4236 22100 4264
rect 15068 4168 15608 4196
rect 15068 4156 15074 4168
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4097 13323 4131
rect 13265 4091 13323 4097
rect 14185 4131 14243 4137
rect 14185 4097 14197 4131
rect 14231 4097 14243 4131
rect 15194 4128 15200 4140
rect 14185 4091 14243 4097
rect 14844 4100 15200 4128
rect 10689 4063 10747 4069
rect 10689 4060 10701 4063
rect 10612 4032 10701 4060
rect 10505 4023 10563 4029
rect 10689 4029 10701 4032
rect 10735 4060 10747 4063
rect 10965 4063 11023 4069
rect 10965 4060 10977 4063
rect 10735 4032 10977 4060
rect 10735 4029 10747 4032
rect 10689 4023 10747 4029
rect 10965 4029 10977 4032
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 8864 3964 9321 3992
rect 9309 3961 9321 3964
rect 9355 3961 9367 3995
rect 10428 3992 10456 4023
rect 11146 4020 11152 4072
rect 11204 4020 11210 4072
rect 11238 4020 11244 4072
rect 11296 4020 11302 4072
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 11885 4063 11943 4069
rect 11885 4060 11897 4063
rect 11379 4032 11897 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11885 4029 11897 4032
rect 11931 4029 11943 4063
rect 11885 4023 11943 4029
rect 12434 4020 12440 4072
rect 12492 4020 12498 4072
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4060 13139 4063
rect 14642 4060 14648 4072
rect 13127 4032 14648 4060
rect 13127 4029 13139 4032
rect 13081 4023 13139 4029
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 14844 4069 14872 4100
rect 15194 4088 15200 4100
rect 15252 4128 15258 4140
rect 15252 4100 15516 4128
rect 15252 4088 15258 4100
rect 14829 4063 14887 4069
rect 14829 4029 14841 4063
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 15010 4020 15016 4072
rect 15068 4020 15074 4072
rect 15488 4069 15516 4100
rect 15289 4063 15347 4069
rect 15289 4060 15301 4063
rect 15120 4032 15301 4060
rect 11256 3992 11284 4020
rect 9309 3955 9367 3961
rect 9968 3964 11284 3992
rect 9968 3924 9996 3964
rect 12066 3952 12072 4004
rect 12124 3992 12130 4004
rect 12989 3995 13047 4001
rect 12989 3992 13001 3995
rect 12124 3964 13001 3992
rect 12124 3952 12130 3964
rect 12989 3961 13001 3964
rect 13035 3961 13047 3995
rect 12989 3955 13047 3961
rect 13909 3995 13967 4001
rect 13909 3961 13921 3995
rect 13955 3992 13967 3995
rect 14182 3992 14188 4004
rect 13955 3964 14188 3992
rect 13955 3961 13967 3964
rect 13909 3955 13967 3961
rect 14182 3952 14188 3964
rect 14240 3952 14246 4004
rect 14274 3952 14280 4004
rect 14332 3992 14338 4004
rect 14921 3995 14979 4001
rect 14921 3992 14933 3995
rect 14332 3964 14933 3992
rect 14332 3952 14338 3964
rect 14921 3961 14933 3964
rect 14967 3961 14979 3995
rect 14921 3955 14979 3961
rect 15120 3992 15148 4032
rect 15289 4029 15301 4032
rect 15335 4029 15347 4063
rect 15289 4023 15347 4029
rect 15473 4063 15531 4069
rect 15473 4029 15485 4063
rect 15519 4029 15531 4063
rect 15580 4060 15608 4168
rect 15841 4199 15899 4205
rect 15841 4165 15853 4199
rect 15887 4196 15899 4199
rect 15887 4168 17724 4196
rect 15887 4165 15899 4168
rect 15841 4159 15899 4165
rect 17696 4128 17724 4168
rect 17770 4156 17776 4208
rect 17828 4196 17834 4208
rect 19306 4196 19334 4236
rect 22094 4224 22100 4236
rect 22152 4224 22158 4276
rect 22830 4224 22836 4276
rect 22888 4224 22894 4276
rect 17828 4168 19334 4196
rect 17828 4156 17834 4168
rect 19076 4137 19104 4168
rect 19061 4131 19119 4137
rect 17696 4100 18184 4128
rect 15657 4063 15715 4069
rect 15657 4060 15669 4063
rect 15580 4032 15669 4060
rect 15473 4023 15531 4029
rect 15657 4029 15669 4032
rect 15703 4029 15715 4063
rect 15657 4023 15715 4029
rect 15930 4020 15936 4072
rect 15988 4020 15994 4072
rect 16298 4020 16304 4072
rect 16356 4060 16362 4072
rect 16574 4060 16580 4072
rect 16356 4032 16580 4060
rect 16356 4020 16362 4032
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 16850 4020 16856 4072
rect 16908 4060 16914 4072
rect 17770 4060 17776 4072
rect 16908 4032 17776 4060
rect 16908 4020 16914 4032
rect 17770 4020 17776 4032
rect 17828 4060 17834 4072
rect 18156 4069 18184 4100
rect 19061 4097 19073 4131
rect 19107 4097 19119 4131
rect 19061 4091 19119 4097
rect 19150 4088 19156 4140
rect 19208 4128 19214 4140
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 19208 4100 19441 4128
rect 19208 4088 19214 4100
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 19429 4091 19487 4097
rect 17957 4063 18015 4069
rect 17957 4060 17969 4063
rect 17828 4032 17969 4060
rect 17828 4020 17834 4032
rect 17957 4029 17969 4032
rect 18003 4029 18015 4063
rect 17957 4023 18015 4029
rect 18141 4063 18199 4069
rect 18141 4029 18153 4063
rect 18187 4029 18199 4063
rect 18141 4023 18199 4029
rect 18877 4063 18935 4069
rect 18877 4029 18889 4063
rect 18923 4029 18935 4063
rect 18877 4023 18935 4029
rect 23017 4063 23075 4069
rect 23017 4029 23029 4063
rect 23063 4060 23075 4063
rect 23658 4060 23664 4072
rect 23063 4032 23664 4060
rect 23063 4029 23075 4032
rect 23017 4023 23075 4029
rect 15120 3964 15516 3992
rect 8772 3896 9996 3924
rect 10042 3884 10048 3936
rect 10100 3884 10106 3936
rect 11606 3884 11612 3936
rect 11664 3884 11670 3936
rect 14001 3927 14059 3933
rect 14001 3893 14013 3927
rect 14047 3924 14059 3927
rect 15120 3924 15148 3964
rect 14047 3896 15148 3924
rect 14047 3893 14059 3896
rect 14001 3887 14059 3893
rect 15194 3884 15200 3936
rect 15252 3884 15258 3936
rect 15488 3924 15516 3964
rect 15562 3952 15568 4004
rect 15620 3952 15626 4004
rect 15838 3952 15844 4004
rect 15896 3992 15902 4004
rect 16117 3995 16175 4001
rect 16117 3992 16129 3995
rect 15896 3964 16129 3992
rect 15896 3952 15902 3964
rect 16117 3961 16129 3964
rect 16163 3961 16175 3995
rect 16117 3955 16175 3961
rect 16022 3924 16028 3936
rect 15488 3896 16028 3924
rect 16022 3884 16028 3896
rect 16080 3884 16086 3936
rect 16132 3924 16160 3955
rect 16206 3952 16212 4004
rect 16264 3952 16270 4004
rect 18892 3992 18920 4023
rect 23658 4020 23664 4032
rect 23716 4020 23722 4072
rect 19674 3995 19732 4001
rect 19674 3992 19686 3995
rect 16500 3964 18920 3992
rect 18984 3964 19686 3992
rect 16298 3924 16304 3936
rect 16132 3896 16304 3924
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 16500 3933 16528 3964
rect 16485 3927 16543 3933
rect 16485 3893 16497 3927
rect 16531 3893 16543 3927
rect 16485 3887 16543 3893
rect 18322 3884 18328 3936
rect 18380 3884 18386 3936
rect 18506 3884 18512 3936
rect 18564 3924 18570 3936
rect 18693 3927 18751 3933
rect 18693 3924 18705 3927
rect 18564 3896 18705 3924
rect 18564 3884 18570 3896
rect 18693 3893 18705 3896
rect 18739 3893 18751 3927
rect 18693 3887 18751 3893
rect 18782 3884 18788 3936
rect 18840 3924 18846 3936
rect 18984 3924 19012 3964
rect 19674 3961 19686 3964
rect 19720 3961 19732 3995
rect 19674 3955 19732 3961
rect 18840 3896 19012 3924
rect 20809 3927 20867 3933
rect 18840 3884 18846 3896
rect 20809 3893 20821 3927
rect 20855 3924 20867 3927
rect 21450 3924 21456 3936
rect 20855 3896 21456 3924
rect 20855 3893 20867 3896
rect 20809 3887 20867 3893
rect 21450 3884 21456 3896
rect 21508 3884 21514 3936
rect 552 3834 27576 3856
rect 552 3782 7114 3834
rect 7166 3782 7178 3834
rect 7230 3782 7242 3834
rect 7294 3782 7306 3834
rect 7358 3782 7370 3834
rect 7422 3782 13830 3834
rect 13882 3782 13894 3834
rect 13946 3782 13958 3834
rect 14010 3782 14022 3834
rect 14074 3782 14086 3834
rect 14138 3782 20546 3834
rect 20598 3782 20610 3834
rect 20662 3782 20674 3834
rect 20726 3782 20738 3834
rect 20790 3782 20802 3834
rect 20854 3782 27262 3834
rect 27314 3782 27326 3834
rect 27378 3782 27390 3834
rect 27442 3782 27454 3834
rect 27506 3782 27518 3834
rect 27570 3782 27576 3834
rect 552 3760 27576 3782
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 5169 3723 5227 3729
rect 5169 3720 5181 3723
rect 4856 3692 5181 3720
rect 4856 3680 4862 3692
rect 5169 3689 5181 3692
rect 5215 3689 5227 3723
rect 5169 3683 5227 3689
rect 7834 3680 7840 3732
rect 7892 3680 7898 3732
rect 10318 3680 10324 3732
rect 10376 3720 10382 3732
rect 10781 3723 10839 3729
rect 10781 3720 10793 3723
rect 10376 3692 10793 3720
rect 10376 3680 10382 3692
rect 10781 3689 10793 3692
rect 10827 3689 10839 3723
rect 10781 3683 10839 3689
rect 12434 3680 12440 3732
rect 12492 3680 12498 3732
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 13909 3723 13967 3729
rect 13909 3720 13921 3723
rect 13780 3692 13921 3720
rect 13780 3680 13786 3692
rect 13909 3689 13921 3692
rect 13955 3689 13967 3723
rect 13909 3683 13967 3689
rect 14366 3680 14372 3732
rect 14424 3720 14430 3732
rect 14737 3723 14795 3729
rect 14737 3720 14749 3723
rect 14424 3692 14749 3720
rect 14424 3680 14430 3692
rect 14737 3689 14749 3692
rect 14783 3689 14795 3723
rect 15930 3720 15936 3732
rect 14737 3683 14795 3689
rect 15120 3692 15936 3720
rect 3418 3612 3424 3664
rect 3476 3652 3482 3664
rect 4034 3655 4092 3661
rect 4034 3652 4046 3655
rect 3476 3624 4046 3652
rect 3476 3612 3482 3624
rect 4034 3621 4046 3624
rect 4080 3621 4092 3655
rect 4034 3615 4092 3621
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 5258 3652 5264 3664
rect 4212 3624 5264 3652
rect 4212 3612 4218 3624
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 6724 3655 6782 3661
rect 6724 3621 6736 3655
rect 6770 3652 6782 3655
rect 6822 3652 6828 3664
rect 6770 3624 6828 3652
rect 6770 3621 6782 3624
rect 6724 3615 6782 3621
rect 6822 3612 6828 3624
rect 6880 3612 6886 3664
rect 11324 3655 11382 3661
rect 8312 3624 9996 3652
rect 3694 3544 3700 3596
rect 3752 3544 3758 3596
rect 3789 3587 3847 3593
rect 3789 3553 3801 3587
rect 3835 3584 3847 3587
rect 3878 3584 3884 3596
rect 3835 3556 3884 3584
rect 3835 3553 3847 3556
rect 3789 3547 3847 3553
rect 3326 3476 3332 3528
rect 3384 3516 3390 3528
rect 3804 3516 3832 3547
rect 3878 3544 3884 3556
rect 3936 3544 3942 3596
rect 5534 3544 5540 3596
rect 5592 3584 5598 3596
rect 6362 3584 6368 3596
rect 5592 3556 6368 3584
rect 5592 3544 5598 3556
rect 6362 3544 6368 3556
rect 6420 3584 6426 3596
rect 8312 3593 8340 3624
rect 9968 3596 9996 3624
rect 11324 3621 11336 3655
rect 11370 3652 11382 3655
rect 11606 3652 11612 3664
rect 11370 3624 11612 3652
rect 11370 3621 11382 3624
rect 11324 3615 11382 3621
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 14277 3655 14335 3661
rect 14277 3652 14289 3655
rect 11716 3624 14289 3652
rect 8570 3593 8576 3596
rect 6457 3587 6515 3593
rect 6457 3584 6469 3587
rect 6420 3556 6469 3584
rect 6420 3544 6426 3556
rect 6457 3553 6469 3556
rect 6503 3553 6515 3587
rect 6457 3547 6515 3553
rect 8297 3587 8355 3593
rect 8297 3553 8309 3587
rect 8343 3553 8355 3587
rect 8564 3584 8576 3593
rect 8531 3556 8576 3584
rect 8297 3547 8355 3553
rect 8564 3547 8576 3556
rect 8570 3544 8576 3547
rect 8628 3544 8634 3596
rect 9950 3544 9956 3596
rect 10008 3584 10014 3596
rect 10962 3584 10968 3596
rect 10008 3556 10968 3584
rect 10008 3544 10014 3556
rect 10962 3544 10968 3556
rect 11020 3584 11026 3596
rect 11057 3587 11115 3593
rect 11057 3584 11069 3587
rect 11020 3556 11069 3584
rect 11020 3544 11026 3556
rect 11057 3553 11069 3556
rect 11103 3553 11115 3587
rect 11716 3584 11744 3624
rect 14277 3621 14289 3624
rect 14323 3621 14335 3655
rect 15120 3652 15148 3692
rect 15930 3680 15936 3692
rect 15988 3720 15994 3732
rect 18693 3723 18751 3729
rect 15988 3692 18092 3720
rect 15988 3680 15994 3692
rect 14277 3615 14335 3621
rect 14384 3624 15148 3652
rect 11057 3547 11115 3553
rect 11164 3556 11744 3584
rect 3384 3488 3832 3516
rect 3384 3476 3390 3488
rect 10134 3476 10140 3528
rect 10192 3476 10198 3528
rect 11164 3516 11192 3556
rect 12158 3544 12164 3596
rect 12216 3584 12222 3596
rect 12216 3556 12664 3584
rect 12216 3544 12222 3556
rect 10244 3488 11192 3516
rect 12529 3519 12587 3525
rect 5166 3408 5172 3460
rect 5224 3448 5230 3460
rect 5442 3448 5448 3460
rect 5224 3420 5448 3448
rect 5224 3408 5230 3420
rect 5442 3408 5448 3420
rect 5500 3448 5506 3460
rect 10244 3448 10272 3488
rect 12529 3485 12541 3519
rect 12575 3485 12587 3519
rect 12636 3516 12664 3556
rect 12710 3544 12716 3596
rect 12768 3544 12774 3596
rect 14384 3593 14412 3624
rect 15194 3612 15200 3664
rect 15252 3652 15258 3664
rect 15252 3624 18000 3652
rect 15252 3612 15258 3624
rect 14369 3587 14427 3593
rect 12820 3556 14320 3584
rect 12820 3516 12848 3556
rect 14292 3528 14320 3556
rect 14369 3553 14381 3587
rect 14415 3553 14427 3587
rect 14369 3547 14427 3553
rect 15102 3544 15108 3596
rect 15160 3544 15166 3596
rect 16117 3587 16175 3593
rect 16117 3584 16129 3587
rect 15212 3556 16129 3584
rect 12636 3488 12848 3516
rect 12529 3479 12587 3485
rect 5500 3420 6316 3448
rect 5500 3408 5506 3420
rect 3513 3383 3571 3389
rect 3513 3349 3525 3383
rect 3559 3380 3571 3383
rect 3602 3380 3608 3392
rect 3559 3352 3608 3380
rect 3559 3349 3571 3352
rect 3513 3343 3571 3349
rect 3602 3340 3608 3352
rect 3660 3340 3666 3392
rect 5534 3340 5540 3392
rect 5592 3380 5598 3392
rect 6178 3380 6184 3392
rect 5592 3352 6184 3380
rect 5592 3340 5598 3352
rect 6178 3340 6184 3352
rect 6236 3340 6242 3392
rect 6288 3380 6316 3420
rect 9232 3420 10272 3448
rect 12544 3448 12572 3479
rect 12894 3476 12900 3528
rect 12952 3476 12958 3528
rect 14274 3476 14280 3528
rect 14332 3476 14338 3528
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 15212 3525 15240 3556
rect 16117 3553 16129 3556
rect 16163 3584 16175 3587
rect 16163 3556 16252 3584
rect 16163 3553 16175 3556
rect 16117 3547 16175 3553
rect 15197 3519 15255 3525
rect 14608 3488 15148 3516
rect 14608 3476 14614 3488
rect 12912 3448 12940 3476
rect 12544 3420 12940 3448
rect 15120 3448 15148 3488
rect 15197 3485 15209 3519
rect 15243 3485 15255 3519
rect 15197 3479 15255 3485
rect 15289 3519 15347 3525
rect 15289 3485 15301 3519
rect 15335 3485 15347 3519
rect 15289 3479 15347 3485
rect 15304 3448 15332 3479
rect 15120 3420 15332 3448
rect 16224 3448 16252 3556
rect 16298 3544 16304 3596
rect 16356 3544 16362 3596
rect 16390 3544 16396 3596
rect 16448 3544 16454 3596
rect 16485 3587 16543 3593
rect 16485 3553 16497 3587
rect 16531 3584 16543 3587
rect 16574 3584 16580 3596
rect 16531 3556 16580 3584
rect 16531 3553 16543 3556
rect 16485 3547 16543 3553
rect 16574 3544 16580 3556
rect 16632 3544 16638 3596
rect 17770 3544 17776 3596
rect 17828 3544 17834 3596
rect 17972 3593 18000 3624
rect 17957 3587 18015 3593
rect 17957 3553 17969 3587
rect 18003 3553 18015 3587
rect 17957 3547 18015 3553
rect 18064 3516 18092 3692
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 18782 3720 18788 3732
rect 18739 3692 18788 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 18782 3680 18788 3692
rect 18840 3680 18846 3732
rect 18969 3723 19027 3729
rect 18969 3689 18981 3723
rect 19015 3689 19027 3723
rect 18969 3683 19027 3689
rect 18322 3612 18328 3664
rect 18380 3652 18386 3664
rect 18984 3652 19012 3683
rect 19306 3655 19364 3661
rect 19306 3652 19318 3655
rect 18380 3624 18828 3652
rect 18984 3624 19318 3652
rect 18380 3612 18386 3624
rect 18506 3544 18512 3596
rect 18564 3544 18570 3596
rect 18800 3593 18828 3624
rect 19306 3621 19318 3624
rect 19352 3621 19364 3655
rect 19306 3615 19364 3621
rect 18785 3587 18843 3593
rect 18785 3553 18797 3587
rect 18831 3553 18843 3587
rect 18785 3547 18843 3553
rect 19058 3544 19064 3596
rect 19116 3544 19122 3596
rect 21450 3584 21456 3596
rect 19168 3556 21456 3584
rect 19168 3516 19196 3556
rect 21450 3544 21456 3556
rect 21508 3544 21514 3596
rect 18064 3488 19196 3516
rect 18046 3448 18052 3460
rect 16224 3420 18052 3448
rect 7466 3380 7472 3392
rect 6288 3352 7472 3380
rect 7466 3340 7472 3352
rect 7524 3380 7530 3392
rect 8202 3380 8208 3392
rect 7524 3352 8208 3380
rect 7524 3340 7530 3352
rect 8202 3340 8208 3352
rect 8260 3340 8266 3392
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 9232 3380 9260 3420
rect 12820 3392 12848 3420
rect 18046 3408 18052 3420
rect 18104 3408 18110 3460
rect 8352 3352 9260 3380
rect 9677 3383 9735 3389
rect 8352 3340 8358 3352
rect 9677 3349 9689 3383
rect 9723 3380 9735 3383
rect 9858 3380 9864 3392
rect 9723 3352 9864 3380
rect 9723 3349 9735 3352
rect 9677 3343 9735 3349
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 12802 3340 12808 3392
rect 12860 3340 12866 3392
rect 12894 3340 12900 3392
rect 12952 3340 12958 3392
rect 13354 3340 13360 3392
rect 13412 3380 13418 3392
rect 16206 3380 16212 3392
rect 13412 3352 16212 3380
rect 13412 3340 13418 3352
rect 16206 3340 16212 3352
rect 16264 3340 16270 3392
rect 16390 3340 16396 3392
rect 16448 3380 16454 3392
rect 16574 3380 16580 3392
rect 16448 3352 16580 3380
rect 16448 3340 16454 3352
rect 16574 3340 16580 3352
rect 16632 3340 16638 3392
rect 16669 3383 16727 3389
rect 16669 3349 16681 3383
rect 16715 3380 16727 3383
rect 17034 3380 17040 3392
rect 16715 3352 17040 3380
rect 16715 3349 16727 3352
rect 16669 3343 16727 3349
rect 17034 3340 17040 3352
rect 17092 3340 17098 3392
rect 18141 3383 18199 3389
rect 18141 3349 18153 3383
rect 18187 3380 18199 3383
rect 18322 3380 18328 3392
rect 18187 3352 18328 3380
rect 18187 3349 18199 3352
rect 18141 3343 18199 3349
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 18598 3340 18604 3392
rect 18656 3380 18662 3392
rect 19978 3380 19984 3392
rect 18656 3352 19984 3380
rect 18656 3340 18662 3352
rect 19978 3340 19984 3352
rect 20036 3380 20042 3392
rect 20441 3383 20499 3389
rect 20441 3380 20453 3383
rect 20036 3352 20453 3380
rect 20036 3340 20042 3352
rect 20441 3349 20453 3352
rect 20487 3349 20499 3383
rect 20441 3343 20499 3349
rect 552 3290 27416 3312
rect 552 3238 3756 3290
rect 3808 3238 3820 3290
rect 3872 3238 3884 3290
rect 3936 3238 3948 3290
rect 4000 3238 4012 3290
rect 4064 3238 10472 3290
rect 10524 3238 10536 3290
rect 10588 3238 10600 3290
rect 10652 3238 10664 3290
rect 10716 3238 10728 3290
rect 10780 3238 17188 3290
rect 17240 3238 17252 3290
rect 17304 3238 17316 3290
rect 17368 3238 17380 3290
rect 17432 3238 17444 3290
rect 17496 3238 23904 3290
rect 23956 3238 23968 3290
rect 24020 3238 24032 3290
rect 24084 3238 24096 3290
rect 24148 3238 24160 3290
rect 24212 3238 27416 3290
rect 552 3216 27416 3238
rect 4709 3179 4767 3185
rect 4709 3145 4721 3179
rect 4755 3176 4767 3179
rect 5534 3176 5540 3188
rect 4755 3148 5540 3176
rect 4755 3145 4767 3148
rect 4709 3139 4767 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 5776 3148 9720 3176
rect 5776 3136 5782 3148
rect 4798 3068 4804 3120
rect 4856 3108 4862 3120
rect 4856 3080 6040 3108
rect 4856 3068 4862 3080
rect 3326 3000 3332 3052
rect 3384 3000 3390 3052
rect 3602 2981 3608 2984
rect 3596 2972 3608 2981
rect 3563 2944 3608 2972
rect 3596 2935 3608 2944
rect 3602 2932 3608 2935
rect 3660 2932 3666 2984
rect 5166 2932 5172 2984
rect 5224 2972 5230 2984
rect 5261 2975 5319 2981
rect 5261 2972 5273 2975
rect 5224 2944 5273 2972
rect 5224 2932 5230 2944
rect 5261 2941 5273 2944
rect 5307 2941 5319 2975
rect 5261 2935 5319 2941
rect 5353 2975 5411 2981
rect 5353 2941 5365 2975
rect 5399 2972 5411 2975
rect 5534 2972 5540 2984
rect 5399 2944 5540 2972
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 5534 2932 5540 2944
rect 5592 2932 5598 2984
rect 5629 2975 5687 2981
rect 5629 2941 5641 2975
rect 5675 2941 5687 2975
rect 5629 2935 5687 2941
rect 5442 2864 5448 2916
rect 5500 2864 5506 2916
rect 5644 2904 5672 2935
rect 5718 2932 5724 2984
rect 5776 2932 5782 2984
rect 5902 2932 5908 2984
rect 5960 2932 5966 2984
rect 6012 2981 6040 3080
rect 7834 3068 7840 3120
rect 7892 3068 7898 3120
rect 9692 3108 9720 3148
rect 10134 3136 10140 3188
rect 10192 3136 10198 3188
rect 15102 3176 15108 3188
rect 10244 3148 15108 3176
rect 10244 3108 10272 3148
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 15654 3136 15660 3188
rect 15712 3176 15718 3188
rect 15933 3179 15991 3185
rect 15933 3176 15945 3179
rect 15712 3148 15945 3176
rect 15712 3136 15718 3148
rect 15933 3145 15945 3148
rect 15979 3145 15991 3179
rect 15933 3139 15991 3145
rect 16022 3136 16028 3188
rect 16080 3176 16086 3188
rect 18598 3176 18604 3188
rect 16080 3148 18604 3176
rect 16080 3136 16086 3148
rect 18598 3136 18604 3148
rect 18656 3136 18662 3188
rect 19058 3176 19064 3188
rect 18708 3148 19064 3176
rect 12434 3108 12440 3120
rect 9692 3080 10272 3108
rect 12360 3080 12440 3108
rect 7852 3040 7880 3068
rect 7576 3012 7880 3040
rect 5997 2975 6055 2981
rect 5997 2941 6009 2975
rect 6043 2941 6055 2975
rect 5997 2935 6055 2941
rect 6089 2975 6147 2981
rect 6089 2941 6101 2975
rect 6135 2972 6147 2975
rect 7466 2972 7472 2984
rect 6135 2944 7472 2972
rect 6135 2941 6147 2944
rect 6089 2935 6147 2941
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 7576 2981 7604 3012
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2941 7619 2975
rect 7561 2935 7619 2941
rect 7837 2975 7895 2981
rect 7837 2941 7849 2975
rect 7883 2972 7895 2975
rect 8294 2972 8300 2984
rect 7883 2944 8300 2972
rect 7883 2941 7895 2944
rect 7837 2935 7895 2941
rect 8294 2932 8300 2944
rect 8352 2932 8358 2984
rect 8757 2975 8815 2981
rect 8757 2941 8769 2975
rect 8803 2972 8815 2975
rect 9950 2972 9956 2984
rect 8803 2944 9956 2972
rect 8803 2941 8815 2944
rect 8757 2935 8815 2941
rect 9950 2932 9956 2944
rect 10008 2932 10014 2984
rect 12066 2932 12072 2984
rect 12124 2932 12130 2984
rect 12360 2981 12388 3080
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 14642 3068 14648 3120
rect 14700 3108 14706 3120
rect 14700 3080 18644 3108
rect 14700 3068 14706 3080
rect 13722 3040 13728 3052
rect 12728 3012 13728 3040
rect 12728 2984 12756 3012
rect 13722 3000 13728 3012
rect 13780 3040 13786 3052
rect 15010 3040 15016 3052
rect 13780 3012 15016 3040
rect 13780 3000 13786 3012
rect 15010 3000 15016 3012
rect 15068 3000 15074 3052
rect 15289 3043 15347 3049
rect 15289 3009 15301 3043
rect 15335 3009 15347 3043
rect 16298 3040 16304 3052
rect 15289 3003 15347 3009
rect 16224 3012 16304 3040
rect 12345 2975 12403 2981
rect 12345 2941 12357 2975
rect 12391 2941 12403 2975
rect 12345 2935 12403 2941
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 12710 2972 12716 2984
rect 12483 2944 12716 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 12894 2932 12900 2984
rect 12952 2932 12958 2984
rect 14550 2932 14556 2984
rect 14608 2972 14614 2984
rect 15304 2972 15332 3003
rect 14608 2944 15332 2972
rect 15473 2975 15531 2981
rect 14608 2932 14614 2944
rect 15473 2941 15485 2975
rect 15519 2972 15531 2975
rect 16022 2972 16028 2984
rect 15519 2944 16028 2972
rect 15519 2941 15531 2944
rect 15473 2935 15531 2941
rect 16022 2932 16028 2944
rect 16080 2932 16086 2984
rect 16224 2981 16252 3012
rect 16298 3000 16304 3012
rect 16356 3000 16362 3052
rect 17497 3043 17555 3049
rect 16592 3012 16896 3040
rect 16209 2975 16267 2981
rect 16209 2941 16221 2975
rect 16255 2941 16267 2975
rect 16209 2935 16267 2941
rect 16390 2932 16396 2984
rect 16448 2932 16454 2984
rect 7653 2907 7711 2913
rect 5644 2876 7604 2904
rect 5644 2848 5672 2876
rect 5074 2796 5080 2848
rect 5132 2796 5138 2848
rect 5626 2796 5632 2848
rect 5684 2796 5690 2848
rect 6270 2796 6276 2848
rect 6328 2796 6334 2848
rect 7285 2839 7343 2845
rect 7285 2805 7297 2839
rect 7331 2836 7343 2839
rect 7466 2836 7472 2848
rect 7331 2808 7472 2836
rect 7331 2805 7343 2808
rect 7285 2799 7343 2805
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 7576 2836 7604 2876
rect 7653 2873 7665 2907
rect 7699 2904 7711 2907
rect 8018 2904 8024 2916
rect 7699 2876 8024 2904
rect 7699 2873 7711 2876
rect 7653 2867 7711 2873
rect 8018 2864 8024 2876
rect 8076 2864 8082 2916
rect 9024 2907 9082 2913
rect 9024 2873 9036 2907
rect 9070 2904 9082 2907
rect 10042 2904 10048 2916
rect 9070 2876 10048 2904
rect 9070 2873 9082 2876
rect 9024 2867 9082 2873
rect 10042 2864 10048 2876
rect 10100 2864 10106 2916
rect 12250 2864 12256 2916
rect 12308 2864 12314 2916
rect 15565 2907 15623 2913
rect 15565 2904 15577 2907
rect 12360 2876 15577 2904
rect 12360 2836 12388 2876
rect 15565 2873 15577 2876
rect 15611 2873 15623 2907
rect 15565 2867 15623 2873
rect 16114 2864 16120 2916
rect 16172 2904 16178 2916
rect 16301 2907 16359 2913
rect 16301 2904 16313 2907
rect 16172 2876 16313 2904
rect 16172 2864 16178 2876
rect 16301 2873 16313 2876
rect 16347 2873 16359 2907
rect 16301 2867 16359 2873
rect 7576 2808 12388 2836
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12621 2839 12679 2845
rect 12621 2836 12633 2839
rect 12492 2808 12633 2836
rect 12492 2796 12498 2808
rect 12621 2805 12633 2808
rect 12667 2805 12679 2839
rect 12621 2799 12679 2805
rect 12710 2796 12716 2848
rect 12768 2796 12774 2848
rect 16592 2845 16620 3012
rect 16868 2981 16896 3012
rect 17497 3009 17509 3043
rect 17543 3040 17555 3043
rect 17770 3040 17776 3052
rect 17543 3012 17776 3040
rect 17543 3009 17555 3012
rect 17497 3003 17555 3009
rect 16761 2975 16819 2981
rect 16761 2941 16773 2975
rect 16807 2941 16819 2975
rect 16761 2935 16819 2941
rect 16853 2975 16911 2981
rect 16853 2941 16865 2975
rect 16899 2941 16911 2975
rect 16853 2935 16911 2941
rect 16776 2904 16804 2935
rect 17034 2932 17040 2984
rect 17092 2972 17098 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 17092 2944 17325 2972
rect 17092 2932 17098 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 17512 2904 17540 3003
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 18322 2932 18328 2984
rect 18380 2932 18386 2984
rect 18616 2972 18644 3080
rect 18708 3049 18736 3148
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 19886 3108 19892 3120
rect 19720 3080 19892 3108
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3009 18751 3043
rect 18693 3003 18751 3009
rect 19720 2972 19748 3080
rect 19886 3068 19892 3080
rect 19944 3108 19950 3120
rect 20073 3111 20131 3117
rect 20073 3108 20085 3111
rect 19944 3080 20085 3108
rect 19944 3068 19950 3080
rect 20073 3077 20085 3080
rect 20119 3077 20131 3111
rect 20073 3071 20131 3077
rect 18616 2944 19748 2972
rect 18938 2907 18996 2913
rect 18938 2904 18950 2907
rect 16776 2876 17540 2904
rect 18524 2876 18950 2904
rect 16577 2839 16635 2845
rect 16577 2805 16589 2839
rect 16623 2805 16635 2839
rect 16577 2799 16635 2805
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 17037 2839 17095 2845
rect 17037 2836 17049 2839
rect 16816 2808 17049 2836
rect 16816 2796 16822 2808
rect 17037 2805 17049 2808
rect 17083 2805 17095 2839
rect 17037 2799 17095 2805
rect 17129 2839 17187 2845
rect 17129 2805 17141 2839
rect 17175 2836 17187 2839
rect 17218 2836 17224 2848
rect 17175 2808 17224 2836
rect 17175 2805 17187 2808
rect 17129 2799 17187 2805
rect 17218 2796 17224 2808
rect 17276 2796 17282 2848
rect 18524 2845 18552 2876
rect 18938 2873 18950 2876
rect 18984 2873 18996 2907
rect 18938 2867 18996 2873
rect 18509 2839 18567 2845
rect 18509 2805 18521 2839
rect 18555 2805 18567 2839
rect 18509 2799 18567 2805
rect 552 2746 27576 2768
rect 552 2694 7114 2746
rect 7166 2694 7178 2746
rect 7230 2694 7242 2746
rect 7294 2694 7306 2746
rect 7358 2694 7370 2746
rect 7422 2694 13830 2746
rect 13882 2694 13894 2746
rect 13946 2694 13958 2746
rect 14010 2694 14022 2746
rect 14074 2694 14086 2746
rect 14138 2694 20546 2746
rect 20598 2694 20610 2746
rect 20662 2694 20674 2746
rect 20726 2694 20738 2746
rect 20790 2694 20802 2746
rect 20854 2694 27262 2746
rect 27314 2694 27326 2746
rect 27378 2694 27390 2746
rect 27442 2694 27454 2746
rect 27506 2694 27518 2746
rect 27570 2694 27576 2746
rect 552 2672 27576 2694
rect 5169 2635 5227 2641
rect 5169 2601 5181 2635
rect 5215 2632 5227 2635
rect 5718 2632 5724 2644
rect 5215 2604 5724 2632
rect 5215 2601 5227 2604
rect 5169 2595 5227 2601
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 9324 2604 9996 2632
rect 5629 2567 5687 2573
rect 5629 2533 5641 2567
rect 5675 2564 5687 2567
rect 5675 2536 6500 2564
rect 5675 2533 5687 2536
rect 5629 2527 5687 2533
rect 3602 2456 3608 2508
rect 3660 2496 3666 2508
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 3660 2468 3801 2496
rect 3660 2456 3666 2468
rect 3789 2465 3801 2468
rect 3835 2465 3847 2499
rect 3789 2459 3847 2465
rect 4056 2499 4114 2505
rect 4056 2465 4068 2499
rect 4102 2496 4114 2499
rect 4338 2496 4344 2508
rect 4102 2468 4344 2496
rect 4102 2465 4114 2468
rect 4056 2459 4114 2465
rect 4338 2456 4344 2468
rect 4396 2456 4402 2508
rect 5074 2456 5080 2508
rect 5132 2496 5138 2508
rect 5445 2499 5503 2505
rect 5445 2496 5457 2499
rect 5132 2468 5457 2496
rect 5132 2456 5138 2468
rect 5445 2465 5457 2468
rect 5491 2465 5503 2499
rect 5445 2459 5503 2465
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2496 6055 2499
rect 6270 2496 6276 2508
rect 6043 2468 6276 2496
rect 6043 2465 6055 2468
rect 5997 2459 6055 2465
rect 6270 2456 6276 2468
rect 6328 2456 6334 2508
rect 6472 2505 6500 2536
rect 6457 2499 6515 2505
rect 6457 2465 6469 2499
rect 6503 2465 6515 2499
rect 6457 2459 6515 2465
rect 7466 2456 7472 2508
rect 7524 2496 7530 2508
rect 7561 2499 7619 2505
rect 7561 2496 7573 2499
rect 7524 2468 7573 2496
rect 7524 2456 7530 2468
rect 7561 2465 7573 2468
rect 7607 2465 7619 2499
rect 7561 2459 7619 2465
rect 8202 2456 8208 2508
rect 8260 2496 8266 2508
rect 8849 2499 8907 2505
rect 8260 2468 8800 2496
rect 8260 2456 8266 2468
rect 5258 2388 5264 2440
rect 5316 2428 5322 2440
rect 6181 2431 6239 2437
rect 6181 2428 6193 2431
rect 5316 2400 6193 2428
rect 5316 2388 5322 2400
rect 6181 2397 6193 2400
rect 6227 2428 6239 2431
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 6227 2400 7389 2428
rect 6227 2397 6239 2400
rect 6181 2391 6239 2397
rect 7377 2397 7389 2400
rect 7423 2428 7435 2431
rect 8662 2428 8668 2440
rect 7423 2400 8668 2428
rect 7423 2397 7435 2400
rect 7377 2391 7435 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 8772 2428 8800 2468
rect 8849 2465 8861 2499
rect 8895 2496 8907 2499
rect 9140 2496 9168 2595
rect 9324 2505 9352 2604
rect 9401 2567 9459 2573
rect 9401 2533 9413 2567
rect 9447 2564 9459 2567
rect 9858 2564 9864 2576
rect 9447 2536 9864 2564
rect 9447 2533 9459 2536
rect 9401 2527 9459 2533
rect 9858 2524 9864 2536
rect 9916 2524 9922 2576
rect 8895 2468 9168 2496
rect 9309 2499 9367 2505
rect 8895 2465 8907 2468
rect 8849 2459 8907 2465
rect 9309 2465 9321 2499
rect 9355 2465 9367 2499
rect 9309 2459 9367 2465
rect 9493 2499 9551 2505
rect 9493 2465 9505 2499
rect 9539 2465 9551 2499
rect 9493 2459 9551 2465
rect 9677 2499 9735 2505
rect 9677 2465 9689 2499
rect 9723 2496 9735 2499
rect 9766 2496 9772 2508
rect 9723 2468 9772 2496
rect 9723 2465 9735 2468
rect 9677 2459 9735 2465
rect 9324 2428 9352 2459
rect 8772 2400 9352 2428
rect 9508 2428 9536 2459
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 9968 2505 9996 2604
rect 10134 2592 10140 2644
rect 10192 2592 10198 2644
rect 12250 2632 12256 2644
rect 10244 2604 12256 2632
rect 10045 2567 10103 2573
rect 10045 2533 10057 2567
rect 10091 2564 10103 2567
rect 10152 2564 10180 2592
rect 10091 2536 10180 2564
rect 10091 2533 10103 2536
rect 10045 2527 10103 2533
rect 9953 2499 10011 2505
rect 9953 2465 9965 2499
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 10137 2499 10195 2505
rect 10137 2465 10149 2499
rect 10183 2496 10195 2499
rect 10244 2496 10272 2604
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 12802 2592 12808 2644
rect 12860 2632 12866 2644
rect 13078 2632 13084 2644
rect 12860 2604 13084 2632
rect 12860 2592 12866 2604
rect 13078 2592 13084 2604
rect 13136 2632 13142 2644
rect 13265 2635 13323 2641
rect 13265 2632 13277 2635
rect 13136 2604 13277 2632
rect 13136 2592 13142 2604
rect 13265 2601 13277 2604
rect 13311 2601 13323 2635
rect 13265 2595 13323 2601
rect 14642 2592 14648 2644
rect 14700 2592 14706 2644
rect 12152 2567 12210 2573
rect 12152 2533 12164 2567
rect 12198 2564 12210 2567
rect 12710 2564 12716 2576
rect 12198 2536 12716 2564
rect 12198 2533 12210 2536
rect 12152 2527 12210 2533
rect 12710 2524 12716 2536
rect 12768 2524 12774 2576
rect 13722 2524 13728 2576
rect 13780 2564 13786 2576
rect 14369 2567 14427 2573
rect 13780 2536 14228 2564
rect 13780 2524 13786 2536
rect 10183 2468 10272 2496
rect 10183 2465 10195 2468
rect 10137 2459 10195 2465
rect 9508 2400 9674 2428
rect 5442 2320 5448 2372
rect 5500 2360 5506 2372
rect 5902 2360 5908 2372
rect 5500 2332 5908 2360
rect 5500 2320 5506 2332
rect 5902 2320 5908 2332
rect 5960 2360 5966 2372
rect 6914 2360 6920 2372
rect 5960 2332 6920 2360
rect 5960 2320 5966 2332
rect 6914 2320 6920 2332
rect 6972 2360 6978 2372
rect 8018 2360 8024 2372
rect 6972 2332 8024 2360
rect 6972 2320 6978 2332
rect 8018 2320 8024 2332
rect 8076 2360 8082 2372
rect 9646 2360 9674 2400
rect 10152 2360 10180 2459
rect 10318 2456 10324 2508
rect 10376 2456 10382 2508
rect 10962 2456 10968 2508
rect 11020 2496 11026 2508
rect 14200 2505 14228 2536
rect 14369 2533 14381 2567
rect 14415 2564 14427 2567
rect 14918 2564 14924 2576
rect 14415 2536 14924 2564
rect 14415 2533 14427 2536
rect 14369 2527 14427 2533
rect 14918 2524 14924 2536
rect 14976 2524 14982 2576
rect 16574 2524 16580 2576
rect 16632 2524 16638 2576
rect 14185 2499 14243 2505
rect 11020 2468 13851 2496
rect 11020 2456 11026 2468
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 11882 2428 11888 2440
rect 10284 2400 11888 2428
rect 10284 2388 10290 2400
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 13823 2428 13851 2468
rect 14185 2465 14197 2499
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 14292 2428 14320 2459
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 14553 2499 14611 2505
rect 14553 2496 14565 2499
rect 14516 2468 14565 2496
rect 14516 2456 14522 2468
rect 14553 2465 14565 2468
rect 14599 2465 14611 2499
rect 14553 2459 14611 2465
rect 13823 2400 14320 2428
rect 14568 2428 14596 2459
rect 15010 2456 15016 2508
rect 15068 2456 15074 2508
rect 16758 2456 16764 2508
rect 16816 2456 16822 2508
rect 17218 2456 17224 2508
rect 17276 2456 17282 2508
rect 15105 2431 15163 2437
rect 15105 2428 15117 2431
rect 14568 2400 15117 2428
rect 15105 2397 15117 2400
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15378 2428 15384 2440
rect 15335 2400 15384 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15378 2388 15384 2400
rect 15436 2428 15442 2440
rect 16298 2428 16304 2440
rect 15436 2400 16304 2428
rect 15436 2388 15442 2400
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 14182 2360 14188 2372
rect 8076 2332 10180 2360
rect 12820 2332 14188 2360
rect 8076 2320 8082 2332
rect 5810 2252 5816 2304
rect 5868 2252 5874 2304
rect 6270 2252 6276 2304
rect 6328 2252 6334 2304
rect 7650 2252 7656 2304
rect 7708 2292 7714 2304
rect 7745 2295 7803 2301
rect 7745 2292 7757 2295
rect 7708 2264 7757 2292
rect 7708 2252 7714 2264
rect 7745 2261 7757 2264
rect 7791 2261 7803 2295
rect 7745 2255 7803 2261
rect 8938 2252 8944 2304
rect 8996 2292 9002 2304
rect 9033 2295 9091 2301
rect 9033 2292 9045 2295
rect 8996 2264 9045 2292
rect 8996 2252 9002 2264
rect 9033 2261 9045 2264
rect 9079 2261 9091 2295
rect 9033 2255 9091 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9769 2295 9827 2301
rect 9769 2292 9781 2295
rect 9732 2264 9781 2292
rect 9732 2252 9738 2264
rect 9769 2261 9781 2264
rect 9815 2261 9827 2295
rect 9769 2255 9827 2261
rect 9858 2252 9864 2304
rect 9916 2292 9922 2304
rect 10870 2292 10876 2304
rect 9916 2264 10876 2292
rect 9916 2252 9922 2264
rect 10870 2252 10876 2264
rect 10928 2292 10934 2304
rect 12820 2292 12848 2332
rect 14182 2320 14188 2332
rect 14240 2320 14246 2372
rect 10928 2264 12848 2292
rect 10928 2252 10934 2264
rect 13906 2252 13912 2304
rect 13964 2292 13970 2304
rect 14001 2295 14059 2301
rect 14001 2292 14013 2295
rect 13964 2264 14013 2292
rect 13964 2252 13970 2264
rect 14001 2261 14013 2264
rect 14047 2261 14059 2295
rect 14001 2255 14059 2261
rect 16942 2252 16948 2304
rect 17000 2252 17006 2304
rect 17034 2252 17040 2304
rect 17092 2252 17098 2304
rect 552 2202 27416 2224
rect 552 2150 3756 2202
rect 3808 2150 3820 2202
rect 3872 2150 3884 2202
rect 3936 2150 3948 2202
rect 4000 2150 4012 2202
rect 4064 2150 10472 2202
rect 10524 2150 10536 2202
rect 10588 2150 10600 2202
rect 10652 2150 10664 2202
rect 10716 2150 10728 2202
rect 10780 2150 17188 2202
rect 17240 2150 17252 2202
rect 17304 2150 17316 2202
rect 17368 2150 17380 2202
rect 17432 2150 17444 2202
rect 17496 2150 23904 2202
rect 23956 2150 23968 2202
rect 24020 2150 24032 2202
rect 24084 2150 24096 2202
rect 24148 2150 24160 2202
rect 24212 2150 27416 2202
rect 552 2128 27416 2150
rect 4338 2048 4344 2100
rect 4396 2048 4402 2100
rect 10318 2048 10324 2100
rect 10376 2088 10382 2100
rect 11333 2091 11391 2097
rect 11333 2088 11345 2091
rect 10376 2060 11345 2088
rect 10376 2048 10382 2060
rect 11333 2057 11345 2060
rect 11379 2088 11391 2091
rect 11379 2060 12434 2088
rect 11379 2057 11391 2060
rect 11333 2051 11391 2057
rect 6362 1912 6368 1964
rect 6420 1912 6426 1964
rect 8662 1912 8668 1964
rect 8720 1952 8726 1964
rect 9950 1961 9956 1964
rect 9942 1955 9956 1961
rect 8720 1924 9904 1952
rect 8720 1912 8726 1924
rect 4525 1887 4583 1893
rect 4525 1853 4537 1887
rect 4571 1884 4583 1887
rect 5810 1884 5816 1896
rect 4571 1856 5816 1884
rect 4571 1853 4583 1856
rect 4525 1847 4583 1853
rect 5810 1844 5816 1856
rect 5868 1844 5874 1896
rect 6109 1887 6167 1893
rect 6109 1853 6121 1887
rect 6155 1884 6167 1887
rect 6270 1884 6276 1896
rect 6155 1856 6276 1884
rect 6155 1853 6167 1856
rect 6109 1847 6167 1853
rect 6270 1844 6276 1856
rect 6328 1844 6334 1896
rect 7650 1844 7656 1896
rect 7708 1844 7714 1896
rect 8938 1844 8944 1896
rect 8996 1844 9002 1896
rect 9217 1887 9275 1893
rect 9217 1853 9229 1887
rect 9263 1884 9275 1887
rect 9493 1887 9551 1893
rect 9493 1884 9505 1887
rect 9263 1856 9505 1884
rect 9263 1853 9275 1856
rect 9217 1847 9275 1853
rect 9493 1853 9505 1856
rect 9539 1853 9551 1887
rect 9493 1847 9551 1853
rect 9674 1844 9680 1896
rect 9732 1844 9738 1896
rect 9876 1893 9904 1924
rect 9942 1921 9954 1955
rect 10008 1952 10014 1964
rect 12406 1952 12434 2060
rect 15010 2020 15016 2032
rect 14200 1992 15016 2020
rect 14200 1961 14228 1992
rect 15010 1980 15016 1992
rect 15068 1980 15074 2032
rect 15286 1980 15292 2032
rect 15344 1980 15350 2032
rect 14185 1955 14243 1961
rect 14185 1952 14197 1955
rect 10008 1924 10042 1952
rect 12406 1924 14197 1952
rect 9942 1915 9956 1921
rect 9950 1912 9956 1915
rect 10008 1912 10014 1924
rect 14185 1921 14197 1924
rect 14231 1921 14243 1955
rect 14185 1915 14243 1921
rect 18506 1912 18512 1964
rect 18564 1952 18570 1964
rect 18564 1924 19840 1952
rect 18564 1912 18570 1924
rect 19812 1896 19840 1924
rect 20254 1912 20260 1964
rect 20312 1912 20318 1964
rect 9861 1887 9919 1893
rect 9861 1853 9873 1887
rect 9907 1884 9919 1887
rect 12345 1887 12403 1893
rect 12345 1884 12357 1887
rect 9907 1880 9996 1884
rect 10060 1880 12357 1884
rect 9907 1856 12357 1880
rect 9907 1853 9919 1856
rect 9861 1847 9919 1853
rect 9968 1852 10088 1856
rect 12345 1853 12357 1856
rect 12391 1853 12403 1887
rect 12345 1847 12403 1853
rect 4890 1776 4896 1828
rect 4948 1816 4954 1828
rect 5994 1816 6000 1828
rect 4948 1788 6000 1816
rect 4948 1776 4954 1788
rect 5994 1776 6000 1788
rect 6052 1776 6058 1828
rect 10198 1819 10256 1825
rect 10198 1816 10210 1819
rect 9784 1788 10210 1816
rect 4985 1751 5043 1757
rect 4985 1717 4997 1751
rect 5031 1748 5043 1751
rect 5626 1748 5632 1760
rect 5031 1720 5632 1748
rect 5031 1717 5043 1720
rect 4985 1711 5043 1717
rect 5626 1708 5632 1720
rect 5684 1748 5690 1760
rect 6822 1748 6828 1760
rect 5684 1720 6828 1748
rect 5684 1708 5690 1720
rect 6822 1708 6828 1720
rect 6880 1708 6886 1760
rect 7469 1751 7527 1757
rect 7469 1717 7481 1751
rect 7515 1748 7527 1751
rect 7558 1748 7564 1760
rect 7515 1720 7564 1748
rect 7515 1717 7527 1720
rect 7469 1711 7527 1717
rect 7558 1708 7564 1720
rect 7616 1708 7622 1760
rect 9122 1708 9128 1760
rect 9180 1708 9186 1760
rect 9401 1751 9459 1757
rect 9401 1717 9413 1751
rect 9447 1748 9459 1751
rect 9784 1748 9812 1788
rect 10198 1785 10210 1788
rect 10244 1785 10256 1819
rect 10198 1779 10256 1785
rect 11514 1776 11520 1828
rect 11572 1816 11578 1828
rect 12066 1816 12072 1828
rect 11572 1788 12072 1816
rect 11572 1776 11578 1788
rect 12066 1776 12072 1788
rect 12124 1776 12130 1828
rect 12360 1816 12388 1847
rect 12434 1844 12440 1896
rect 12492 1844 12498 1896
rect 12621 1887 12679 1893
rect 12621 1853 12633 1887
rect 12667 1884 12679 1887
rect 12713 1887 12771 1893
rect 12713 1884 12725 1887
rect 12667 1856 12725 1884
rect 12667 1853 12679 1856
rect 12621 1847 12679 1853
rect 12713 1853 12725 1856
rect 12759 1853 12771 1887
rect 12713 1847 12771 1853
rect 12894 1844 12900 1896
rect 12952 1884 12958 1896
rect 13725 1887 13783 1893
rect 13725 1884 13737 1887
rect 12952 1856 13737 1884
rect 12952 1844 12958 1856
rect 13725 1853 13737 1856
rect 13771 1853 13783 1887
rect 13725 1847 13783 1853
rect 13906 1844 13912 1896
rect 13964 1844 13970 1896
rect 14366 1884 14372 1896
rect 14016 1856 14372 1884
rect 12912 1816 12940 1844
rect 12360 1788 12940 1816
rect 12986 1776 12992 1828
rect 13044 1816 13050 1828
rect 14016 1816 14044 1856
rect 14366 1844 14372 1856
rect 14424 1884 14430 1896
rect 14550 1884 14556 1896
rect 14424 1856 14556 1884
rect 14424 1844 14430 1856
rect 14550 1844 14556 1856
rect 14608 1844 14614 1896
rect 14921 1887 14979 1893
rect 14921 1853 14933 1887
rect 14967 1884 14979 1887
rect 15010 1884 15016 1896
rect 14967 1856 15016 1884
rect 14967 1853 14979 1856
rect 14921 1847 14979 1853
rect 15010 1844 15016 1856
rect 15068 1844 15074 1896
rect 15105 1887 15163 1893
rect 15105 1853 15117 1887
rect 15151 1884 15163 1887
rect 15378 1884 15384 1896
rect 15151 1856 15384 1884
rect 15151 1853 15163 1856
rect 15105 1847 15163 1853
rect 15378 1844 15384 1856
rect 15436 1844 15442 1896
rect 15841 1887 15899 1893
rect 15841 1853 15853 1887
rect 15887 1853 15899 1887
rect 15841 1847 15899 1853
rect 13044 1788 14044 1816
rect 14093 1819 14151 1825
rect 13044 1776 13050 1788
rect 14093 1785 14105 1819
rect 14139 1816 14151 1819
rect 15856 1816 15884 1847
rect 16758 1844 16764 1896
rect 16816 1884 16822 1896
rect 17405 1887 17463 1893
rect 17405 1884 17417 1887
rect 16816 1856 17417 1884
rect 16816 1844 16822 1856
rect 17405 1853 17417 1856
rect 17451 1884 17463 1887
rect 17862 1884 17868 1896
rect 17451 1856 17868 1884
rect 17451 1853 17463 1856
rect 17405 1847 17463 1853
rect 17862 1844 17868 1856
rect 17920 1844 17926 1896
rect 18414 1844 18420 1896
rect 18472 1884 18478 1896
rect 18874 1884 18880 1896
rect 18472 1856 18880 1884
rect 18472 1844 18478 1856
rect 18874 1844 18880 1856
rect 18932 1844 18938 1896
rect 19794 1844 19800 1896
rect 19852 1844 19858 1896
rect 19978 1844 19984 1896
rect 20036 1844 20042 1896
rect 20346 1844 20352 1896
rect 20404 1884 20410 1896
rect 21726 1884 21732 1896
rect 20404 1856 21732 1884
rect 20404 1844 20410 1856
rect 21726 1844 21732 1856
rect 21784 1844 21790 1896
rect 14139 1788 15884 1816
rect 14139 1785 14151 1788
rect 14093 1779 14151 1785
rect 16942 1776 16948 1828
rect 17000 1816 17006 1828
rect 17138 1819 17196 1825
rect 17138 1816 17150 1819
rect 17000 1788 17150 1816
rect 17000 1776 17006 1788
rect 17138 1785 17150 1788
rect 17184 1785 17196 1819
rect 17138 1779 17196 1785
rect 17954 1776 17960 1828
rect 18012 1816 18018 1828
rect 20993 1819 21051 1825
rect 18012 1788 18552 1816
rect 18012 1776 18018 1788
rect 9447 1720 9812 1748
rect 9447 1717 9459 1720
rect 9401 1711 9459 1717
rect 12894 1708 12900 1760
rect 12952 1708 12958 1760
rect 15654 1708 15660 1760
rect 15712 1708 15718 1760
rect 16022 1708 16028 1760
rect 16080 1748 16086 1760
rect 16390 1748 16396 1760
rect 16080 1720 16396 1748
rect 16080 1708 16086 1720
rect 16390 1708 16396 1720
rect 16448 1708 16454 1760
rect 16482 1708 16488 1760
rect 16540 1748 16546 1760
rect 18414 1748 18420 1760
rect 16540 1720 18420 1748
rect 16540 1708 16546 1720
rect 18414 1708 18420 1720
rect 18472 1708 18478 1760
rect 18524 1748 18552 1788
rect 20993 1785 21005 1819
rect 21039 1816 21051 1819
rect 23566 1816 23572 1828
rect 21039 1788 23572 1816
rect 21039 1785 21051 1788
rect 20993 1779 21051 1785
rect 23566 1776 23572 1788
rect 23624 1776 23630 1828
rect 21542 1748 21548 1760
rect 18524 1720 21548 1748
rect 21542 1708 21548 1720
rect 21600 1708 21606 1760
rect 552 1658 27576 1680
rect 552 1606 7114 1658
rect 7166 1606 7178 1658
rect 7230 1606 7242 1658
rect 7294 1606 7306 1658
rect 7358 1606 7370 1658
rect 7422 1606 13830 1658
rect 13882 1606 13894 1658
rect 13946 1606 13958 1658
rect 14010 1606 14022 1658
rect 14074 1606 14086 1658
rect 14138 1606 20546 1658
rect 20598 1606 20610 1658
rect 20662 1606 20674 1658
rect 20726 1606 20738 1658
rect 20790 1606 20802 1658
rect 20854 1606 27262 1658
rect 27314 1606 27326 1658
rect 27378 1606 27390 1658
rect 27442 1606 27454 1658
rect 27506 1606 27518 1658
rect 27570 1606 27576 1658
rect 552 1584 27576 1606
rect 2590 1504 2596 1556
rect 2648 1544 2654 1556
rect 5905 1547 5963 1553
rect 5905 1544 5917 1547
rect 2648 1516 5917 1544
rect 2648 1504 2654 1516
rect 5905 1513 5917 1516
rect 5951 1513 5963 1547
rect 6454 1544 6460 1556
rect 5905 1507 5963 1513
rect 6196 1516 6460 1544
rect 6196 1476 6224 1516
rect 6454 1504 6460 1516
rect 6512 1504 6518 1556
rect 8294 1504 8300 1556
rect 8352 1544 8358 1556
rect 8665 1547 8723 1553
rect 8665 1544 8677 1547
rect 8352 1516 8677 1544
rect 8352 1504 8358 1516
rect 8665 1513 8677 1516
rect 8711 1513 8723 1547
rect 8665 1507 8723 1513
rect 10689 1547 10747 1553
rect 10689 1513 10701 1547
rect 10735 1544 10747 1547
rect 10870 1544 10876 1556
rect 10735 1516 10876 1544
rect 10735 1513 10747 1516
rect 10689 1507 10747 1513
rect 10870 1504 10876 1516
rect 10928 1504 10934 1556
rect 11256 1516 11836 1544
rect 7742 1476 7748 1488
rect 5092 1448 6224 1476
rect 6288 1448 7748 1476
rect 4338 1368 4344 1420
rect 4396 1408 4402 1420
rect 4433 1411 4491 1417
rect 4433 1408 4445 1411
rect 4396 1380 4445 1408
rect 4396 1368 4402 1380
rect 4433 1377 4445 1380
rect 4479 1377 4491 1411
rect 4433 1371 4491 1377
rect 4890 1368 4896 1420
rect 4948 1368 4954 1420
rect 5092 1417 5120 1448
rect 5077 1411 5135 1417
rect 5077 1377 5089 1411
rect 5123 1377 5135 1411
rect 5077 1371 5135 1377
rect 5445 1411 5503 1417
rect 5445 1377 5457 1411
rect 5491 1408 5503 1411
rect 5718 1408 5724 1420
rect 5491 1380 5724 1408
rect 5491 1377 5503 1380
rect 5445 1371 5503 1377
rect 5718 1368 5724 1380
rect 5776 1368 5782 1420
rect 6288 1417 6316 1448
rect 7742 1436 7748 1448
rect 7800 1436 7806 1488
rect 9122 1436 9128 1488
rect 9180 1476 9186 1488
rect 9554 1479 9612 1485
rect 9554 1476 9566 1479
rect 9180 1448 9566 1476
rect 9180 1436 9186 1448
rect 9554 1445 9566 1448
rect 9600 1445 9612 1479
rect 9554 1439 9612 1445
rect 6273 1411 6331 1417
rect 6273 1377 6285 1411
rect 6319 1377 6331 1411
rect 6273 1371 6331 1377
rect 6454 1368 6460 1420
rect 6512 1368 6518 1420
rect 6822 1368 6828 1420
rect 6880 1368 6886 1420
rect 7558 1417 7564 1420
rect 7552 1408 7564 1417
rect 7519 1380 7564 1408
rect 7552 1371 7564 1380
rect 7558 1368 7564 1371
rect 7616 1368 7622 1420
rect 8386 1368 8392 1420
rect 8444 1408 8450 1420
rect 11256 1408 11284 1516
rect 11514 1436 11520 1488
rect 11572 1436 11578 1488
rect 11422 1417 11428 1420
rect 11420 1408 11428 1417
rect 8444 1380 11284 1408
rect 11383 1380 11428 1408
rect 8444 1368 8450 1380
rect 11420 1371 11428 1380
rect 11422 1368 11428 1371
rect 11480 1368 11486 1420
rect 11606 1368 11612 1420
rect 11664 1368 11670 1420
rect 11808 1417 11836 1516
rect 12066 1504 12072 1556
rect 12124 1504 12130 1556
rect 17954 1544 17960 1556
rect 12176 1516 17960 1544
rect 11793 1411 11851 1417
rect 11793 1377 11805 1411
rect 11839 1408 11851 1411
rect 12176 1408 12204 1516
rect 17954 1504 17960 1516
rect 18012 1504 18018 1556
rect 18046 1504 18052 1556
rect 18104 1544 18110 1556
rect 18141 1547 18199 1553
rect 18141 1544 18153 1547
rect 18104 1516 18153 1544
rect 18104 1504 18110 1516
rect 18141 1513 18153 1516
rect 18187 1513 18199 1547
rect 20346 1544 20352 1556
rect 18141 1507 18199 1513
rect 19168 1516 20352 1544
rect 12894 1436 12900 1488
rect 12952 1476 12958 1488
rect 13182 1479 13240 1485
rect 13182 1476 13194 1479
rect 12952 1448 13194 1476
rect 12952 1436 12958 1448
rect 13182 1445 13194 1448
rect 13228 1445 13240 1479
rect 15378 1476 15384 1488
rect 13182 1439 13240 1445
rect 14292 1448 15384 1476
rect 14292 1417 14320 1448
rect 15378 1436 15384 1448
rect 15436 1436 15442 1488
rect 17034 1485 17040 1488
rect 17028 1476 17040 1485
rect 16995 1448 17040 1476
rect 17028 1439 17040 1448
rect 17034 1436 17040 1439
rect 17092 1436 17098 1488
rect 18156 1476 18184 1507
rect 18601 1479 18659 1485
rect 18601 1476 18613 1479
rect 18156 1448 18613 1476
rect 18601 1445 18613 1448
rect 18647 1445 18659 1479
rect 18601 1439 18659 1445
rect 18693 1479 18751 1485
rect 18693 1445 18705 1479
rect 18739 1476 18751 1479
rect 19168 1476 19196 1516
rect 18739 1448 19196 1476
rect 18739 1445 18751 1448
rect 18693 1439 18751 1445
rect 14185 1411 14243 1417
rect 14185 1408 14197 1411
rect 11839 1380 12204 1408
rect 12406 1380 14197 1408
rect 11839 1377 11851 1380
rect 11793 1371 11851 1377
rect 5353 1343 5411 1349
rect 5353 1309 5365 1343
rect 5399 1340 5411 1343
rect 6730 1340 6736 1352
rect 5399 1312 6736 1340
rect 5399 1309 5411 1312
rect 5353 1303 5411 1309
rect 6730 1300 6736 1312
rect 6788 1300 6794 1352
rect 7285 1343 7343 1349
rect 7285 1309 7297 1343
rect 7331 1309 7343 1343
rect 7285 1303 7343 1309
rect 9309 1343 9367 1349
rect 9309 1309 9321 1343
rect 9355 1309 9367 1343
rect 11624 1340 11652 1368
rect 12406 1340 12434 1380
rect 11624 1312 12434 1340
rect 13449 1343 13507 1349
rect 9309 1303 9367 1309
rect 13449 1309 13461 1343
rect 13495 1309 13507 1343
rect 13449 1303 13507 1309
rect 6362 1232 6368 1284
rect 6420 1272 6426 1284
rect 7300 1272 7328 1303
rect 6420 1244 7328 1272
rect 6420 1232 6426 1244
rect 9324 1204 9352 1303
rect 9950 1204 9956 1216
rect 9324 1176 9956 1204
rect 9950 1164 9956 1176
rect 10008 1164 10014 1216
rect 11241 1207 11299 1213
rect 11241 1173 11253 1207
rect 11287 1204 11299 1207
rect 11330 1204 11336 1216
rect 11287 1176 11336 1204
rect 11287 1173 11299 1176
rect 11241 1167 11299 1173
rect 11330 1164 11336 1176
rect 11388 1164 11394 1216
rect 11882 1164 11888 1216
rect 11940 1204 11946 1216
rect 13464 1204 13492 1303
rect 14016 1272 14044 1380
rect 14185 1377 14197 1380
rect 14231 1377 14243 1411
rect 14185 1371 14243 1377
rect 14277 1411 14335 1417
rect 14277 1377 14289 1411
rect 14323 1377 14335 1411
rect 14277 1371 14335 1377
rect 14550 1368 14556 1420
rect 14608 1368 14614 1420
rect 15013 1411 15071 1417
rect 15013 1408 15025 1411
rect 14660 1380 15025 1408
rect 14090 1300 14096 1352
rect 14148 1340 14154 1352
rect 14369 1343 14427 1349
rect 14369 1340 14381 1343
rect 14148 1312 14381 1340
rect 14148 1300 14154 1312
rect 14369 1309 14381 1312
rect 14415 1340 14427 1343
rect 14458 1340 14464 1352
rect 14415 1312 14464 1340
rect 14415 1309 14427 1312
rect 14369 1303 14427 1309
rect 14458 1300 14464 1312
rect 14516 1300 14522 1352
rect 14660 1272 14688 1380
rect 15013 1377 15025 1380
rect 15059 1377 15071 1411
rect 15013 1371 15071 1377
rect 15105 1411 15163 1417
rect 15105 1377 15117 1411
rect 15151 1408 15163 1411
rect 15194 1408 15200 1420
rect 15151 1380 15200 1408
rect 15151 1377 15163 1380
rect 15105 1371 15163 1377
rect 15194 1368 15200 1380
rect 15252 1408 15258 1420
rect 15838 1408 15844 1420
rect 15252 1380 15844 1408
rect 15252 1368 15258 1380
rect 15838 1368 15844 1380
rect 15896 1368 15902 1420
rect 16298 1368 16304 1420
rect 16356 1408 16362 1420
rect 16356 1380 18368 1408
rect 16356 1368 16362 1380
rect 16758 1300 16764 1352
rect 16816 1300 16822 1352
rect 18340 1340 18368 1380
rect 18414 1368 18420 1420
rect 18472 1417 18478 1420
rect 18472 1411 18515 1417
rect 18503 1377 18515 1411
rect 18472 1371 18515 1377
rect 18472 1368 18478 1371
rect 18708 1340 18736 1439
rect 18874 1368 18880 1420
rect 18932 1368 18938 1420
rect 18966 1368 18972 1420
rect 19024 1368 19030 1420
rect 19168 1417 19196 1448
rect 19538 1479 19596 1485
rect 19538 1445 19550 1479
rect 19584 1476 19596 1479
rect 20070 1476 20076 1488
rect 19584 1448 20076 1476
rect 19584 1445 19596 1448
rect 19538 1439 19596 1445
rect 20070 1436 20076 1448
rect 20128 1436 20134 1488
rect 19153 1411 19211 1417
rect 19153 1377 19165 1411
rect 19199 1377 19211 1411
rect 19153 1371 19211 1377
rect 19242 1368 19248 1420
rect 19300 1368 19306 1420
rect 19342 1411 19400 1417
rect 19342 1377 19354 1411
rect 19388 1408 19400 1411
rect 19794 1408 19800 1420
rect 19388 1380 19800 1408
rect 19388 1377 19400 1380
rect 19342 1371 19400 1377
rect 19794 1368 19800 1380
rect 19852 1368 19858 1420
rect 19886 1368 19892 1420
rect 19944 1368 19950 1420
rect 20272 1417 20300 1516
rect 20346 1504 20352 1516
rect 20404 1504 20410 1556
rect 21542 1544 21548 1556
rect 20548 1516 21548 1544
rect 20257 1411 20315 1417
rect 20257 1377 20269 1411
rect 20303 1377 20315 1411
rect 20257 1371 20315 1377
rect 18340 1312 18736 1340
rect 20441 1343 20499 1349
rect 20441 1309 20453 1343
rect 20487 1340 20499 1343
rect 20548 1340 20576 1516
rect 21542 1504 21548 1516
rect 21600 1504 21606 1556
rect 21818 1504 21824 1556
rect 21876 1544 21882 1556
rect 22189 1547 22247 1553
rect 22189 1544 22201 1547
rect 21876 1516 22201 1544
rect 21876 1504 21882 1516
rect 22189 1513 22201 1516
rect 22235 1513 22247 1547
rect 22189 1507 22247 1513
rect 20901 1479 20959 1485
rect 20901 1445 20913 1479
rect 20947 1476 20959 1479
rect 25314 1476 25320 1488
rect 20947 1448 25320 1476
rect 20947 1445 20959 1448
rect 20901 1439 20959 1445
rect 25314 1436 25320 1448
rect 25372 1436 25378 1488
rect 21450 1368 21456 1420
rect 21508 1368 21514 1420
rect 21726 1368 21732 1420
rect 21784 1408 21790 1420
rect 21821 1411 21879 1417
rect 21821 1408 21833 1411
rect 21784 1380 21833 1408
rect 21784 1368 21790 1380
rect 21821 1377 21833 1380
rect 21867 1377 21879 1411
rect 21821 1371 21879 1377
rect 22002 1368 22008 1420
rect 22060 1408 22066 1420
rect 22922 1408 22928 1420
rect 22060 1380 22928 1408
rect 22060 1368 22066 1380
rect 22922 1368 22928 1380
rect 22980 1368 22986 1420
rect 20487 1312 20576 1340
rect 21545 1343 21603 1349
rect 20487 1309 20499 1312
rect 20441 1303 20499 1309
rect 21545 1309 21557 1343
rect 21591 1309 21603 1343
rect 21545 1303 21603 1309
rect 14016 1244 14688 1272
rect 19794 1232 19800 1284
rect 19852 1272 19858 1284
rect 21560 1272 21588 1303
rect 19852 1244 21588 1272
rect 19852 1232 19858 1244
rect 11940 1176 13492 1204
rect 11940 1164 11946 1176
rect 14826 1164 14832 1216
rect 14884 1204 14890 1216
rect 15565 1207 15623 1213
rect 15565 1204 15577 1207
rect 14884 1176 15577 1204
rect 14884 1164 14890 1176
rect 15565 1173 15577 1176
rect 15611 1173 15623 1207
rect 15565 1167 15623 1173
rect 18322 1164 18328 1216
rect 18380 1164 18386 1216
rect 552 1114 27416 1136
rect 552 1062 3756 1114
rect 3808 1062 3820 1114
rect 3872 1062 3884 1114
rect 3936 1062 3948 1114
rect 4000 1062 4012 1114
rect 4064 1062 10472 1114
rect 10524 1062 10536 1114
rect 10588 1062 10600 1114
rect 10652 1062 10664 1114
rect 10716 1062 10728 1114
rect 10780 1062 17188 1114
rect 17240 1062 17252 1114
rect 17304 1062 17316 1114
rect 17368 1062 17380 1114
rect 17432 1062 17444 1114
rect 17496 1062 23904 1114
rect 23956 1062 23968 1114
rect 24020 1062 24032 1114
rect 24084 1062 24096 1114
rect 24148 1062 24160 1114
rect 24212 1062 27416 1114
rect 552 1040 27416 1062
rect 11422 960 11428 1012
rect 11480 1000 11486 1012
rect 12986 1000 12992 1012
rect 11480 972 12992 1000
rect 11480 960 11486 972
rect 12986 960 12992 972
rect 13044 960 13050 1012
rect 14090 960 14096 1012
rect 14148 960 14154 1012
rect 14384 972 19656 1000
rect 5905 935 5963 941
rect 5905 901 5917 935
rect 5951 932 5963 935
rect 6086 932 6092 944
rect 5951 904 6092 932
rect 5951 901 5963 904
rect 5905 895 5963 901
rect 6086 892 6092 904
rect 6144 892 6150 944
rect 7834 892 7840 944
rect 7892 932 7898 944
rect 8021 935 8079 941
rect 8021 932 8033 935
rect 7892 904 8033 932
rect 7892 892 7898 904
rect 8021 901 8033 904
rect 8067 901 8079 935
rect 8021 895 8079 901
rect 9582 892 9588 944
rect 9640 892 9646 944
rect 13078 892 13084 944
rect 13136 892 13142 944
rect 6730 864 6736 876
rect 6104 836 6736 864
rect 6104 805 6132 836
rect 6730 824 6736 836
rect 6788 864 6794 876
rect 14384 864 14412 972
rect 19628 944 19656 972
rect 16574 892 16580 944
rect 16632 932 16638 944
rect 16669 935 16727 941
rect 16669 932 16681 935
rect 16632 904 16681 932
rect 16632 892 16638 904
rect 16669 901 16681 904
rect 16715 901 16727 935
rect 16669 895 16727 901
rect 19610 892 19616 944
rect 19668 932 19674 944
rect 19668 904 20208 932
rect 19668 892 19674 904
rect 6788 836 7604 864
rect 6788 824 6794 836
rect 6084 799 6142 805
rect 6084 765 6096 799
rect 6130 765 6142 799
rect 6084 759 6142 765
rect 6178 756 6184 808
rect 6236 756 6242 808
rect 6273 799 6331 805
rect 6273 765 6285 799
rect 6319 796 6331 799
rect 6362 796 6368 808
rect 6319 768 6368 796
rect 6319 765 6331 768
rect 6273 759 6331 765
rect 6362 756 6368 768
rect 6420 756 6426 808
rect 6457 799 6515 805
rect 6457 765 6469 799
rect 6503 796 6515 799
rect 6546 796 6552 808
rect 6503 768 6552 796
rect 6503 765 6515 768
rect 6457 759 6515 765
rect 6546 756 6552 768
rect 6604 756 6610 808
rect 7466 756 7472 808
rect 7524 756 7530 808
rect 7576 796 7604 836
rect 12544 836 14412 864
rect 15473 867 15531 873
rect 7889 799 7947 805
rect 7889 796 7901 799
rect 7576 768 7901 796
rect 7889 765 7901 768
rect 7935 796 7947 799
rect 7935 768 8524 796
rect 7935 765 7947 768
rect 7889 759 7947 765
rect 6380 728 6408 756
rect 7653 731 7711 737
rect 7653 728 7665 731
rect 6380 700 7665 728
rect 7653 697 7665 700
rect 7699 697 7711 731
rect 7653 691 7711 697
rect 7745 731 7803 737
rect 7745 697 7757 731
rect 7791 728 7803 731
rect 8294 728 8300 740
rect 7791 700 8300 728
rect 7791 697 7803 700
rect 7745 691 7803 697
rect 7668 660 7696 691
rect 8294 688 8300 700
rect 8352 688 8358 740
rect 8496 728 8524 768
rect 9030 756 9036 808
rect 9088 756 9094 808
rect 9453 799 9511 805
rect 9453 796 9465 799
rect 9140 768 9465 796
rect 9140 728 9168 768
rect 9453 765 9465 768
rect 9499 796 9511 799
rect 11422 796 11428 808
rect 9499 768 11428 796
rect 9499 765 9511 768
rect 9453 759 9511 765
rect 11422 756 11428 768
rect 11480 756 11486 808
rect 11974 756 11980 808
rect 12032 796 12038 808
rect 12544 805 12572 836
rect 15473 833 15485 867
rect 15519 864 15531 867
rect 16758 864 16764 876
rect 15519 836 16764 864
rect 15519 833 15531 836
rect 15473 827 15531 833
rect 16758 824 16764 836
rect 16816 824 16822 876
rect 19702 824 19708 876
rect 19760 864 19766 876
rect 20180 873 20208 904
rect 20165 867 20223 873
rect 19760 836 19932 864
rect 19760 824 19766 836
rect 12529 799 12587 805
rect 12529 796 12541 799
rect 12032 768 12541 796
rect 12032 756 12038 768
rect 12529 765 12541 768
rect 12575 765 12587 799
rect 12529 759 12587 765
rect 12802 756 12808 808
rect 12860 756 12866 808
rect 12986 805 12992 808
rect 12949 799 12992 805
rect 12949 765 12961 799
rect 12949 759 12992 765
rect 12986 756 12992 759
rect 13044 756 13050 808
rect 15217 799 15275 805
rect 15217 765 15229 799
rect 15263 796 15275 799
rect 15654 796 15660 808
rect 15263 768 15660 796
rect 15263 765 15275 768
rect 15217 759 15275 765
rect 15654 756 15660 768
rect 15712 756 15718 808
rect 16114 756 16120 808
rect 16172 756 16178 808
rect 16298 756 16304 808
rect 16356 756 16362 808
rect 16390 756 16396 808
rect 16448 756 16454 808
rect 16482 756 16488 808
rect 16540 805 16546 808
rect 16540 759 16548 805
rect 16540 756 16546 759
rect 19794 756 19800 808
rect 19852 756 19858 808
rect 19904 805 19932 836
rect 20165 833 20177 867
rect 20211 833 20223 867
rect 20165 827 20223 833
rect 19889 799 19947 805
rect 19889 765 19901 799
rect 19935 765 19947 799
rect 19889 759 19947 765
rect 20257 799 20315 805
rect 20257 765 20269 799
rect 20303 796 20315 799
rect 20346 796 20352 808
rect 20303 768 20352 796
rect 20303 765 20315 768
rect 20257 759 20315 765
rect 20346 756 20352 768
rect 20404 756 20410 808
rect 8496 700 9168 728
rect 9217 731 9275 737
rect 9217 697 9229 731
rect 9263 697 9275 731
rect 9217 691 9275 697
rect 9309 731 9367 737
rect 9309 697 9321 731
rect 9355 728 9367 731
rect 9858 728 9864 740
rect 9355 700 9864 728
rect 9355 697 9367 700
rect 9309 691 9367 697
rect 9232 660 9260 691
rect 9858 688 9864 700
rect 9916 688 9922 740
rect 12713 731 12771 737
rect 12713 697 12725 731
rect 12759 697 12771 731
rect 12713 691 12771 697
rect 20901 731 20959 737
rect 20901 697 20913 731
rect 20947 728 20959 731
rect 27062 728 27068 740
rect 20947 700 27068 728
rect 20947 697 20959 700
rect 20901 691 20959 697
rect 11606 660 11612 672
rect 7668 632 11612 660
rect 11606 620 11612 632
rect 11664 660 11670 672
rect 12728 660 12756 691
rect 27062 688 27068 700
rect 27120 688 27126 740
rect 11664 632 12756 660
rect 11664 620 11670 632
rect 552 570 27576 592
rect 552 518 7114 570
rect 7166 518 7178 570
rect 7230 518 7242 570
rect 7294 518 7306 570
rect 7358 518 7370 570
rect 7422 518 13830 570
rect 13882 518 13894 570
rect 13946 518 13958 570
rect 14010 518 14022 570
rect 14074 518 14086 570
rect 14138 518 20546 570
rect 20598 518 20610 570
rect 20662 518 20674 570
rect 20726 518 20738 570
rect 20790 518 20802 570
rect 20854 518 27262 570
rect 27314 518 27326 570
rect 27378 518 27390 570
rect 27442 518 27454 570
rect 27506 518 27518 570
rect 27570 518 27576 570
rect 552 496 27576 518
<< via1 >>
rect 10232 17552 10284 17604
rect 10416 17552 10468 17604
rect 16764 17552 16816 17604
rect 25136 17552 25188 17604
rect 3608 17484 3660 17536
rect 3976 17484 4028 17536
rect 18972 17484 19024 17536
rect 24676 17484 24728 17536
rect 3756 17382 3808 17434
rect 3820 17382 3872 17434
rect 3884 17382 3936 17434
rect 3948 17382 4000 17434
rect 4012 17382 4064 17434
rect 10472 17382 10524 17434
rect 10536 17382 10588 17434
rect 10600 17382 10652 17434
rect 10664 17382 10716 17434
rect 10728 17382 10780 17434
rect 17188 17382 17240 17434
rect 17252 17382 17304 17434
rect 17316 17382 17368 17434
rect 17380 17382 17432 17434
rect 17444 17382 17496 17434
rect 23904 17382 23956 17434
rect 23968 17382 24020 17434
rect 24032 17382 24084 17434
rect 24096 17382 24148 17434
rect 24160 17382 24212 17434
rect 848 17323 900 17332
rect 848 17289 857 17323
rect 857 17289 891 17323
rect 891 17289 900 17323
rect 848 17280 900 17289
rect 1492 17323 1544 17332
rect 1492 17289 1501 17323
rect 1501 17289 1535 17323
rect 1535 17289 1544 17323
rect 1492 17280 1544 17289
rect 3608 17280 3660 17332
rect 5908 17280 5960 17332
rect 6552 17280 6604 17332
rect 8484 17280 8536 17332
rect 9128 17280 9180 17332
rect 10232 17280 10284 17332
rect 11704 17280 11756 17332
rect 13636 17280 13688 17332
rect 20352 17280 20404 17332
rect 24676 17323 24728 17332
rect 24676 17289 24685 17323
rect 24685 17289 24719 17323
rect 24719 17289 24728 17323
rect 24676 17280 24728 17289
rect 25136 17323 25188 17332
rect 25136 17289 25145 17323
rect 25145 17289 25179 17323
rect 25179 17289 25188 17323
rect 25136 17280 25188 17289
rect 12164 17212 12216 17264
rect 19064 17212 19116 17264
rect 2688 17144 2740 17196
rect 3424 17187 3476 17196
rect 3424 17153 3433 17187
rect 3433 17153 3467 17187
rect 3467 17153 3476 17187
rect 3424 17144 3476 17153
rect 4712 17187 4764 17196
rect 4712 17153 4721 17187
rect 4721 17153 4755 17187
rect 4755 17153 4764 17187
rect 4712 17144 4764 17153
rect 5264 17144 5316 17196
rect 7840 17076 7892 17128
rect 9956 17076 10008 17128
rect 10784 17119 10836 17128
rect 10784 17085 10793 17119
rect 10793 17085 10827 17119
rect 10827 17085 10836 17119
rect 10784 17076 10836 17085
rect 11888 17119 11940 17128
rect 11888 17085 11897 17119
rect 11897 17085 11931 17119
rect 11931 17085 11940 17119
rect 11888 17076 11940 17085
rect 14556 17076 14608 17128
rect 16488 17119 16540 17128
rect 16488 17085 16497 17119
rect 16497 17085 16531 17119
rect 16531 17085 16540 17119
rect 16488 17076 16540 17085
rect 16856 17076 16908 17128
rect 17776 17119 17828 17128
rect 17776 17085 17785 17119
rect 17785 17085 17819 17119
rect 17819 17085 17828 17119
rect 17776 17076 17828 17085
rect 19432 17144 19484 17196
rect 19984 17144 20036 17196
rect 20168 17144 20220 17196
rect 20720 17212 20772 17264
rect 18972 17119 19024 17128
rect 18972 17085 18981 17119
rect 18981 17085 19015 17119
rect 19015 17085 19024 17119
rect 18972 17076 19024 17085
rect 19064 17119 19116 17128
rect 19064 17085 19073 17119
rect 19073 17085 19107 17119
rect 19107 17085 19116 17119
rect 19064 17076 19116 17085
rect 19524 17119 19576 17128
rect 19524 17085 19533 17119
rect 19533 17085 19567 17119
rect 19567 17085 19576 17119
rect 19524 17076 19576 17085
rect 20352 17076 20404 17128
rect 20720 17119 20772 17128
rect 20720 17085 20729 17119
rect 20729 17085 20763 17119
rect 20763 17085 20772 17119
rect 24032 17255 24084 17264
rect 24032 17221 24041 17255
rect 24041 17221 24075 17255
rect 24075 17221 24084 17255
rect 24032 17212 24084 17221
rect 20720 17076 20772 17085
rect 21364 17076 21416 17128
rect 25872 17144 25924 17196
rect 9404 16940 9456 16992
rect 15108 16940 15160 16992
rect 17592 16983 17644 16992
rect 17592 16949 17601 16983
rect 17601 16949 17635 16983
rect 17635 16949 17644 16983
rect 17592 16940 17644 16949
rect 17776 16940 17828 16992
rect 18420 16940 18472 16992
rect 19340 16983 19392 16992
rect 19340 16949 19349 16983
rect 19349 16949 19383 16983
rect 19383 16949 19392 16983
rect 19340 16940 19392 16949
rect 19892 16983 19944 16992
rect 19892 16949 19901 16983
rect 19901 16949 19935 16983
rect 19935 16949 19944 16983
rect 19892 16940 19944 16949
rect 19984 16940 20036 16992
rect 21456 16940 21508 16992
rect 22284 17076 22336 17128
rect 22652 17076 22704 17128
rect 23296 17076 23348 17128
rect 23756 17076 23808 17128
rect 24584 17076 24636 17128
rect 25228 17076 25280 17128
rect 25504 17076 25556 17128
rect 26332 17076 26384 17128
rect 24124 17008 24176 17060
rect 24676 17008 24728 17060
rect 26976 17008 27028 17060
rect 23112 16940 23164 16992
rect 26700 16940 26752 16992
rect 7114 16838 7166 16890
rect 7178 16838 7230 16890
rect 7242 16838 7294 16890
rect 7306 16838 7358 16890
rect 7370 16838 7422 16890
rect 13830 16838 13882 16890
rect 13894 16838 13946 16890
rect 13958 16838 14010 16890
rect 14022 16838 14074 16890
rect 14086 16838 14138 16890
rect 20546 16838 20598 16890
rect 20610 16838 20662 16890
rect 20674 16838 20726 16890
rect 20738 16838 20790 16890
rect 20802 16838 20854 16890
rect 27262 16838 27314 16890
rect 27326 16838 27378 16890
rect 27390 16838 27442 16890
rect 27454 16838 27506 16890
rect 27518 16838 27570 16890
rect 9680 16736 9732 16788
rect 9772 16779 9824 16788
rect 9772 16745 9781 16779
rect 9781 16745 9815 16779
rect 9815 16745 9824 16779
rect 9772 16736 9824 16745
rect 10784 16736 10836 16788
rect 12992 16736 13044 16788
rect 12716 16668 12768 16720
rect 14280 16736 14332 16788
rect 15844 16779 15896 16788
rect 15844 16745 15853 16779
rect 15853 16745 15887 16779
rect 15887 16745 15896 16779
rect 15844 16736 15896 16745
rect 19800 16736 19852 16788
rect 17592 16668 17644 16720
rect 20720 16668 20772 16720
rect 24124 16736 24176 16788
rect 25964 16736 26016 16788
rect 8484 16643 8536 16652
rect 8484 16609 8518 16643
rect 8518 16609 8536 16643
rect 8484 16600 8536 16609
rect 9956 16643 10008 16652
rect 5816 16532 5868 16584
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 10784 16643 10836 16652
rect 10784 16609 10793 16643
rect 10793 16609 10827 16643
rect 10827 16609 10836 16643
rect 10784 16600 10836 16609
rect 11152 16600 11204 16652
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 12992 16643 13044 16652
rect 12992 16609 13001 16643
rect 13001 16609 13035 16643
rect 13035 16609 13044 16643
rect 12992 16600 13044 16609
rect 14004 16643 14056 16652
rect 14004 16609 14013 16643
rect 14013 16609 14047 16643
rect 14047 16609 14056 16643
rect 14004 16600 14056 16609
rect 14280 16600 14332 16652
rect 15200 16600 15252 16652
rect 15568 16600 15620 16652
rect 16580 16643 16632 16652
rect 16580 16609 16589 16643
rect 16589 16609 16623 16643
rect 16623 16609 16632 16643
rect 16580 16600 16632 16609
rect 16764 16643 16816 16652
rect 16764 16609 16773 16643
rect 16773 16609 16807 16643
rect 16807 16609 16816 16643
rect 16764 16600 16816 16609
rect 14832 16532 14884 16584
rect 15108 16575 15160 16584
rect 15108 16541 15117 16575
rect 15117 16541 15151 16575
rect 15151 16541 15160 16575
rect 15108 16532 15160 16541
rect 19064 16600 19116 16652
rect 18512 16575 18564 16584
rect 18512 16541 18521 16575
rect 18521 16541 18555 16575
rect 18555 16541 18564 16575
rect 18512 16532 18564 16541
rect 19616 16643 19668 16652
rect 19616 16609 19625 16643
rect 19625 16609 19659 16643
rect 19659 16609 19668 16643
rect 19616 16600 19668 16609
rect 19800 16600 19852 16652
rect 20904 16532 20956 16584
rect 22652 16643 22704 16652
rect 22652 16609 22661 16643
rect 22661 16609 22695 16643
rect 22695 16609 22704 16643
rect 22652 16600 22704 16609
rect 7840 16439 7892 16448
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 10140 16439 10192 16448
rect 10140 16405 10149 16439
rect 10149 16405 10183 16439
rect 10183 16405 10192 16439
rect 10140 16396 10192 16405
rect 13360 16396 13412 16448
rect 19064 16439 19116 16448
rect 19064 16405 19073 16439
rect 19073 16405 19107 16439
rect 19107 16405 19116 16439
rect 19064 16396 19116 16405
rect 19616 16396 19668 16448
rect 21364 16396 21416 16448
rect 22100 16464 22152 16516
rect 24124 16643 24176 16652
rect 24124 16609 24133 16643
rect 24133 16609 24167 16643
rect 24167 16609 24176 16643
rect 24124 16600 24176 16609
rect 24308 16643 24360 16652
rect 24308 16609 24317 16643
rect 24317 16609 24351 16643
rect 24351 16609 24360 16643
rect 24308 16600 24360 16609
rect 25320 16600 25372 16652
rect 25596 16668 25648 16720
rect 26240 16643 26292 16652
rect 26240 16609 26249 16643
rect 26249 16609 26283 16643
rect 26283 16609 26292 16643
rect 26240 16600 26292 16609
rect 26700 16643 26752 16652
rect 26700 16609 26709 16643
rect 26709 16609 26743 16643
rect 26743 16609 26752 16643
rect 26700 16600 26752 16609
rect 26884 16643 26936 16652
rect 26884 16609 26893 16643
rect 26893 16609 26927 16643
rect 26927 16609 26936 16643
rect 26884 16600 26936 16609
rect 26976 16600 27028 16652
rect 23480 16575 23532 16584
rect 23480 16541 23489 16575
rect 23489 16541 23523 16575
rect 23523 16541 23532 16575
rect 23480 16532 23532 16541
rect 24952 16439 25004 16448
rect 24952 16405 24961 16439
rect 24961 16405 24995 16439
rect 24995 16405 25004 16439
rect 24952 16396 25004 16405
rect 25688 16396 25740 16448
rect 3756 16294 3808 16346
rect 3820 16294 3872 16346
rect 3884 16294 3936 16346
rect 3948 16294 4000 16346
rect 4012 16294 4064 16346
rect 10472 16294 10524 16346
rect 10536 16294 10588 16346
rect 10600 16294 10652 16346
rect 10664 16294 10716 16346
rect 10728 16294 10780 16346
rect 17188 16294 17240 16346
rect 17252 16294 17304 16346
rect 17316 16294 17368 16346
rect 17380 16294 17432 16346
rect 17444 16294 17496 16346
rect 23904 16294 23956 16346
rect 23968 16294 24020 16346
rect 24032 16294 24084 16346
rect 24096 16294 24148 16346
rect 24160 16294 24212 16346
rect 7472 16192 7524 16244
rect 8484 16235 8536 16244
rect 8484 16201 8493 16235
rect 8493 16201 8527 16235
rect 8527 16201 8536 16235
rect 8484 16192 8536 16201
rect 9680 16192 9732 16244
rect 10324 16235 10376 16244
rect 10324 16201 10333 16235
rect 10333 16201 10367 16235
rect 10367 16201 10376 16235
rect 10324 16192 10376 16201
rect 11060 16192 11112 16244
rect 12256 16192 12308 16244
rect 14924 16192 14976 16244
rect 22652 16192 22704 16244
rect 6460 16167 6512 16176
rect 6460 16133 6469 16167
rect 6469 16133 6503 16167
rect 6503 16133 6512 16167
rect 6460 16124 6512 16133
rect 7564 15988 7616 16040
rect 8760 16031 8812 16040
rect 8760 15997 8769 16031
rect 8769 15997 8803 16031
rect 8803 15997 8812 16031
rect 8760 15988 8812 15997
rect 8852 16031 8904 16040
rect 8852 15997 8861 16031
rect 8861 15997 8895 16031
rect 8895 15997 8904 16031
rect 8852 15988 8904 15997
rect 6736 15920 6788 15972
rect 7656 15963 7708 15972
rect 7656 15929 7665 15963
rect 7665 15929 7699 15963
rect 7699 15929 7708 15963
rect 7656 15920 7708 15929
rect 7840 15963 7892 15972
rect 7840 15929 7849 15963
rect 7849 15929 7883 15963
rect 7883 15929 7892 15963
rect 7840 15920 7892 15929
rect 8668 15920 8720 15972
rect 9404 16031 9456 16040
rect 9404 15997 9413 16031
rect 9413 15997 9447 16031
rect 9447 15997 9456 16031
rect 9404 15988 9456 15997
rect 9680 16031 9732 16040
rect 9680 15997 9689 16031
rect 9689 15997 9723 16031
rect 9723 15997 9732 16031
rect 9680 15988 9732 15997
rect 23480 16124 23532 16176
rect 10140 15988 10192 16040
rect 10876 16031 10928 16040
rect 10876 15997 10885 16031
rect 10885 15997 10919 16031
rect 10919 15997 10928 16031
rect 10876 15988 10928 15997
rect 11060 15988 11112 16040
rect 11244 16056 11296 16108
rect 11152 15963 11204 15972
rect 11152 15929 11161 15963
rect 11161 15929 11195 15963
rect 11195 15929 11204 15963
rect 11152 15920 11204 15929
rect 7472 15852 7524 15904
rect 9680 15852 9732 15904
rect 10140 15852 10192 15904
rect 10968 15852 11020 15904
rect 11520 15988 11572 16040
rect 20720 16099 20772 16108
rect 20720 16065 20729 16099
rect 20729 16065 20763 16099
rect 20763 16065 20772 16099
rect 20720 16056 20772 16065
rect 22928 16056 22980 16108
rect 25320 16235 25372 16244
rect 25320 16201 25329 16235
rect 25329 16201 25363 16235
rect 25363 16201 25372 16235
rect 25320 16192 25372 16201
rect 25688 16124 25740 16176
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 12624 15988 12676 16040
rect 13360 16031 13412 16040
rect 13360 15997 13369 16031
rect 13369 15997 13403 16031
rect 13403 15997 13412 16031
rect 13360 15988 13412 15997
rect 14280 15988 14332 16040
rect 14648 16031 14700 16040
rect 14648 15997 14657 16031
rect 14657 15997 14691 16031
rect 14691 15997 14700 16031
rect 14648 15988 14700 15997
rect 14740 15988 14792 16040
rect 15108 16031 15160 16040
rect 15108 15997 15117 16031
rect 15117 15997 15151 16031
rect 15151 15997 15160 16031
rect 15108 15988 15160 15997
rect 17040 15988 17092 16040
rect 18328 15988 18380 16040
rect 21088 16031 21140 16040
rect 21088 15997 21097 16031
rect 21097 15997 21131 16031
rect 21131 15997 21140 16031
rect 21088 15988 21140 15997
rect 21364 16031 21416 16040
rect 21364 15997 21398 16031
rect 21398 15997 21416 16031
rect 21364 15988 21416 15997
rect 22284 15988 22336 16040
rect 11796 15920 11848 15972
rect 24584 15988 24636 16040
rect 11704 15852 11756 15904
rect 13084 15895 13136 15904
rect 13084 15861 13093 15895
rect 13093 15861 13127 15895
rect 13127 15861 13136 15895
rect 13084 15852 13136 15861
rect 14924 15852 14976 15904
rect 18880 15852 18932 15904
rect 20904 15852 20956 15904
rect 22836 15852 22888 15904
rect 23296 15852 23348 15904
rect 24860 15920 24912 15972
rect 24952 15963 25004 15972
rect 24952 15929 24970 15963
rect 24970 15929 25004 15963
rect 24952 15920 25004 15929
rect 26240 16031 26292 16040
rect 26240 15997 26249 16031
rect 26249 15997 26283 16031
rect 26283 15997 26292 16031
rect 26240 15988 26292 15997
rect 26608 15852 26660 15904
rect 7114 15750 7166 15802
rect 7178 15750 7230 15802
rect 7242 15750 7294 15802
rect 7306 15750 7358 15802
rect 7370 15750 7422 15802
rect 13830 15750 13882 15802
rect 13894 15750 13946 15802
rect 13958 15750 14010 15802
rect 14022 15750 14074 15802
rect 14086 15750 14138 15802
rect 20546 15750 20598 15802
rect 20610 15750 20662 15802
rect 20674 15750 20726 15802
rect 20738 15750 20790 15802
rect 20802 15750 20854 15802
rect 27262 15750 27314 15802
rect 27326 15750 27378 15802
rect 27390 15750 27442 15802
rect 27454 15750 27506 15802
rect 27518 15750 27570 15802
rect 4620 15512 4672 15564
rect 8668 15648 8720 15700
rect 8760 15691 8812 15700
rect 8760 15657 8769 15691
rect 8769 15657 8803 15691
rect 8803 15657 8812 15691
rect 8760 15648 8812 15657
rect 8852 15648 8904 15700
rect 11612 15648 11664 15700
rect 12440 15648 12492 15700
rect 18512 15648 18564 15700
rect 22100 15691 22152 15700
rect 22100 15657 22109 15691
rect 22109 15657 22143 15691
rect 22143 15657 22152 15691
rect 22100 15648 22152 15657
rect 23296 15648 23348 15700
rect 26884 15648 26936 15700
rect 7472 15580 7524 15632
rect 7656 15580 7708 15632
rect 5816 15555 5868 15564
rect 5816 15521 5825 15555
rect 5825 15521 5859 15555
rect 5859 15521 5868 15555
rect 5816 15512 5868 15521
rect 6368 15512 6420 15564
rect 8208 15512 8260 15564
rect 9680 15580 9732 15632
rect 5172 15351 5224 15360
rect 5172 15317 5181 15351
rect 5181 15317 5215 15351
rect 5215 15317 5224 15351
rect 5172 15308 5224 15317
rect 9864 15444 9916 15496
rect 10968 15555 11020 15564
rect 10968 15521 10977 15555
rect 10977 15521 11011 15555
rect 11011 15521 11020 15555
rect 10968 15512 11020 15521
rect 11336 15512 11388 15564
rect 12624 15580 12676 15632
rect 13084 15580 13136 15632
rect 11796 15555 11848 15564
rect 11796 15521 11805 15555
rect 11805 15521 11839 15555
rect 11839 15521 11848 15555
rect 11796 15512 11848 15521
rect 12348 15512 12400 15564
rect 16672 15512 16724 15564
rect 18328 15580 18380 15632
rect 22468 15623 22520 15632
rect 22468 15589 22477 15623
rect 22477 15589 22511 15623
rect 22511 15589 22520 15623
rect 22468 15580 22520 15589
rect 6920 15376 6972 15428
rect 10048 15376 10100 15428
rect 10968 15376 11020 15428
rect 11796 15376 11848 15428
rect 15476 15444 15528 15496
rect 14280 15376 14332 15428
rect 7012 15308 7064 15360
rect 8668 15308 8720 15360
rect 11152 15308 11204 15360
rect 11428 15351 11480 15360
rect 11428 15317 11437 15351
rect 11437 15317 11471 15351
rect 11471 15317 11480 15351
rect 11428 15308 11480 15317
rect 14464 15308 14516 15360
rect 19064 15555 19116 15564
rect 19064 15521 19073 15555
rect 19073 15521 19107 15555
rect 19107 15521 19116 15555
rect 19064 15512 19116 15521
rect 19616 15512 19668 15564
rect 21272 15512 21324 15564
rect 22284 15512 22336 15564
rect 23480 15580 23532 15632
rect 25596 15580 25648 15632
rect 19156 15444 19208 15496
rect 20076 15444 20128 15496
rect 21364 15487 21416 15496
rect 21364 15453 21373 15487
rect 21373 15453 21407 15487
rect 21407 15453 21416 15487
rect 22744 15555 22796 15564
rect 22744 15521 22753 15555
rect 22753 15521 22787 15555
rect 22787 15521 22796 15555
rect 22744 15512 22796 15521
rect 21364 15444 21416 15453
rect 19892 15376 19944 15428
rect 23020 15555 23072 15564
rect 23020 15521 23029 15555
rect 23029 15521 23063 15555
rect 23063 15521 23072 15555
rect 23020 15512 23072 15521
rect 22928 15444 22980 15496
rect 26424 15555 26476 15564
rect 26424 15521 26433 15555
rect 26433 15521 26467 15555
rect 26467 15521 26476 15555
rect 26424 15512 26476 15521
rect 26608 15555 26660 15564
rect 26608 15521 26615 15555
rect 26615 15521 26660 15555
rect 26608 15512 26660 15521
rect 26700 15555 26752 15564
rect 26700 15521 26709 15555
rect 26709 15521 26743 15555
rect 26743 15521 26752 15555
rect 26700 15512 26752 15521
rect 26792 15555 26844 15564
rect 26792 15521 26801 15555
rect 26801 15521 26835 15555
rect 26835 15521 26844 15555
rect 26792 15512 26844 15521
rect 26884 15555 26936 15564
rect 26884 15521 26898 15555
rect 26898 15521 26932 15555
rect 26932 15521 26936 15555
rect 26884 15512 26936 15521
rect 24768 15444 24820 15496
rect 24860 15487 24912 15496
rect 24860 15453 24869 15487
rect 24869 15453 24903 15487
rect 24903 15453 24912 15487
rect 24860 15444 24912 15453
rect 23572 15376 23624 15428
rect 19248 15308 19300 15360
rect 20720 15308 20772 15360
rect 22100 15308 22152 15360
rect 23480 15351 23532 15360
rect 23480 15317 23489 15351
rect 23489 15317 23523 15351
rect 23523 15317 23532 15351
rect 23480 15308 23532 15317
rect 26332 15308 26384 15360
rect 3756 15206 3808 15258
rect 3820 15206 3872 15258
rect 3884 15206 3936 15258
rect 3948 15206 4000 15258
rect 4012 15206 4064 15258
rect 10472 15206 10524 15258
rect 10536 15206 10588 15258
rect 10600 15206 10652 15258
rect 10664 15206 10716 15258
rect 10728 15206 10780 15258
rect 17188 15206 17240 15258
rect 17252 15206 17304 15258
rect 17316 15206 17368 15258
rect 17380 15206 17432 15258
rect 17444 15206 17496 15258
rect 23904 15206 23956 15258
rect 23968 15206 24020 15258
rect 24032 15206 24084 15258
rect 24096 15206 24148 15258
rect 24160 15206 24212 15258
rect 6460 15147 6512 15156
rect 6460 15113 6469 15147
rect 6469 15113 6503 15147
rect 6503 15113 6512 15147
rect 6460 15104 6512 15113
rect 7472 15147 7524 15156
rect 7472 15113 7481 15147
rect 7481 15113 7515 15147
rect 7515 15113 7524 15147
rect 7472 15104 7524 15113
rect 9956 15104 10008 15156
rect 3608 14968 3660 15020
rect 10232 15036 10284 15088
rect 11060 15104 11112 15156
rect 11336 15104 11388 15156
rect 13360 15104 13412 15156
rect 15476 15147 15528 15156
rect 15476 15113 15485 15147
rect 15485 15113 15519 15147
rect 15519 15113 15528 15147
rect 15476 15104 15528 15113
rect 17040 15147 17092 15156
rect 17040 15113 17049 15147
rect 17049 15113 17083 15147
rect 17083 15113 17092 15147
rect 17040 15104 17092 15113
rect 10968 15036 11020 15088
rect 11152 15036 11204 15088
rect 2044 14832 2096 14884
rect 3792 14900 3844 14952
rect 4160 14900 4212 14952
rect 5816 14900 5868 14952
rect 6828 14900 6880 14952
rect 7012 14900 7064 14952
rect 8484 14900 8536 14952
rect 11428 14968 11480 15020
rect 9680 14900 9732 14952
rect 2320 14764 2372 14816
rect 5172 14832 5224 14884
rect 7656 14832 7708 14884
rect 9864 14875 9916 14884
rect 9864 14841 9873 14875
rect 9873 14841 9907 14875
rect 9907 14841 9916 14875
rect 9864 14832 9916 14841
rect 10048 14943 10100 14952
rect 10048 14909 10057 14943
rect 10057 14909 10091 14943
rect 10091 14909 10100 14943
rect 10048 14900 10100 14909
rect 11152 14900 11204 14952
rect 11704 14968 11756 15020
rect 11980 14943 12032 14952
rect 11980 14909 11989 14943
rect 11989 14909 12023 14943
rect 12023 14909 12032 14943
rect 11980 14900 12032 14909
rect 14188 14900 14240 14952
rect 16672 14900 16724 14952
rect 16948 14900 17000 14952
rect 19064 15104 19116 15156
rect 19892 15104 19944 15156
rect 18604 14900 18656 14952
rect 18880 14900 18932 14952
rect 19064 14943 19116 14952
rect 19064 14909 19073 14943
rect 19073 14909 19107 14943
rect 19107 14909 19116 14943
rect 19064 14900 19116 14909
rect 19800 14968 19852 15020
rect 20260 14968 20312 15020
rect 19248 14900 19300 14952
rect 20168 14900 20220 14952
rect 20352 14943 20404 14952
rect 20352 14909 20356 14943
rect 20356 14909 20390 14943
rect 20390 14909 20404 14943
rect 20352 14900 20404 14909
rect 20628 14900 20680 14952
rect 20904 14968 20956 15020
rect 22744 15104 22796 15156
rect 24492 15104 24544 15156
rect 24768 15104 24820 15156
rect 21088 14968 21140 15020
rect 23848 15011 23900 15020
rect 20996 14900 21048 14952
rect 21732 14900 21784 14952
rect 22744 14900 22796 14952
rect 23848 14977 23857 15011
rect 23857 14977 23891 15011
rect 23891 14977 23900 15011
rect 23848 14968 23900 14977
rect 23204 14943 23256 14952
rect 23204 14909 23213 14943
rect 23213 14909 23247 14943
rect 23247 14909 23256 14943
rect 23204 14900 23256 14909
rect 12348 14832 12400 14884
rect 14372 14875 14424 14884
rect 14372 14841 14406 14875
rect 14406 14841 14424 14875
rect 14372 14832 14424 14841
rect 6552 14807 6604 14816
rect 6552 14773 6561 14807
rect 6561 14773 6595 14807
rect 6595 14773 6604 14807
rect 6552 14764 6604 14773
rect 6644 14764 6696 14816
rect 9036 14764 9088 14816
rect 10048 14764 10100 14816
rect 10324 14764 10376 14816
rect 10600 14764 10652 14816
rect 11152 14764 11204 14816
rect 11336 14764 11388 14816
rect 13544 14764 13596 14816
rect 13728 14764 13780 14816
rect 16120 14764 16172 14816
rect 17868 14875 17920 14884
rect 17868 14841 17877 14875
rect 17877 14841 17911 14875
rect 17911 14841 17920 14875
rect 17868 14832 17920 14841
rect 18236 14832 18288 14884
rect 18788 14832 18840 14884
rect 19432 14807 19484 14816
rect 19432 14773 19441 14807
rect 19441 14773 19475 14807
rect 19475 14773 19484 14807
rect 19432 14764 19484 14773
rect 22284 14832 22336 14884
rect 22376 14832 22428 14884
rect 23480 14832 23532 14884
rect 24676 14832 24728 14884
rect 25872 14943 25924 14952
rect 25872 14909 25881 14943
rect 25881 14909 25915 14943
rect 25915 14909 25924 14943
rect 25872 14900 25924 14909
rect 25964 14943 26016 14952
rect 25964 14909 25973 14943
rect 25973 14909 26007 14943
rect 26007 14909 26016 14943
rect 25964 14900 26016 14909
rect 26608 14900 26660 14952
rect 25044 14832 25096 14884
rect 21180 14764 21232 14816
rect 22468 14764 22520 14816
rect 22836 14764 22888 14816
rect 23296 14764 23348 14816
rect 24400 14764 24452 14816
rect 26424 14807 26476 14816
rect 26424 14773 26433 14807
rect 26433 14773 26467 14807
rect 26467 14773 26476 14807
rect 26424 14764 26476 14773
rect 7114 14662 7166 14714
rect 7178 14662 7230 14714
rect 7242 14662 7294 14714
rect 7306 14662 7358 14714
rect 7370 14662 7422 14714
rect 13830 14662 13882 14714
rect 13894 14662 13946 14714
rect 13958 14662 14010 14714
rect 14022 14662 14074 14714
rect 14086 14662 14138 14714
rect 20546 14662 20598 14714
rect 20610 14662 20662 14714
rect 20674 14662 20726 14714
rect 20738 14662 20790 14714
rect 20802 14662 20854 14714
rect 27262 14662 27314 14714
rect 27326 14662 27378 14714
rect 27390 14662 27442 14714
rect 27454 14662 27506 14714
rect 27518 14662 27570 14714
rect 3792 14603 3844 14612
rect 3792 14569 3801 14603
rect 3801 14569 3835 14603
rect 3835 14569 3844 14603
rect 3792 14560 3844 14569
rect 6368 14603 6420 14612
rect 6368 14569 6377 14603
rect 6377 14569 6411 14603
rect 6411 14569 6420 14603
rect 6368 14560 6420 14569
rect 6460 14560 6512 14612
rect 2320 14467 2372 14476
rect 2320 14433 2329 14467
rect 2329 14433 2363 14467
rect 2363 14433 2372 14467
rect 2320 14424 2372 14433
rect 3240 14424 3292 14476
rect 6644 14492 6696 14544
rect 4252 14424 4304 14476
rect 6552 14467 6604 14476
rect 6552 14433 6561 14467
rect 6561 14433 6595 14467
rect 6595 14433 6604 14467
rect 6552 14424 6604 14433
rect 10600 14560 10652 14612
rect 10876 14560 10928 14612
rect 11612 14560 11664 14612
rect 14372 14560 14424 14612
rect 14464 14560 14516 14612
rect 8300 14492 8352 14544
rect 2412 14399 2464 14408
rect 2412 14365 2421 14399
rect 2421 14365 2455 14399
rect 2455 14365 2464 14399
rect 2412 14356 2464 14365
rect 3424 14356 3476 14408
rect 4620 14356 4672 14408
rect 4804 14356 4856 14408
rect 6644 14399 6696 14408
rect 6644 14365 6653 14399
rect 6653 14365 6687 14399
rect 6687 14365 6696 14399
rect 6644 14356 6696 14365
rect 7748 14424 7800 14476
rect 8484 14467 8536 14476
rect 8484 14433 8493 14467
rect 8493 14433 8527 14467
rect 8527 14433 8536 14467
rect 8484 14424 8536 14433
rect 1768 14220 1820 14272
rect 2228 14263 2280 14272
rect 2228 14229 2237 14263
rect 2237 14229 2271 14263
rect 2271 14229 2280 14263
rect 2228 14220 2280 14229
rect 3516 14288 3568 14340
rect 2688 14220 2740 14272
rect 3608 14220 3660 14272
rect 4620 14263 4672 14272
rect 4620 14229 4629 14263
rect 4629 14229 4663 14263
rect 4663 14229 4672 14263
rect 4620 14220 4672 14229
rect 5908 14288 5960 14340
rect 7012 14288 7064 14340
rect 9036 14467 9088 14476
rect 9036 14433 9045 14467
rect 9045 14433 9079 14467
rect 9079 14433 9088 14467
rect 9036 14424 9088 14433
rect 9588 14492 9640 14544
rect 9864 14492 9916 14544
rect 9404 14356 9456 14408
rect 10140 14465 10192 14474
rect 10140 14431 10149 14465
rect 10149 14431 10183 14465
rect 10183 14431 10192 14465
rect 10140 14422 10192 14431
rect 10416 14424 10468 14476
rect 10876 14424 10928 14476
rect 11152 14467 11204 14476
rect 11152 14433 11161 14467
rect 11161 14433 11195 14467
rect 11195 14433 11204 14467
rect 11152 14424 11204 14433
rect 11336 14467 11388 14476
rect 11336 14433 11345 14467
rect 11345 14433 11379 14467
rect 11379 14433 11388 14467
rect 11336 14424 11388 14433
rect 13084 14424 13136 14476
rect 13360 14467 13412 14476
rect 13360 14433 13369 14467
rect 13369 14433 13403 14467
rect 13403 14433 13412 14467
rect 13360 14424 13412 14433
rect 13544 14467 13596 14476
rect 13544 14433 13553 14467
rect 13553 14433 13587 14467
rect 13587 14433 13596 14467
rect 13544 14424 13596 14433
rect 16396 14560 16448 14612
rect 17868 14560 17920 14612
rect 18144 14560 18196 14612
rect 18788 14560 18840 14612
rect 20076 14560 20128 14612
rect 20812 14560 20864 14612
rect 20996 14560 21048 14612
rect 21364 14560 21416 14612
rect 22284 14560 22336 14612
rect 26240 14603 26292 14612
rect 26240 14569 26249 14603
rect 26249 14569 26283 14603
rect 26283 14569 26292 14603
rect 26240 14560 26292 14569
rect 26792 14560 26844 14612
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 14004 14356 14056 14408
rect 14372 14356 14424 14408
rect 4896 14220 4948 14272
rect 7840 14220 7892 14272
rect 9956 14220 10008 14272
rect 10968 14263 11020 14272
rect 10968 14229 10977 14263
rect 10977 14229 11011 14263
rect 11011 14229 11020 14263
rect 10968 14220 11020 14229
rect 13728 14288 13780 14340
rect 14832 14467 14884 14476
rect 14832 14433 14841 14467
rect 14841 14433 14875 14467
rect 14875 14433 14884 14467
rect 14832 14424 14884 14433
rect 16028 14424 16080 14476
rect 18328 14467 18380 14476
rect 18328 14433 18337 14467
rect 18337 14433 18371 14467
rect 18371 14433 18380 14467
rect 18328 14424 18380 14433
rect 19432 14492 19484 14544
rect 20352 14492 20404 14544
rect 22836 14492 22888 14544
rect 19064 14424 19116 14476
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 18052 14399 18104 14408
rect 18052 14365 18061 14399
rect 18061 14365 18095 14399
rect 18095 14365 18104 14399
rect 18052 14356 18104 14365
rect 15476 14288 15528 14340
rect 14832 14220 14884 14272
rect 15292 14263 15344 14272
rect 15292 14229 15301 14263
rect 15301 14229 15335 14263
rect 15335 14229 15344 14263
rect 15292 14220 15344 14229
rect 16120 14220 16172 14272
rect 16948 14220 17000 14272
rect 17592 14220 17644 14272
rect 18512 14220 18564 14272
rect 18604 14220 18656 14272
rect 20628 14424 20680 14476
rect 22008 14424 22060 14476
rect 22376 14467 22428 14476
rect 22376 14433 22394 14467
rect 22394 14433 22428 14467
rect 22376 14424 22428 14433
rect 20076 14356 20128 14408
rect 22744 14356 22796 14408
rect 19524 14220 19576 14272
rect 20352 14220 20404 14272
rect 21364 14220 21416 14272
rect 22652 14220 22704 14272
rect 22928 14288 22980 14340
rect 23296 14424 23348 14476
rect 23572 14424 23624 14476
rect 26424 14492 26476 14544
rect 23848 14356 23900 14408
rect 24860 14399 24912 14408
rect 24860 14365 24869 14399
rect 24869 14365 24903 14399
rect 24903 14365 24912 14399
rect 24860 14356 24912 14365
rect 26424 14399 26476 14408
rect 26424 14365 26433 14399
rect 26433 14365 26467 14399
rect 26467 14365 26476 14399
rect 26424 14356 26476 14365
rect 24400 14220 24452 14272
rect 26608 14220 26660 14272
rect 3756 14118 3808 14170
rect 3820 14118 3872 14170
rect 3884 14118 3936 14170
rect 3948 14118 4000 14170
rect 4012 14118 4064 14170
rect 10472 14118 10524 14170
rect 10536 14118 10588 14170
rect 10600 14118 10652 14170
rect 10664 14118 10716 14170
rect 10728 14118 10780 14170
rect 17188 14118 17240 14170
rect 17252 14118 17304 14170
rect 17316 14118 17368 14170
rect 17380 14118 17432 14170
rect 17444 14118 17496 14170
rect 23904 14118 23956 14170
rect 23968 14118 24020 14170
rect 24032 14118 24084 14170
rect 24096 14118 24148 14170
rect 24160 14118 24212 14170
rect 3240 14059 3292 14068
rect 3240 14025 3249 14059
rect 3249 14025 3283 14059
rect 3283 14025 3292 14059
rect 3240 14016 3292 14025
rect 4160 14016 4212 14068
rect 4712 14016 4764 14068
rect 2688 13812 2740 13864
rect 3424 13812 3476 13864
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 5172 13948 5224 14000
rect 6736 14016 6788 14068
rect 4620 13880 4672 13932
rect 1768 13787 1820 13796
rect 1768 13753 1802 13787
rect 1802 13753 1820 13787
rect 1768 13744 1820 13753
rect 2412 13744 2464 13796
rect 4160 13855 4212 13864
rect 4160 13821 4169 13855
rect 4169 13821 4203 13855
rect 4203 13821 4212 13855
rect 4160 13812 4212 13821
rect 4252 13812 4304 13864
rect 4344 13812 4396 13864
rect 4896 13855 4948 13864
rect 4896 13821 4905 13855
rect 4905 13821 4939 13855
rect 4939 13821 4948 13855
rect 4896 13812 4948 13821
rect 6184 13855 6236 13864
rect 6184 13821 6193 13855
rect 6193 13821 6227 13855
rect 6227 13821 6236 13855
rect 6184 13812 6236 13821
rect 1952 13676 2004 13728
rect 3608 13676 3660 13728
rect 4160 13676 4212 13728
rect 5080 13676 5132 13728
rect 5264 13676 5316 13728
rect 6920 13812 6972 13864
rect 7748 14016 7800 14068
rect 7564 13991 7616 14000
rect 7564 13957 7573 13991
rect 7573 13957 7607 13991
rect 7607 13957 7616 13991
rect 7564 13948 7616 13957
rect 8208 13991 8260 14000
rect 8208 13957 8217 13991
rect 8217 13957 8251 13991
rect 8251 13957 8260 13991
rect 8208 13948 8260 13957
rect 8300 13812 8352 13864
rect 9864 14016 9916 14068
rect 12072 14016 12124 14068
rect 14372 14016 14424 14068
rect 16396 14059 16448 14068
rect 16396 14025 16405 14059
rect 16405 14025 16439 14059
rect 16439 14025 16448 14059
rect 16396 14016 16448 14025
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 7748 13719 7800 13728
rect 7748 13685 7757 13719
rect 7757 13685 7791 13719
rect 7791 13685 7800 13719
rect 7748 13676 7800 13685
rect 8392 13744 8444 13796
rect 16672 13948 16724 14000
rect 18604 14016 18656 14068
rect 20168 14059 20220 14068
rect 20168 14025 20177 14059
rect 20177 14025 20211 14059
rect 20211 14025 20220 14059
rect 20168 14016 20220 14025
rect 22008 14016 22060 14068
rect 17040 13948 17092 14000
rect 9680 13812 9732 13864
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 9772 13744 9824 13796
rect 10140 13787 10192 13796
rect 10140 13753 10149 13787
rect 10149 13753 10183 13787
rect 10183 13753 10192 13787
rect 10140 13744 10192 13753
rect 11980 13812 12032 13864
rect 8484 13676 8536 13728
rect 9404 13676 9456 13728
rect 10508 13719 10560 13728
rect 10508 13685 10517 13719
rect 10517 13685 10551 13719
rect 10551 13685 10560 13719
rect 10508 13676 10560 13685
rect 10876 13787 10928 13796
rect 10876 13753 10910 13787
rect 10910 13753 10928 13787
rect 10876 13744 10928 13753
rect 11520 13744 11572 13796
rect 14096 13812 14148 13864
rect 15292 13812 15344 13864
rect 16028 13855 16080 13864
rect 16028 13821 16036 13855
rect 16036 13821 16070 13855
rect 16070 13821 16080 13855
rect 16028 13812 16080 13821
rect 16120 13855 16172 13864
rect 16120 13821 16129 13855
rect 16129 13821 16163 13855
rect 16163 13821 16172 13855
rect 16120 13812 16172 13821
rect 16672 13855 16724 13864
rect 16672 13821 16681 13855
rect 16681 13821 16715 13855
rect 16715 13821 16724 13855
rect 16672 13812 16724 13821
rect 18236 13880 18288 13932
rect 20904 13948 20956 14000
rect 22928 14016 22980 14068
rect 24308 14016 24360 14068
rect 25872 14016 25924 14068
rect 11060 13676 11112 13728
rect 11336 13676 11388 13728
rect 15752 13787 15804 13796
rect 15752 13753 15761 13787
rect 15761 13753 15795 13787
rect 15795 13753 15804 13787
rect 15752 13744 15804 13753
rect 17040 13855 17092 13864
rect 17040 13821 17049 13855
rect 17049 13821 17083 13855
rect 17083 13821 17092 13855
rect 17040 13812 17092 13821
rect 17960 13812 18012 13864
rect 18328 13812 18380 13864
rect 18512 13812 18564 13864
rect 19524 13812 19576 13864
rect 19800 13855 19852 13864
rect 19800 13821 19809 13855
rect 19809 13821 19843 13855
rect 19843 13821 19852 13855
rect 19800 13812 19852 13821
rect 19892 13855 19944 13864
rect 19892 13821 19901 13855
rect 19901 13821 19935 13855
rect 19935 13821 19944 13855
rect 19892 13812 19944 13821
rect 20260 13812 20312 13864
rect 12072 13676 12124 13728
rect 17224 13744 17276 13796
rect 17592 13744 17644 13796
rect 18604 13744 18656 13796
rect 19248 13744 19300 13796
rect 20536 13855 20588 13864
rect 20536 13821 20545 13855
rect 20545 13821 20579 13855
rect 20579 13821 20588 13855
rect 20536 13812 20588 13821
rect 20720 13812 20772 13864
rect 21088 13855 21140 13864
rect 21088 13821 21095 13855
rect 21095 13821 21140 13855
rect 19432 13719 19484 13728
rect 19432 13685 19441 13719
rect 19441 13685 19475 13719
rect 19475 13685 19484 13719
rect 19432 13676 19484 13685
rect 20260 13676 20312 13728
rect 20812 13676 20864 13728
rect 21088 13812 21140 13821
rect 21180 13855 21232 13864
rect 21180 13821 21189 13855
rect 21189 13821 21223 13855
rect 21223 13821 21232 13855
rect 21180 13812 21232 13821
rect 21272 13855 21324 13864
rect 21272 13821 21281 13855
rect 21281 13821 21315 13855
rect 21315 13821 21324 13855
rect 21272 13812 21324 13821
rect 21364 13855 21416 13864
rect 21364 13821 21378 13855
rect 21378 13821 21412 13855
rect 21412 13821 21416 13855
rect 21364 13812 21416 13821
rect 21732 13812 21784 13864
rect 21824 13855 21876 13864
rect 21824 13821 21833 13855
rect 21833 13821 21867 13855
rect 21867 13821 21876 13855
rect 21824 13812 21876 13821
rect 22100 13812 22152 13864
rect 23204 13880 23256 13932
rect 22744 13812 22796 13864
rect 22652 13744 22704 13796
rect 24216 13812 24268 13864
rect 24492 13880 24544 13932
rect 24400 13855 24452 13864
rect 24400 13821 24409 13855
rect 24409 13821 24443 13855
rect 24443 13821 24452 13855
rect 24400 13812 24452 13821
rect 26332 13948 26384 14000
rect 26516 13948 26568 14000
rect 21732 13676 21784 13728
rect 22376 13719 22428 13728
rect 22376 13685 22385 13719
rect 22385 13685 22419 13719
rect 22419 13685 22428 13719
rect 22376 13676 22428 13685
rect 23204 13676 23256 13728
rect 24952 13855 25004 13864
rect 24952 13821 24961 13855
rect 24961 13821 24995 13855
rect 24995 13821 25004 13855
rect 24952 13812 25004 13821
rect 25964 13855 26016 13864
rect 25964 13821 25973 13855
rect 25973 13821 26007 13855
rect 26007 13821 26016 13855
rect 25964 13812 26016 13821
rect 26056 13855 26108 13864
rect 26056 13821 26070 13855
rect 26070 13821 26104 13855
rect 26104 13821 26108 13855
rect 26056 13812 26108 13821
rect 26516 13855 26568 13864
rect 26516 13821 26523 13855
rect 26523 13821 26568 13855
rect 26516 13812 26568 13821
rect 26608 13855 26660 13864
rect 26608 13821 26617 13855
rect 26617 13821 26651 13855
rect 26651 13821 26660 13855
rect 26608 13812 26660 13821
rect 26700 13855 26752 13864
rect 26700 13821 26709 13855
rect 26709 13821 26743 13855
rect 26743 13821 26752 13855
rect 26700 13812 26752 13821
rect 26792 13855 26844 13864
rect 26792 13821 26806 13855
rect 26806 13821 26840 13855
rect 26840 13821 26844 13855
rect 26792 13812 26844 13821
rect 25412 13676 25464 13728
rect 26240 13719 26292 13728
rect 26240 13685 26249 13719
rect 26249 13685 26283 13719
rect 26283 13685 26292 13719
rect 26240 13676 26292 13685
rect 7114 13574 7166 13626
rect 7178 13574 7230 13626
rect 7242 13574 7294 13626
rect 7306 13574 7358 13626
rect 7370 13574 7422 13626
rect 13830 13574 13882 13626
rect 13894 13574 13946 13626
rect 13958 13574 14010 13626
rect 14022 13574 14074 13626
rect 14086 13574 14138 13626
rect 20546 13574 20598 13626
rect 20610 13574 20662 13626
rect 20674 13574 20726 13626
rect 20738 13574 20790 13626
rect 20802 13574 20854 13626
rect 27262 13574 27314 13626
rect 27326 13574 27378 13626
rect 27390 13574 27442 13626
rect 27454 13574 27506 13626
rect 27518 13574 27570 13626
rect 4160 13472 4212 13524
rect 5908 13515 5960 13524
rect 1952 13447 2004 13456
rect 1952 13413 1961 13447
rect 1961 13413 1995 13447
rect 1995 13413 2004 13447
rect 1952 13404 2004 13413
rect 3608 13404 3660 13456
rect 5264 13447 5316 13456
rect 5264 13413 5273 13447
rect 5273 13413 5307 13447
rect 5307 13413 5316 13447
rect 5264 13404 5316 13413
rect 5908 13481 5917 13515
rect 5917 13481 5951 13515
rect 5951 13481 5960 13515
rect 5908 13472 5960 13481
rect 6920 13472 6972 13524
rect 5540 13404 5592 13456
rect 2228 13268 2280 13320
rect 2688 13379 2740 13388
rect 2688 13345 2697 13379
rect 2697 13345 2731 13379
rect 2731 13345 2740 13379
rect 2688 13336 2740 13345
rect 2964 13336 3016 13388
rect 5172 13379 5224 13388
rect 5172 13345 5181 13379
rect 5181 13345 5215 13379
rect 5215 13345 5224 13379
rect 5172 13336 5224 13345
rect 7564 13404 7616 13456
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 3424 13311 3476 13320
rect 3424 13277 3433 13311
rect 3433 13277 3467 13311
rect 3467 13277 3476 13311
rect 3424 13268 3476 13277
rect 4804 13268 4856 13320
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 2044 13175 2096 13184
rect 2044 13141 2053 13175
rect 2053 13141 2087 13175
rect 2087 13141 2096 13175
rect 2044 13132 2096 13141
rect 5080 13200 5132 13252
rect 6828 13336 6880 13388
rect 7196 13379 7248 13388
rect 7196 13345 7230 13379
rect 7230 13345 7248 13379
rect 7196 13336 7248 13345
rect 3332 13132 3384 13184
rect 4160 13132 4212 13184
rect 4988 13175 5040 13184
rect 4988 13141 4997 13175
rect 4997 13141 5031 13175
rect 5031 13141 5040 13175
rect 4988 13132 5040 13141
rect 7564 13132 7616 13184
rect 9680 13336 9732 13388
rect 10508 13404 10560 13456
rect 10876 13472 10928 13524
rect 11336 13472 11388 13524
rect 10876 13336 10928 13388
rect 11060 13379 11112 13388
rect 11060 13345 11069 13379
rect 11069 13345 11103 13379
rect 11103 13345 11112 13379
rect 11060 13336 11112 13345
rect 15476 13472 15528 13524
rect 15752 13472 15804 13524
rect 18052 13472 18104 13524
rect 18144 13472 18196 13524
rect 21088 13515 21140 13524
rect 21088 13481 21097 13515
rect 21097 13481 21131 13515
rect 21131 13481 21140 13515
rect 21088 13472 21140 13481
rect 24952 13472 25004 13524
rect 11336 13379 11388 13388
rect 11336 13345 11345 13379
rect 11345 13345 11379 13379
rect 11379 13345 11388 13379
rect 11336 13336 11388 13345
rect 9772 13268 9824 13320
rect 9680 13200 9732 13252
rect 10692 13268 10744 13320
rect 12164 13336 12216 13388
rect 13360 13311 13412 13320
rect 13360 13277 13369 13311
rect 13369 13277 13403 13311
rect 13403 13277 13412 13311
rect 13360 13268 13412 13277
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 15016 13379 15068 13388
rect 15016 13345 15025 13379
rect 15025 13345 15059 13379
rect 15059 13345 15068 13379
rect 15016 13336 15068 13345
rect 18236 13404 18288 13456
rect 19340 13404 19392 13456
rect 18052 13379 18104 13388
rect 18052 13345 18061 13379
rect 18061 13345 18095 13379
rect 18095 13345 18104 13379
rect 18052 13336 18104 13345
rect 18144 13379 18196 13388
rect 18144 13345 18153 13379
rect 18153 13345 18187 13379
rect 18187 13345 18196 13379
rect 18144 13336 18196 13345
rect 18328 13379 18380 13388
rect 18328 13345 18337 13379
rect 18337 13345 18371 13379
rect 18371 13345 18380 13379
rect 18328 13336 18380 13345
rect 15108 13268 15160 13320
rect 15476 13268 15528 13320
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 16948 13311 17000 13320
rect 16948 13277 16957 13311
rect 16957 13277 16991 13311
rect 16991 13277 17000 13311
rect 16948 13268 17000 13277
rect 17224 13268 17276 13320
rect 19432 13336 19484 13388
rect 22376 13404 22428 13456
rect 19984 13379 20036 13388
rect 19984 13345 20018 13379
rect 20018 13345 20036 13379
rect 19984 13336 20036 13345
rect 21180 13336 21232 13388
rect 21640 13379 21692 13388
rect 21640 13345 21649 13379
rect 21649 13345 21683 13379
rect 21683 13345 21692 13379
rect 21640 13336 21692 13345
rect 22836 13336 22888 13388
rect 26516 13336 26568 13388
rect 25228 13268 25280 13320
rect 8392 13175 8444 13184
rect 8392 13141 8401 13175
rect 8401 13141 8435 13175
rect 8435 13141 8444 13175
rect 8392 13132 8444 13141
rect 8852 13132 8904 13184
rect 10048 13132 10100 13184
rect 10784 13132 10836 13184
rect 11704 13175 11756 13184
rect 11704 13141 11713 13175
rect 11713 13141 11747 13175
rect 11747 13141 11756 13175
rect 11704 13132 11756 13141
rect 13636 13175 13688 13184
rect 13636 13141 13645 13175
rect 13645 13141 13679 13175
rect 13679 13141 13688 13175
rect 13636 13132 13688 13141
rect 14372 13132 14424 13184
rect 17592 13175 17644 13184
rect 17592 13141 17601 13175
rect 17601 13141 17635 13175
rect 17635 13141 17644 13175
rect 17592 13132 17644 13141
rect 18972 13175 19024 13184
rect 18972 13141 18981 13175
rect 18981 13141 19015 13175
rect 19015 13141 19024 13175
rect 18972 13132 19024 13141
rect 23480 13132 23532 13184
rect 25780 13132 25832 13184
rect 3756 13030 3808 13082
rect 3820 13030 3872 13082
rect 3884 13030 3936 13082
rect 3948 13030 4000 13082
rect 4012 13030 4064 13082
rect 10472 13030 10524 13082
rect 10536 13030 10588 13082
rect 10600 13030 10652 13082
rect 10664 13030 10716 13082
rect 10728 13030 10780 13082
rect 17188 13030 17240 13082
rect 17252 13030 17304 13082
rect 17316 13030 17368 13082
rect 17380 13030 17432 13082
rect 17444 13030 17496 13082
rect 23904 13030 23956 13082
rect 23968 13030 24020 13082
rect 24032 13030 24084 13082
rect 24096 13030 24148 13082
rect 24160 13030 24212 13082
rect 2964 12971 3016 12980
rect 2964 12937 2973 12971
rect 2973 12937 3007 12971
rect 3007 12937 3016 12971
rect 2964 12928 3016 12937
rect 3424 12928 3476 12980
rect 5080 12928 5132 12980
rect 7196 12928 7248 12980
rect 2412 12724 2464 12776
rect 3608 12792 3660 12844
rect 4712 12903 4764 12912
rect 4712 12869 4721 12903
rect 4721 12869 4755 12903
rect 4755 12869 4764 12903
rect 4712 12860 4764 12869
rect 6460 12860 6512 12912
rect 6828 12860 6880 12912
rect 10876 12928 10928 12980
rect 11796 12928 11848 12980
rect 13176 12928 13228 12980
rect 7748 12860 7800 12912
rect 8392 12860 8444 12912
rect 3424 12767 3476 12776
rect 2044 12656 2096 12708
rect 2688 12656 2740 12708
rect 3424 12733 3430 12767
rect 3430 12733 3464 12767
rect 3464 12733 3476 12767
rect 3424 12724 3476 12733
rect 3700 12724 3752 12776
rect 3332 12656 3384 12708
rect 4160 12724 4212 12776
rect 4344 12656 4396 12708
rect 3240 12631 3292 12640
rect 3240 12597 3249 12631
rect 3249 12597 3283 12631
rect 3283 12597 3292 12631
rect 3240 12588 3292 12597
rect 3424 12631 3476 12640
rect 3424 12597 3433 12631
rect 3433 12597 3467 12631
rect 3467 12597 3476 12631
rect 3424 12588 3476 12597
rect 3700 12588 3752 12640
rect 6092 12724 6144 12776
rect 6736 12724 6788 12776
rect 7564 12767 7616 12776
rect 7564 12733 7573 12767
rect 7573 12733 7607 12767
rect 7607 12733 7616 12767
rect 7564 12724 7616 12733
rect 8668 12792 8720 12844
rect 5264 12656 5316 12708
rect 8116 12724 8168 12776
rect 10968 12860 11020 12912
rect 15476 12971 15528 12980
rect 15476 12937 15485 12971
rect 15485 12937 15519 12971
rect 15519 12937 15528 12971
rect 15476 12928 15528 12937
rect 16948 12928 17000 12980
rect 17316 12928 17368 12980
rect 18052 12928 18104 12980
rect 20444 12928 20496 12980
rect 22836 12928 22888 12980
rect 25228 12971 25280 12980
rect 25228 12937 25237 12971
rect 25237 12937 25271 12971
rect 25271 12937 25280 12971
rect 25228 12928 25280 12937
rect 26516 12928 26568 12980
rect 24400 12860 24452 12912
rect 24860 12860 24912 12912
rect 9680 12792 9732 12844
rect 9864 12792 9916 12844
rect 12072 12792 12124 12844
rect 17960 12835 18012 12844
rect 17960 12801 17969 12835
rect 17969 12801 18003 12835
rect 18003 12801 18012 12835
rect 18696 12835 18748 12844
rect 17960 12792 18012 12801
rect 18696 12801 18705 12835
rect 18705 12801 18739 12835
rect 18739 12801 18748 12835
rect 18696 12792 18748 12801
rect 21088 12835 21140 12844
rect 21088 12801 21097 12835
rect 21097 12801 21131 12835
rect 21131 12801 21140 12835
rect 21088 12792 21140 12801
rect 23480 12792 23532 12844
rect 9956 12767 10008 12776
rect 9956 12733 9965 12767
rect 9965 12733 9999 12767
rect 9999 12733 10008 12767
rect 9956 12724 10008 12733
rect 10140 12724 10192 12776
rect 11980 12724 12032 12776
rect 14188 12724 14240 12776
rect 14372 12767 14424 12776
rect 14372 12733 14406 12767
rect 14406 12733 14424 12767
rect 14372 12724 14424 12733
rect 14832 12724 14884 12776
rect 16120 12724 16172 12776
rect 17132 12724 17184 12776
rect 20260 12724 20312 12776
rect 23204 12724 23256 12776
rect 24308 12767 24360 12776
rect 24308 12733 24322 12767
rect 24322 12733 24356 12767
rect 24356 12733 24360 12767
rect 24308 12724 24360 12733
rect 24676 12724 24728 12776
rect 25044 12792 25096 12844
rect 6276 12631 6328 12640
rect 6276 12597 6285 12631
rect 6285 12597 6319 12631
rect 6319 12597 6328 12631
rect 6276 12588 6328 12597
rect 13176 12656 13228 12708
rect 8668 12588 8720 12640
rect 9772 12631 9824 12640
rect 9772 12597 9781 12631
rect 9781 12597 9815 12631
rect 9815 12597 9824 12631
rect 9772 12588 9824 12597
rect 10048 12588 10100 12640
rect 16948 12656 17000 12708
rect 21640 12699 21692 12708
rect 21640 12665 21649 12699
rect 21649 12665 21683 12699
rect 21683 12665 21692 12699
rect 21640 12656 21692 12665
rect 22928 12656 22980 12708
rect 23388 12656 23440 12708
rect 25412 12724 25464 12776
rect 19432 12588 19484 12640
rect 20260 12588 20312 12640
rect 20352 12588 20404 12640
rect 23572 12588 23624 12640
rect 24308 12588 24360 12640
rect 24400 12588 24452 12640
rect 25596 12699 25648 12708
rect 25596 12665 25630 12699
rect 25630 12665 25648 12699
rect 25596 12656 25648 12665
rect 25044 12588 25096 12640
rect 25872 12588 25924 12640
rect 7114 12486 7166 12538
rect 7178 12486 7230 12538
rect 7242 12486 7294 12538
rect 7306 12486 7358 12538
rect 7370 12486 7422 12538
rect 13830 12486 13882 12538
rect 13894 12486 13946 12538
rect 13958 12486 14010 12538
rect 14022 12486 14074 12538
rect 14086 12486 14138 12538
rect 20546 12486 20598 12538
rect 20610 12486 20662 12538
rect 20674 12486 20726 12538
rect 20738 12486 20790 12538
rect 20802 12486 20854 12538
rect 27262 12486 27314 12538
rect 27326 12486 27378 12538
rect 27390 12486 27442 12538
rect 27454 12486 27506 12538
rect 27518 12486 27570 12538
rect 3424 12384 3476 12436
rect 5264 12427 5316 12436
rect 5264 12393 5273 12427
rect 5273 12393 5307 12427
rect 5307 12393 5316 12427
rect 5264 12384 5316 12393
rect 7196 12384 7248 12436
rect 8116 12384 8168 12436
rect 9680 12384 9732 12436
rect 12164 12384 12216 12436
rect 2688 12291 2740 12300
rect 2688 12257 2697 12291
rect 2697 12257 2731 12291
rect 2731 12257 2740 12291
rect 2688 12248 2740 12257
rect 3240 12316 3292 12368
rect 3516 12248 3568 12300
rect 5632 12316 5684 12368
rect 6276 12316 6328 12368
rect 8668 12359 8720 12368
rect 8668 12325 8677 12359
rect 8677 12325 8711 12359
rect 8711 12325 8720 12359
rect 8668 12316 8720 12325
rect 4988 12291 5040 12300
rect 4988 12257 4997 12291
rect 4997 12257 5031 12291
rect 5031 12257 5040 12291
rect 4988 12248 5040 12257
rect 7196 12291 7248 12300
rect 7196 12257 7205 12291
rect 7205 12257 7239 12291
rect 7239 12257 7248 12291
rect 7196 12248 7248 12257
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 3608 12223 3660 12232
rect 3608 12189 3617 12223
rect 3617 12189 3651 12223
rect 3651 12189 3660 12223
rect 3608 12180 3660 12189
rect 4804 12223 4856 12232
rect 4804 12189 4813 12223
rect 4813 12189 4847 12223
rect 4847 12189 4856 12223
rect 4804 12180 4856 12189
rect 6644 12112 6696 12164
rect 2320 12087 2372 12096
rect 2320 12053 2329 12087
rect 2329 12053 2363 12087
rect 2363 12053 2372 12087
rect 2320 12044 2372 12053
rect 3608 12044 3660 12096
rect 6920 12044 6972 12096
rect 7564 12155 7616 12164
rect 7564 12121 7573 12155
rect 7573 12121 7607 12155
rect 7607 12121 7616 12155
rect 7564 12112 7616 12121
rect 7656 12155 7708 12164
rect 7656 12121 7665 12155
rect 7665 12121 7699 12155
rect 7699 12121 7708 12155
rect 7656 12112 7708 12121
rect 8944 12291 8996 12300
rect 8944 12257 8953 12291
rect 8953 12257 8987 12291
rect 8987 12257 8996 12291
rect 8944 12248 8996 12257
rect 9404 12248 9456 12300
rect 9864 12248 9916 12300
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 9588 12180 9640 12232
rect 10140 12223 10192 12232
rect 10140 12189 10149 12223
rect 10149 12189 10183 12223
rect 10183 12189 10192 12223
rect 11520 12248 11572 12300
rect 12072 12248 12124 12300
rect 10140 12180 10192 12189
rect 8760 12112 8812 12164
rect 9680 12087 9732 12096
rect 9680 12053 9689 12087
rect 9689 12053 9723 12087
rect 9723 12053 9732 12087
rect 9680 12044 9732 12053
rect 11612 12044 11664 12096
rect 12164 12044 12216 12096
rect 12716 12044 12768 12096
rect 13820 12384 13872 12436
rect 14280 12384 14332 12436
rect 14188 12316 14240 12368
rect 16212 12427 16264 12436
rect 16212 12393 16221 12427
rect 16221 12393 16255 12427
rect 16255 12393 16264 12427
rect 16212 12384 16264 12393
rect 16948 12427 17000 12436
rect 16948 12393 16957 12427
rect 16957 12393 16991 12427
rect 16991 12393 17000 12427
rect 16948 12384 17000 12393
rect 13636 12291 13688 12300
rect 13636 12257 13670 12291
rect 13670 12257 13688 12291
rect 13636 12248 13688 12257
rect 13912 12248 13964 12300
rect 16672 12316 16724 12368
rect 14464 12180 14516 12232
rect 14924 12180 14976 12232
rect 15936 12291 15988 12300
rect 15936 12257 15945 12291
rect 15945 12257 15979 12291
rect 15979 12257 15988 12291
rect 15936 12248 15988 12257
rect 17592 12384 17644 12436
rect 19984 12384 20036 12436
rect 22744 12427 22796 12436
rect 22744 12393 22753 12427
rect 22753 12393 22787 12427
rect 22787 12393 22796 12427
rect 22744 12384 22796 12393
rect 18972 12316 19024 12368
rect 19800 12316 19852 12368
rect 17316 12291 17368 12300
rect 17316 12257 17325 12291
rect 17325 12257 17359 12291
rect 17359 12257 17368 12291
rect 17316 12248 17368 12257
rect 18328 12248 18380 12300
rect 18696 12248 18748 12300
rect 19984 12248 20036 12300
rect 20352 12291 20404 12300
rect 20352 12257 20361 12291
rect 20361 12257 20395 12291
rect 20395 12257 20404 12291
rect 20352 12248 20404 12257
rect 21732 12316 21784 12368
rect 25044 12384 25096 12436
rect 25596 12384 25648 12436
rect 20536 12291 20588 12300
rect 20536 12257 20545 12291
rect 20545 12257 20579 12291
rect 20579 12257 20588 12291
rect 20536 12248 20588 12257
rect 23388 12316 23440 12368
rect 21272 12180 21324 12232
rect 17592 12112 17644 12164
rect 20076 12112 20128 12164
rect 23480 12291 23532 12300
rect 23480 12257 23489 12291
rect 23489 12257 23523 12291
rect 23523 12257 23532 12291
rect 23480 12248 23532 12257
rect 23480 12112 23532 12164
rect 24308 12248 24360 12300
rect 24768 12112 24820 12164
rect 25044 12291 25096 12300
rect 25044 12257 25053 12291
rect 25053 12257 25087 12291
rect 25087 12257 25096 12291
rect 25044 12248 25096 12257
rect 25964 12384 26016 12436
rect 25780 12291 25832 12300
rect 25780 12257 25789 12291
rect 25789 12257 25823 12291
rect 25823 12257 25832 12291
rect 25780 12248 25832 12257
rect 25872 12291 25924 12300
rect 25872 12257 25881 12291
rect 25881 12257 25915 12291
rect 25915 12257 25924 12291
rect 25872 12248 25924 12257
rect 26240 12316 26292 12368
rect 26240 12180 26292 12232
rect 15016 12044 15068 12096
rect 15844 12087 15896 12096
rect 15844 12053 15853 12087
rect 15853 12053 15887 12087
rect 15887 12053 15896 12087
rect 15844 12044 15896 12053
rect 16028 12044 16080 12096
rect 18972 12044 19024 12096
rect 21364 12087 21416 12096
rect 21364 12053 21373 12087
rect 21373 12053 21407 12087
rect 21407 12053 21416 12087
rect 21364 12044 21416 12053
rect 24676 12044 24728 12096
rect 25412 12087 25464 12096
rect 25412 12053 25421 12087
rect 25421 12053 25455 12087
rect 25455 12053 25464 12087
rect 25412 12044 25464 12053
rect 3756 11942 3808 11994
rect 3820 11942 3872 11994
rect 3884 11942 3936 11994
rect 3948 11942 4000 11994
rect 4012 11942 4064 11994
rect 10472 11942 10524 11994
rect 10536 11942 10588 11994
rect 10600 11942 10652 11994
rect 10664 11942 10716 11994
rect 10728 11942 10780 11994
rect 17188 11942 17240 11994
rect 17252 11942 17304 11994
rect 17316 11942 17368 11994
rect 17380 11942 17432 11994
rect 17444 11942 17496 11994
rect 23904 11942 23956 11994
rect 23968 11942 24020 11994
rect 24032 11942 24084 11994
rect 24096 11942 24148 11994
rect 24160 11942 24212 11994
rect 3608 11840 3660 11892
rect 7564 11840 7616 11892
rect 7840 11840 7892 11892
rect 9220 11840 9272 11892
rect 12072 11883 12124 11892
rect 12072 11849 12081 11883
rect 12081 11849 12115 11883
rect 12115 11849 12124 11883
rect 12072 11840 12124 11849
rect 13820 11840 13872 11892
rect 14648 11840 14700 11892
rect 4804 11772 4856 11824
rect 12440 11772 12492 11824
rect 12716 11772 12768 11824
rect 15568 11840 15620 11892
rect 17592 11840 17644 11892
rect 18144 11840 18196 11892
rect 19892 11840 19944 11892
rect 20536 11840 20588 11892
rect 21456 11840 21508 11892
rect 23480 11883 23532 11892
rect 23480 11849 23489 11883
rect 23489 11849 23523 11883
rect 23523 11849 23532 11883
rect 23480 11840 23532 11849
rect 24676 11840 24728 11892
rect 26240 11883 26292 11892
rect 26240 11849 26249 11883
rect 26249 11849 26283 11883
rect 26283 11849 26292 11883
rect 26240 11840 26292 11849
rect 2412 11636 2464 11688
rect 9956 11704 10008 11756
rect 11520 11704 11572 11756
rect 8484 11679 8536 11688
rect 8484 11645 8493 11679
rect 8493 11645 8527 11679
rect 8527 11645 8536 11679
rect 8484 11636 8536 11645
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 8852 11636 8904 11688
rect 9312 11636 9364 11688
rect 11612 11679 11664 11688
rect 11612 11645 11621 11679
rect 11621 11645 11655 11679
rect 11655 11645 11664 11679
rect 11612 11636 11664 11645
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 12164 11636 12216 11688
rect 13176 11704 13228 11756
rect 13728 11704 13780 11756
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 14372 11704 14424 11756
rect 2320 11568 2372 11620
rect 5816 11568 5868 11620
rect 6092 11568 6144 11620
rect 9588 11611 9640 11620
rect 9588 11577 9597 11611
rect 9597 11577 9631 11611
rect 9631 11577 9640 11611
rect 9588 11568 9640 11577
rect 12072 11568 12124 11620
rect 4804 11500 4856 11552
rect 8944 11500 8996 11552
rect 9956 11500 10008 11552
rect 12440 11611 12492 11620
rect 12440 11577 12449 11611
rect 12449 11577 12483 11611
rect 12483 11577 12492 11611
rect 12440 11568 12492 11577
rect 12808 11568 12860 11620
rect 13912 11636 13964 11688
rect 16120 11636 16172 11688
rect 17132 11636 17184 11688
rect 12624 11500 12676 11552
rect 14648 11543 14700 11552
rect 14648 11509 14657 11543
rect 14657 11509 14691 11543
rect 14691 11509 14700 11543
rect 14648 11500 14700 11509
rect 15016 11500 15068 11552
rect 15568 11543 15620 11552
rect 15568 11509 15577 11543
rect 15577 11509 15611 11543
rect 15611 11509 15620 11543
rect 15568 11500 15620 11509
rect 15660 11543 15712 11552
rect 15660 11509 15669 11543
rect 15669 11509 15703 11543
rect 15703 11509 15712 11543
rect 15660 11500 15712 11509
rect 16948 11500 17000 11552
rect 17040 11543 17092 11552
rect 17040 11509 17049 11543
rect 17049 11509 17083 11543
rect 17083 11509 17092 11543
rect 17040 11500 17092 11509
rect 17132 11500 17184 11552
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 18972 11772 19024 11824
rect 18788 11679 18840 11688
rect 18788 11645 18798 11679
rect 18798 11645 18832 11679
rect 18832 11645 18840 11679
rect 18788 11636 18840 11645
rect 19340 11636 19392 11688
rect 19432 11679 19484 11688
rect 19432 11645 19441 11679
rect 19441 11645 19475 11679
rect 19475 11645 19484 11679
rect 19432 11636 19484 11645
rect 19524 11679 19576 11688
rect 19524 11645 19534 11679
rect 19534 11645 19568 11679
rect 19568 11645 19576 11679
rect 19524 11636 19576 11645
rect 24400 11747 24452 11756
rect 24400 11713 24409 11747
rect 24409 11713 24443 11747
rect 24443 11713 24452 11747
rect 24400 11704 24452 11713
rect 24860 11747 24912 11756
rect 24860 11713 24869 11747
rect 24869 11713 24903 11747
rect 24903 11713 24912 11747
rect 24860 11704 24912 11713
rect 19892 11679 19944 11688
rect 19892 11645 19906 11679
rect 19906 11645 19940 11679
rect 19940 11645 19944 11679
rect 19892 11636 19944 11645
rect 20444 11636 20496 11688
rect 21180 11636 21232 11688
rect 22836 11636 22888 11688
rect 25412 11636 25464 11688
rect 26240 11636 26292 11688
rect 26700 11636 26752 11688
rect 18972 11500 19024 11552
rect 19800 11611 19852 11620
rect 19800 11577 19809 11611
rect 19809 11577 19843 11611
rect 19843 11577 19852 11611
rect 19800 11568 19852 11577
rect 21364 11611 21416 11620
rect 21364 11577 21398 11611
rect 21398 11577 21416 11611
rect 21364 11568 21416 11577
rect 20260 11500 20312 11552
rect 23664 11500 23716 11552
rect 25136 11500 25188 11552
rect 7114 11398 7166 11450
rect 7178 11398 7230 11450
rect 7242 11398 7294 11450
rect 7306 11398 7358 11450
rect 7370 11398 7422 11450
rect 13830 11398 13882 11450
rect 13894 11398 13946 11450
rect 13958 11398 14010 11450
rect 14022 11398 14074 11450
rect 14086 11398 14138 11450
rect 20546 11398 20598 11450
rect 20610 11398 20662 11450
rect 20674 11398 20726 11450
rect 20738 11398 20790 11450
rect 20802 11398 20854 11450
rect 27262 11398 27314 11450
rect 27326 11398 27378 11450
rect 27390 11398 27442 11450
rect 27454 11398 27506 11450
rect 27518 11398 27570 11450
rect 3516 11339 3568 11348
rect 3516 11305 3525 11339
rect 3525 11305 3559 11339
rect 3559 11305 3568 11339
rect 3516 11296 3568 11305
rect 6920 11228 6972 11280
rect 3424 11160 3476 11212
rect 8024 11296 8076 11348
rect 9036 11296 9088 11348
rect 9404 11296 9456 11348
rect 8116 11228 8168 11280
rect 5816 11135 5868 11144
rect 5816 11101 5825 11135
rect 5825 11101 5859 11135
rect 5859 11101 5868 11135
rect 5816 11092 5868 11101
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 8208 11203 8260 11212
rect 8208 11169 8217 11203
rect 8217 11169 8251 11203
rect 8251 11169 8260 11203
rect 8208 11160 8260 11169
rect 9312 11228 9364 11280
rect 9680 11228 9732 11280
rect 8300 11092 8352 11144
rect 8668 11203 8720 11212
rect 8668 11169 8677 11203
rect 8677 11169 8711 11203
rect 8711 11169 8720 11203
rect 8668 11160 8720 11169
rect 8760 11203 8812 11212
rect 8760 11169 8769 11203
rect 8769 11169 8803 11203
rect 8803 11169 8812 11203
rect 8760 11160 8812 11169
rect 8576 11092 8628 11144
rect 4804 11067 4856 11076
rect 4804 11033 4813 11067
rect 4813 11033 4847 11067
rect 4847 11033 4856 11067
rect 4804 11024 4856 11033
rect 6828 11024 6880 11076
rect 6736 10956 6788 11008
rect 7472 10956 7524 11008
rect 7932 10999 7984 11008
rect 7932 10965 7941 10999
rect 7941 10965 7975 10999
rect 7975 10965 7984 10999
rect 7932 10956 7984 10965
rect 9128 10999 9180 11008
rect 9128 10965 9137 10999
rect 9137 10965 9171 10999
rect 9171 10965 9180 10999
rect 9128 10956 9180 10965
rect 13728 11339 13780 11348
rect 13728 11305 13737 11339
rect 13737 11305 13771 11339
rect 13771 11305 13780 11339
rect 13728 11296 13780 11305
rect 18052 11296 18104 11348
rect 12716 11228 12768 11280
rect 18512 11339 18564 11348
rect 18512 11305 18521 11339
rect 18521 11305 18555 11339
rect 18555 11305 18564 11339
rect 18512 11296 18564 11305
rect 19248 11296 19300 11348
rect 19708 11296 19760 11348
rect 19800 11296 19852 11348
rect 21272 11339 21324 11348
rect 21272 11305 21281 11339
rect 21281 11305 21315 11339
rect 21315 11305 21324 11339
rect 21272 11296 21324 11305
rect 24400 11296 24452 11348
rect 26240 11339 26292 11348
rect 26240 11305 26249 11339
rect 26249 11305 26283 11339
rect 26283 11305 26292 11339
rect 26240 11296 26292 11305
rect 11520 11160 11572 11212
rect 14188 11160 14240 11212
rect 14832 11160 14884 11212
rect 15568 11160 15620 11212
rect 17132 11160 17184 11212
rect 19432 11228 19484 11280
rect 14464 11092 14516 11144
rect 14924 11092 14976 11144
rect 15752 11092 15804 11144
rect 16212 11092 16264 11144
rect 16948 11092 17000 11144
rect 9588 10956 9640 11008
rect 18052 11024 18104 11076
rect 18604 11203 18656 11212
rect 18604 11169 18613 11203
rect 18613 11169 18647 11203
rect 18647 11169 18656 11203
rect 18604 11160 18656 11169
rect 18788 11203 18840 11212
rect 18788 11169 18797 11203
rect 18797 11169 18831 11203
rect 18831 11169 18840 11203
rect 18788 11160 18840 11169
rect 18880 11203 18932 11212
rect 18880 11169 18889 11203
rect 18889 11169 18923 11203
rect 18923 11169 18932 11203
rect 18880 11160 18932 11169
rect 19892 11228 19944 11280
rect 20444 11160 20496 11212
rect 20720 11135 20772 11144
rect 20720 11101 20729 11135
rect 20729 11101 20763 11135
rect 20763 11101 20772 11135
rect 20720 11092 20772 11101
rect 21456 11160 21508 11212
rect 21732 11203 21784 11212
rect 21732 11169 21741 11203
rect 21741 11169 21775 11203
rect 21775 11169 21784 11203
rect 21732 11160 21784 11169
rect 21364 11024 21416 11076
rect 22284 11160 22336 11212
rect 22836 11160 22888 11212
rect 23756 11160 23808 11212
rect 24860 11203 24912 11212
rect 24860 11169 24869 11203
rect 24869 11169 24903 11203
rect 24903 11169 24912 11203
rect 24860 11160 24912 11169
rect 22744 11135 22796 11144
rect 22744 11101 22753 11135
rect 22753 11101 22787 11135
rect 22787 11101 22796 11135
rect 22744 11092 22796 11101
rect 25872 11092 25924 11144
rect 22652 11024 22704 11076
rect 14372 10956 14424 11008
rect 17592 10956 17644 11008
rect 19340 10999 19392 11008
rect 19340 10965 19349 10999
rect 19349 10965 19383 10999
rect 19383 10965 19392 10999
rect 19340 10956 19392 10965
rect 22928 10956 22980 11008
rect 3756 10854 3808 10906
rect 3820 10854 3872 10906
rect 3884 10854 3936 10906
rect 3948 10854 4000 10906
rect 4012 10854 4064 10906
rect 10472 10854 10524 10906
rect 10536 10854 10588 10906
rect 10600 10854 10652 10906
rect 10664 10854 10716 10906
rect 10728 10854 10780 10906
rect 17188 10854 17240 10906
rect 17252 10854 17304 10906
rect 17316 10854 17368 10906
rect 17380 10854 17432 10906
rect 17444 10854 17496 10906
rect 23904 10854 23956 10906
rect 23968 10854 24020 10906
rect 24032 10854 24084 10906
rect 24096 10854 24148 10906
rect 24160 10854 24212 10906
rect 7288 10752 7340 10804
rect 8668 10752 8720 10804
rect 8852 10684 8904 10736
rect 2412 10548 2464 10600
rect 5816 10591 5868 10600
rect 5816 10557 5825 10591
rect 5825 10557 5859 10591
rect 5859 10557 5868 10591
rect 5816 10548 5868 10557
rect 7748 10591 7800 10600
rect 7748 10557 7755 10591
rect 7755 10557 7800 10591
rect 5632 10480 5684 10532
rect 6092 10523 6144 10532
rect 6092 10489 6126 10523
rect 6126 10489 6144 10523
rect 6092 10480 6144 10489
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 7748 10548 7800 10557
rect 7932 10591 7984 10600
rect 7932 10557 7941 10591
rect 7941 10557 7975 10591
rect 7975 10557 7984 10591
rect 7932 10548 7984 10557
rect 8300 10548 8352 10600
rect 8576 10548 8628 10600
rect 8944 10548 8996 10600
rect 8484 10480 8536 10532
rect 8760 10480 8812 10532
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 12716 10752 12768 10804
rect 15200 10752 15252 10804
rect 12532 10684 12584 10736
rect 16948 10752 17000 10804
rect 19984 10752 20036 10804
rect 20720 10752 20772 10804
rect 21732 10752 21784 10804
rect 12624 10548 12676 10600
rect 14372 10616 14424 10668
rect 14832 10616 14884 10668
rect 15108 10616 15160 10668
rect 18696 10659 18748 10668
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 13084 10591 13136 10600
rect 13084 10557 13093 10591
rect 13093 10557 13127 10591
rect 13127 10557 13136 10591
rect 13084 10548 13136 10557
rect 15200 10591 15252 10600
rect 15200 10557 15209 10591
rect 15209 10557 15243 10591
rect 15243 10557 15252 10591
rect 15200 10548 15252 10557
rect 15292 10591 15344 10600
rect 15292 10557 15301 10591
rect 15301 10557 15335 10591
rect 15335 10557 15344 10591
rect 15292 10548 15344 10557
rect 15384 10591 15436 10600
rect 15384 10557 15393 10591
rect 15393 10557 15427 10591
rect 15427 10557 15436 10591
rect 15384 10548 15436 10557
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 17868 10591 17920 10600
rect 17868 10557 17877 10591
rect 17877 10557 17911 10591
rect 17911 10557 17920 10591
rect 17868 10548 17920 10557
rect 19340 10548 19392 10600
rect 19432 10548 19484 10600
rect 22192 10591 22244 10600
rect 8300 10412 8352 10464
rect 9220 10412 9272 10464
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 15752 10480 15804 10532
rect 15936 10480 15988 10532
rect 22192 10557 22201 10591
rect 22201 10557 22235 10591
rect 22235 10557 22244 10591
rect 22192 10548 22244 10557
rect 23572 10752 23624 10804
rect 23756 10752 23808 10804
rect 26424 10752 26476 10804
rect 22652 10684 22704 10736
rect 22008 10480 22060 10532
rect 22928 10591 22980 10600
rect 22928 10557 22937 10591
rect 22937 10557 22971 10591
rect 22971 10557 22980 10591
rect 22928 10548 22980 10557
rect 25044 10684 25096 10736
rect 24860 10616 24912 10668
rect 15016 10412 15068 10464
rect 16672 10412 16724 10464
rect 17316 10455 17368 10464
rect 17316 10421 17325 10455
rect 17325 10421 17359 10455
rect 17359 10421 17368 10455
rect 17316 10412 17368 10421
rect 19892 10412 19944 10464
rect 21732 10412 21784 10464
rect 23664 10548 23716 10600
rect 24492 10548 24544 10600
rect 24952 10548 25004 10600
rect 24676 10480 24728 10532
rect 24124 10412 24176 10464
rect 25320 10412 25372 10464
rect 7114 10310 7166 10362
rect 7178 10310 7230 10362
rect 7242 10310 7294 10362
rect 7306 10310 7358 10362
rect 7370 10310 7422 10362
rect 13830 10310 13882 10362
rect 13894 10310 13946 10362
rect 13958 10310 14010 10362
rect 14022 10310 14074 10362
rect 14086 10310 14138 10362
rect 20546 10310 20598 10362
rect 20610 10310 20662 10362
rect 20674 10310 20726 10362
rect 20738 10310 20790 10362
rect 20802 10310 20854 10362
rect 27262 10310 27314 10362
rect 27326 10310 27378 10362
rect 27390 10310 27442 10362
rect 27454 10310 27506 10362
rect 27518 10310 27570 10362
rect 3608 10208 3660 10260
rect 6092 10208 6144 10260
rect 8208 10208 8260 10260
rect 8576 10208 8628 10260
rect 8760 10208 8812 10260
rect 8944 10251 8996 10260
rect 8944 10217 8953 10251
rect 8953 10217 8987 10251
rect 8987 10217 8996 10251
rect 8944 10208 8996 10217
rect 12164 10208 12216 10260
rect 12900 10208 12952 10260
rect 12992 10208 13044 10260
rect 14556 10208 14608 10260
rect 15384 10208 15436 10260
rect 15936 10208 15988 10260
rect 17316 10208 17368 10260
rect 20260 10251 20312 10260
rect 20260 10217 20269 10251
rect 20269 10217 20303 10251
rect 20303 10217 20312 10251
rect 20260 10208 20312 10217
rect 21824 10208 21876 10260
rect 22100 10251 22152 10260
rect 22100 10217 22109 10251
rect 22109 10217 22143 10251
rect 22143 10217 22152 10251
rect 22100 10208 22152 10217
rect 23020 10208 23072 10260
rect 23296 10208 23348 10260
rect 25872 10208 25924 10260
rect 2872 10140 2924 10192
rect 5724 10140 5776 10192
rect 2412 10115 2464 10124
rect 2412 10081 2421 10115
rect 2421 10081 2455 10115
rect 2455 10081 2464 10115
rect 2412 10072 2464 10081
rect 3424 10072 3476 10124
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 6092 10072 6144 10124
rect 1860 9936 1912 9988
rect 6644 10115 6696 10124
rect 6644 10081 6653 10115
rect 6653 10081 6687 10115
rect 6687 10081 6696 10115
rect 6644 10072 6696 10081
rect 4988 9936 5040 9988
rect 3056 9868 3108 9920
rect 4160 9868 4212 9920
rect 5540 9868 5592 9920
rect 6368 9979 6420 9988
rect 6368 9945 6377 9979
rect 6377 9945 6411 9979
rect 6411 9945 6420 9979
rect 6368 9936 6420 9945
rect 7196 10115 7248 10124
rect 7196 10081 7205 10115
rect 7205 10081 7239 10115
rect 7239 10081 7248 10115
rect 7196 10072 7248 10081
rect 8300 10115 8352 10124
rect 8300 10081 8309 10115
rect 8309 10081 8343 10115
rect 8343 10081 8352 10115
rect 8300 10072 8352 10081
rect 7932 10004 7984 10056
rect 7656 9936 7708 9988
rect 8576 10115 8628 10124
rect 8576 10081 8585 10115
rect 8585 10081 8619 10115
rect 8619 10081 8628 10115
rect 8576 10072 8628 10081
rect 8852 10072 8904 10124
rect 9588 10140 9640 10192
rect 9128 10072 9180 10124
rect 12348 10140 12400 10192
rect 14280 10140 14332 10192
rect 12256 10115 12308 10124
rect 12256 10081 12266 10115
rect 12266 10081 12300 10115
rect 12300 10081 12308 10115
rect 12256 10072 12308 10081
rect 8944 10004 8996 10056
rect 12624 10115 12676 10124
rect 12624 10081 12638 10115
rect 12638 10081 12672 10115
rect 12672 10081 12676 10115
rect 12624 10072 12676 10081
rect 13360 10072 13412 10124
rect 13452 10004 13504 10056
rect 9036 9936 9088 9988
rect 13728 9936 13780 9988
rect 6460 9868 6512 9920
rect 7196 9868 7248 9920
rect 8208 9868 8260 9920
rect 8668 9868 8720 9920
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 14832 10004 14884 10056
rect 16580 10072 16632 10124
rect 16672 10115 16724 10124
rect 16672 10081 16681 10115
rect 16681 10081 16715 10115
rect 16715 10081 16724 10115
rect 16672 10072 16724 10081
rect 16856 10072 16908 10124
rect 15108 10004 15160 10056
rect 17592 10072 17644 10124
rect 18696 10072 18748 10124
rect 22376 10140 22428 10192
rect 24124 10140 24176 10192
rect 17776 10004 17828 10056
rect 18236 10047 18288 10056
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 20168 10004 20220 10056
rect 21732 10115 21784 10124
rect 21732 10081 21741 10115
rect 21741 10081 21775 10115
rect 21775 10081 21784 10115
rect 21732 10072 21784 10081
rect 22008 10115 22060 10124
rect 22008 10081 22017 10115
rect 22017 10081 22051 10115
rect 22051 10081 22060 10115
rect 22008 10072 22060 10081
rect 22192 10072 22244 10124
rect 17868 9936 17920 9988
rect 23296 10115 23348 10124
rect 23296 10081 23305 10115
rect 23305 10081 23339 10115
rect 23339 10081 23348 10115
rect 23296 10072 23348 10081
rect 23388 10115 23440 10124
rect 23388 10081 23397 10115
rect 23397 10081 23431 10115
rect 23431 10081 23440 10115
rect 23388 10072 23440 10081
rect 23756 10072 23808 10124
rect 24308 10115 24360 10124
rect 24308 10081 24317 10115
rect 24317 10081 24351 10115
rect 24351 10081 24360 10115
rect 24308 10072 24360 10081
rect 24400 10115 24452 10124
rect 24400 10081 24409 10115
rect 24409 10081 24443 10115
rect 24443 10081 24452 10115
rect 24400 10072 24452 10081
rect 24860 10004 24912 10056
rect 25044 10115 25096 10124
rect 25044 10081 25053 10115
rect 25053 10081 25087 10115
rect 25087 10081 25096 10115
rect 25044 10072 25096 10081
rect 25136 10115 25188 10124
rect 25136 10081 25145 10115
rect 25145 10081 25179 10115
rect 25179 10081 25188 10115
rect 25136 10072 25188 10081
rect 25228 10072 25280 10124
rect 25872 10115 25924 10124
rect 25872 10081 25881 10115
rect 25881 10081 25915 10115
rect 25915 10081 25924 10115
rect 25872 10072 25924 10081
rect 15476 9868 15528 9920
rect 17040 9868 17092 9920
rect 19524 9868 19576 9920
rect 24492 9936 24544 9988
rect 24676 9979 24728 9988
rect 24676 9945 24685 9979
rect 24685 9945 24719 9979
rect 24719 9945 24728 9979
rect 24676 9936 24728 9945
rect 24952 9936 25004 9988
rect 26424 10072 26476 10124
rect 26424 9979 26476 9988
rect 26424 9945 26433 9979
rect 26433 9945 26467 9979
rect 26467 9945 26476 9979
rect 26424 9936 26476 9945
rect 24308 9868 24360 9920
rect 25044 9868 25096 9920
rect 3756 9766 3808 9818
rect 3820 9766 3872 9818
rect 3884 9766 3936 9818
rect 3948 9766 4000 9818
rect 4012 9766 4064 9818
rect 10472 9766 10524 9818
rect 10536 9766 10588 9818
rect 10600 9766 10652 9818
rect 10664 9766 10716 9818
rect 10728 9766 10780 9818
rect 17188 9766 17240 9818
rect 17252 9766 17304 9818
rect 17316 9766 17368 9818
rect 17380 9766 17432 9818
rect 17444 9766 17496 9818
rect 23904 9766 23956 9818
rect 23968 9766 24020 9818
rect 24032 9766 24084 9818
rect 24096 9766 24148 9818
rect 24160 9766 24212 9818
rect 6368 9664 6420 9716
rect 13452 9664 13504 9716
rect 16028 9664 16080 9716
rect 2872 9639 2924 9648
rect 2872 9605 2881 9639
rect 2881 9605 2915 9639
rect 2915 9605 2924 9639
rect 2872 9596 2924 9605
rect 3608 9596 3660 9648
rect 5540 9596 5592 9648
rect 5632 9528 5684 9580
rect 2412 9460 2464 9512
rect 3056 9503 3108 9512
rect 3056 9469 3065 9503
rect 3065 9469 3099 9503
rect 3099 9469 3108 9503
rect 3056 9460 3108 9469
rect 3608 9460 3660 9512
rect 4160 9503 4212 9512
rect 4160 9469 4169 9503
rect 4169 9469 4203 9503
rect 4203 9469 4212 9503
rect 4160 9460 4212 9469
rect 4436 9503 4488 9512
rect 4436 9469 4445 9503
rect 4445 9469 4479 9503
rect 4479 9469 4488 9503
rect 4436 9460 4488 9469
rect 1676 9435 1728 9444
rect 1676 9401 1710 9435
rect 1710 9401 1728 9435
rect 1676 9392 1728 9401
rect 3148 9392 3200 9444
rect 5448 9503 5500 9512
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 4988 9392 5040 9444
rect 5724 9392 5776 9444
rect 6000 9503 6052 9512
rect 6000 9469 6009 9503
rect 6009 9469 6043 9503
rect 6043 9469 6052 9503
rect 6000 9460 6052 9469
rect 6828 9528 6880 9580
rect 6276 9460 6328 9512
rect 6644 9460 6696 9512
rect 8116 9460 8168 9512
rect 8760 9460 8812 9512
rect 9312 9596 9364 9648
rect 14464 9639 14516 9648
rect 14464 9605 14473 9639
rect 14473 9605 14507 9639
rect 14507 9605 14516 9639
rect 14464 9596 14516 9605
rect 15752 9596 15804 9648
rect 11520 9528 11572 9580
rect 15292 9528 15344 9580
rect 6092 9392 6144 9444
rect 6736 9392 6788 9444
rect 9220 9503 9272 9512
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9220 9460 9272 9469
rect 9496 9460 9548 9512
rect 9588 9460 9640 9512
rect 12992 9460 13044 9512
rect 13176 9460 13228 9512
rect 16120 9503 16172 9512
rect 16120 9469 16129 9503
rect 16129 9469 16163 9503
rect 16163 9469 16172 9503
rect 16120 9460 16172 9469
rect 16580 9596 16632 9648
rect 16948 9571 17000 9580
rect 16948 9537 16957 9571
rect 16957 9537 16991 9571
rect 16991 9537 17000 9571
rect 16948 9528 17000 9537
rect 17592 9596 17644 9648
rect 18236 9664 18288 9716
rect 22376 9664 22428 9716
rect 18604 9596 18656 9648
rect 17224 9528 17276 9580
rect 17500 9571 17552 9580
rect 17500 9537 17509 9571
rect 17509 9537 17543 9571
rect 17543 9537 17552 9571
rect 17500 9528 17552 9537
rect 9404 9392 9456 9444
rect 2872 9324 2924 9376
rect 4620 9324 4672 9376
rect 8392 9324 8444 9376
rect 11888 9435 11940 9444
rect 11888 9401 11922 9435
rect 11922 9401 11940 9435
rect 11888 9392 11940 9401
rect 12348 9392 12400 9444
rect 13268 9392 13320 9444
rect 15752 9435 15804 9444
rect 15752 9401 15761 9435
rect 15761 9401 15795 9435
rect 15795 9401 15804 9435
rect 15752 9392 15804 9401
rect 15936 9392 15988 9444
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 17132 9503 17184 9512
rect 17132 9469 17141 9503
rect 17141 9469 17175 9503
rect 17175 9469 17184 9503
rect 17132 9460 17184 9469
rect 17960 9460 18012 9512
rect 19524 9528 19576 9580
rect 20444 9596 20496 9648
rect 21364 9639 21416 9648
rect 21364 9605 21373 9639
rect 21373 9605 21407 9639
rect 21407 9605 21416 9639
rect 21364 9596 21416 9605
rect 21640 9596 21692 9648
rect 19340 9503 19392 9512
rect 19340 9469 19349 9503
rect 19349 9469 19383 9503
rect 19383 9469 19392 9503
rect 19340 9460 19392 9469
rect 22744 9571 22796 9580
rect 22744 9537 22753 9571
rect 22753 9537 22787 9571
rect 22787 9537 22796 9571
rect 22744 9528 22796 9537
rect 24768 9596 24820 9648
rect 24860 9639 24912 9648
rect 24860 9605 24869 9639
rect 24869 9605 24903 9639
rect 24903 9605 24912 9639
rect 24860 9596 24912 9605
rect 17500 9392 17552 9444
rect 19892 9503 19944 9512
rect 19892 9469 19901 9503
rect 19901 9469 19935 9503
rect 19935 9469 19944 9503
rect 19892 9460 19944 9469
rect 20168 9503 20220 9512
rect 9680 9324 9732 9376
rect 12440 9324 12492 9376
rect 13176 9324 13228 9376
rect 16028 9324 16080 9376
rect 17040 9324 17092 9376
rect 18052 9324 18104 9376
rect 20168 9469 20177 9503
rect 20177 9469 20211 9503
rect 20211 9469 20220 9503
rect 20168 9460 20220 9469
rect 21180 9460 21232 9512
rect 22100 9460 22152 9512
rect 22192 9392 22244 9444
rect 23388 9460 23440 9512
rect 23756 9460 23808 9512
rect 24952 9528 25004 9580
rect 24492 9503 24544 9512
rect 24492 9469 24501 9503
rect 24501 9469 24535 9503
rect 24535 9469 24544 9503
rect 24492 9460 24544 9469
rect 25228 9460 25280 9512
rect 23296 9392 23348 9444
rect 20444 9324 20496 9376
rect 21180 9324 21232 9376
rect 22284 9324 22336 9376
rect 22744 9324 22796 9376
rect 24492 9324 24544 9376
rect 24952 9324 25004 9376
rect 7114 9222 7166 9274
rect 7178 9222 7230 9274
rect 7242 9222 7294 9274
rect 7306 9222 7358 9274
rect 7370 9222 7422 9274
rect 13830 9222 13882 9274
rect 13894 9222 13946 9274
rect 13958 9222 14010 9274
rect 14022 9222 14074 9274
rect 14086 9222 14138 9274
rect 20546 9222 20598 9274
rect 20610 9222 20662 9274
rect 20674 9222 20726 9274
rect 20738 9222 20790 9274
rect 20802 9222 20854 9274
rect 27262 9222 27314 9274
rect 27326 9222 27378 9274
rect 27390 9222 27442 9274
rect 27454 9222 27506 9274
rect 27518 9222 27570 9274
rect 1676 9163 1728 9172
rect 1676 9129 1691 9163
rect 1691 9129 1725 9163
rect 1725 9129 1728 9163
rect 1676 9120 1728 9129
rect 2044 9120 2096 9172
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 8116 9163 8168 9172
rect 8116 9129 8125 9163
rect 8125 9129 8159 9163
rect 8159 9129 8168 9163
rect 8116 9120 8168 9129
rect 8300 9120 8352 9172
rect 8760 9120 8812 9172
rect 8852 9120 8904 9172
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 5172 9095 5224 9104
rect 5172 9061 5181 9095
rect 5181 9061 5215 9095
rect 5215 9061 5224 9095
rect 5172 9052 5224 9061
rect 8392 9095 8444 9104
rect 8392 9061 8401 9095
rect 8401 9061 8435 9095
rect 8435 9061 8444 9095
rect 8392 9052 8444 9061
rect 9312 9163 9364 9172
rect 9312 9129 9321 9163
rect 9321 9129 9355 9163
rect 9355 9129 9364 9163
rect 9312 9120 9364 9129
rect 11888 9163 11940 9172
rect 11888 9129 11897 9163
rect 11897 9129 11931 9163
rect 11931 9129 11940 9163
rect 11888 9120 11940 9129
rect 12164 9120 12216 9172
rect 14280 9120 14332 9172
rect 17776 9120 17828 9172
rect 2872 8984 2924 9036
rect 2044 8891 2096 8900
rect 2044 8857 2053 8891
rect 2053 8857 2087 8891
rect 2087 8857 2096 8891
rect 2044 8848 2096 8857
rect 2320 8916 2372 8968
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 5816 8984 5868 9036
rect 7012 9027 7064 9036
rect 7012 8993 7046 9027
rect 7046 8993 7064 9027
rect 7012 8984 7064 8993
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 8208 8916 8260 8968
rect 2228 8780 2280 8832
rect 4436 8780 4488 8832
rect 4804 8780 4856 8832
rect 7472 8780 7524 8832
rect 8760 8848 8812 8900
rect 8944 9027 8996 9036
rect 8944 8993 8953 9027
rect 8953 8993 8987 9027
rect 8987 8993 8996 9027
rect 8944 8984 8996 8993
rect 9772 9052 9824 9104
rect 10968 9052 11020 9104
rect 9312 8984 9364 9036
rect 11336 8984 11388 9036
rect 12348 8984 12400 9036
rect 11888 8916 11940 8968
rect 13268 9052 13320 9104
rect 13176 9027 13228 9036
rect 13176 8993 13185 9027
rect 13185 8993 13219 9027
rect 13219 8993 13228 9027
rect 13176 8984 13228 8993
rect 13544 9027 13596 9036
rect 13544 8993 13548 9027
rect 13548 8993 13582 9027
rect 13582 8993 13596 9027
rect 13544 8984 13596 8993
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 15476 9095 15528 9104
rect 15476 9061 15494 9095
rect 15494 9061 15528 9095
rect 15476 9052 15528 9061
rect 16764 9027 16816 9036
rect 16764 8993 16798 9027
rect 16798 8993 16816 9027
rect 13452 8916 13504 8968
rect 16764 8984 16816 8993
rect 18788 9120 18840 9172
rect 22376 9120 22428 9172
rect 18052 9052 18104 9104
rect 18788 9027 18840 9036
rect 18788 8993 18797 9027
rect 18797 8993 18831 9027
rect 18831 8993 18840 9027
rect 18788 8984 18840 8993
rect 19892 9052 19944 9104
rect 20076 8984 20128 9036
rect 20904 8984 20956 9036
rect 21732 9052 21784 9104
rect 14280 8916 14332 8968
rect 16304 8916 16356 8968
rect 9036 8848 9088 8900
rect 9404 8848 9456 8900
rect 10048 8848 10100 8900
rect 12348 8848 12400 8900
rect 22100 8984 22152 9036
rect 21640 8916 21692 8968
rect 23296 9027 23348 9036
rect 23296 8993 23305 9027
rect 23305 8993 23339 9027
rect 23339 8993 23348 9027
rect 23296 8984 23348 8993
rect 23388 9027 23440 9036
rect 23388 8993 23397 9027
rect 23397 8993 23431 9027
rect 23431 8993 23440 9027
rect 23388 8984 23440 8993
rect 23204 8916 23256 8968
rect 23296 8848 23348 8900
rect 23572 8848 23624 8900
rect 26424 9052 26476 9104
rect 23756 9027 23808 9036
rect 23756 8993 23765 9027
rect 23765 8993 23799 9027
rect 23799 8993 23808 9027
rect 23756 8984 23808 8993
rect 24308 8984 24360 9036
rect 25780 9027 25832 9036
rect 25780 8993 25789 9027
rect 25789 8993 25823 9027
rect 25823 8993 25832 9027
rect 25780 8984 25832 8993
rect 25412 8959 25464 8968
rect 25412 8925 25421 8959
rect 25421 8925 25455 8959
rect 25455 8925 25464 8959
rect 25412 8916 25464 8925
rect 25688 8916 25740 8968
rect 12256 8780 12308 8832
rect 17960 8823 18012 8832
rect 17960 8789 17969 8823
rect 17969 8789 18003 8823
rect 18003 8789 18012 8823
rect 17960 8780 18012 8789
rect 19524 8780 19576 8832
rect 21640 8780 21692 8832
rect 21916 8780 21968 8832
rect 23112 8823 23164 8832
rect 23112 8789 23121 8823
rect 23121 8789 23155 8823
rect 23155 8789 23164 8823
rect 23112 8780 23164 8789
rect 24400 8780 24452 8832
rect 25596 8848 25648 8900
rect 25504 8823 25556 8832
rect 25504 8789 25513 8823
rect 25513 8789 25547 8823
rect 25547 8789 25556 8823
rect 25504 8780 25556 8789
rect 3756 8678 3808 8730
rect 3820 8678 3872 8730
rect 3884 8678 3936 8730
rect 3948 8678 4000 8730
rect 4012 8678 4064 8730
rect 10472 8678 10524 8730
rect 10536 8678 10588 8730
rect 10600 8678 10652 8730
rect 10664 8678 10716 8730
rect 10728 8678 10780 8730
rect 17188 8678 17240 8730
rect 17252 8678 17304 8730
rect 17316 8678 17368 8730
rect 17380 8678 17432 8730
rect 17444 8678 17496 8730
rect 23904 8678 23956 8730
rect 23968 8678 24020 8730
rect 24032 8678 24084 8730
rect 24096 8678 24148 8730
rect 24160 8678 24212 8730
rect 3148 8576 3200 8628
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 8668 8576 8720 8628
rect 9036 8576 9088 8628
rect 10968 8576 11020 8628
rect 1492 8372 1544 8424
rect 2688 8372 2740 8424
rect 4344 8508 4396 8560
rect 8944 8508 8996 8560
rect 9588 8508 9640 8560
rect 9772 8508 9824 8560
rect 12624 8576 12676 8628
rect 13544 8576 13596 8628
rect 13636 8576 13688 8628
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 4436 8440 4488 8492
rect 9220 8440 9272 8492
rect 10416 8440 10468 8492
rect 2228 8304 2280 8356
rect 4068 8372 4120 8424
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 8484 8372 8536 8424
rect 8760 8372 8812 8424
rect 9312 8415 9364 8424
rect 9312 8381 9321 8415
rect 9321 8381 9355 8415
rect 9355 8381 9364 8415
rect 9312 8372 9364 8381
rect 9404 8415 9456 8424
rect 9404 8381 9414 8415
rect 9414 8381 9448 8415
rect 9448 8381 9456 8415
rect 9404 8372 9456 8381
rect 9588 8415 9640 8424
rect 9588 8381 9597 8415
rect 9597 8381 9631 8415
rect 9631 8381 9640 8415
rect 9588 8372 9640 8381
rect 9772 8415 9824 8424
rect 11336 8440 11388 8492
rect 9772 8381 9786 8415
rect 9786 8381 9820 8415
rect 9820 8381 9824 8415
rect 9772 8372 9824 8381
rect 11244 8415 11296 8424
rect 11244 8381 11254 8415
rect 11254 8381 11288 8415
rect 11288 8381 11296 8415
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 12532 8508 12584 8560
rect 11244 8372 11296 8381
rect 12164 8415 12216 8424
rect 12164 8381 12173 8415
rect 12173 8381 12207 8415
rect 12207 8381 12216 8415
rect 12164 8372 12216 8381
rect 4528 8304 4580 8356
rect 7012 8304 7064 8356
rect 8208 8304 8260 8356
rect 8576 8347 8628 8356
rect 8576 8313 8585 8347
rect 8585 8313 8619 8347
rect 8619 8313 8628 8347
rect 8576 8304 8628 8313
rect 3424 8279 3476 8288
rect 3424 8245 3433 8279
rect 3433 8245 3467 8279
rect 3467 8245 3476 8279
rect 3424 8236 3476 8245
rect 3608 8236 3660 8288
rect 4344 8279 4396 8288
rect 4344 8245 4353 8279
rect 4353 8245 4387 8279
rect 4387 8245 4396 8279
rect 4344 8236 4396 8245
rect 4436 8279 4488 8288
rect 4436 8245 4445 8279
rect 4445 8245 4479 8279
rect 4479 8245 4488 8279
rect 4436 8236 4488 8245
rect 7748 8279 7800 8288
rect 7748 8245 7757 8279
rect 7757 8245 7791 8279
rect 7791 8245 7800 8279
rect 7748 8236 7800 8245
rect 8852 8236 8904 8288
rect 10968 8304 11020 8356
rect 12072 8304 12124 8356
rect 12348 8415 12400 8424
rect 12348 8381 12357 8415
rect 12357 8381 12391 8415
rect 12391 8381 12400 8415
rect 12348 8372 12400 8381
rect 12532 8415 12584 8424
rect 12532 8381 12541 8415
rect 12541 8381 12575 8415
rect 12575 8381 12584 8415
rect 12532 8372 12584 8381
rect 10324 8236 10376 8288
rect 10416 8236 10468 8288
rect 12440 8304 12492 8356
rect 12992 8415 13044 8424
rect 12992 8381 13001 8415
rect 13001 8381 13035 8415
rect 13035 8381 13044 8415
rect 12992 8372 13044 8381
rect 14280 8372 14332 8424
rect 13084 8304 13136 8356
rect 16120 8576 16172 8628
rect 16764 8576 16816 8628
rect 19432 8576 19484 8628
rect 17776 8551 17828 8560
rect 17776 8517 17785 8551
rect 17785 8517 17819 8551
rect 17819 8517 17828 8551
rect 17776 8508 17828 8517
rect 22192 8619 22244 8628
rect 22192 8585 22201 8619
rect 22201 8585 22235 8619
rect 22235 8585 22244 8619
rect 22192 8576 22244 8585
rect 22284 8576 22336 8628
rect 23756 8576 23808 8628
rect 24308 8576 24360 8628
rect 16304 8483 16356 8492
rect 16304 8449 16313 8483
rect 16313 8449 16347 8483
rect 16347 8449 16356 8483
rect 16304 8440 16356 8449
rect 20904 8483 20956 8492
rect 20904 8449 20913 8483
rect 20913 8449 20947 8483
rect 20947 8449 20956 8483
rect 20904 8440 20956 8449
rect 21364 8440 21416 8492
rect 23112 8508 23164 8560
rect 23572 8508 23624 8560
rect 16028 8415 16080 8424
rect 16028 8381 16046 8415
rect 16046 8381 16080 8415
rect 16028 8372 16080 8381
rect 17040 8372 17092 8424
rect 17408 8415 17460 8424
rect 17408 8381 17417 8415
rect 17417 8381 17451 8415
rect 17451 8381 17460 8415
rect 17408 8372 17460 8381
rect 17592 8415 17644 8424
rect 17592 8381 17601 8415
rect 17601 8381 17635 8415
rect 17635 8381 17644 8415
rect 17592 8372 17644 8381
rect 19340 8372 19392 8424
rect 19524 8415 19576 8424
rect 19524 8381 19558 8415
rect 19558 8381 19576 8415
rect 19524 8372 19576 8381
rect 20996 8415 21048 8424
rect 20996 8381 21005 8415
rect 21005 8381 21039 8415
rect 21039 8381 21048 8415
rect 20996 8372 21048 8381
rect 17960 8304 18012 8356
rect 18052 8304 18104 8356
rect 21180 8304 21232 8356
rect 21456 8372 21508 8424
rect 21640 8372 21692 8424
rect 23848 8440 23900 8492
rect 24400 8440 24452 8492
rect 24952 8483 25004 8492
rect 24952 8449 24961 8483
rect 24961 8449 24995 8483
rect 24995 8449 25004 8483
rect 24952 8440 25004 8449
rect 25412 8576 25464 8628
rect 21916 8415 21968 8424
rect 21916 8381 21925 8415
rect 21925 8381 21959 8415
rect 21959 8381 21968 8415
rect 21916 8372 21968 8381
rect 22744 8347 22796 8356
rect 22744 8313 22753 8347
rect 22753 8313 22787 8347
rect 22787 8313 22796 8347
rect 22744 8304 22796 8313
rect 22836 8304 22888 8356
rect 23296 8304 23348 8356
rect 24124 8372 24176 8424
rect 25504 8304 25556 8356
rect 13268 8279 13320 8288
rect 13268 8245 13277 8279
rect 13277 8245 13311 8279
rect 13311 8245 13320 8279
rect 13268 8236 13320 8245
rect 20904 8236 20956 8288
rect 21824 8236 21876 8288
rect 23020 8236 23072 8288
rect 25688 8236 25740 8288
rect 26516 8279 26568 8288
rect 26516 8245 26525 8279
rect 26525 8245 26559 8279
rect 26559 8245 26568 8279
rect 26516 8236 26568 8245
rect 7114 8134 7166 8186
rect 7178 8134 7230 8186
rect 7242 8134 7294 8186
rect 7306 8134 7358 8186
rect 7370 8134 7422 8186
rect 13830 8134 13882 8186
rect 13894 8134 13946 8186
rect 13958 8134 14010 8186
rect 14022 8134 14074 8186
rect 14086 8134 14138 8186
rect 20546 8134 20598 8186
rect 20610 8134 20662 8186
rect 20674 8134 20726 8186
rect 20738 8134 20790 8186
rect 20802 8134 20854 8186
rect 27262 8134 27314 8186
rect 27326 8134 27378 8186
rect 27390 8134 27442 8186
rect 27454 8134 27506 8186
rect 27518 8134 27570 8186
rect 4068 8075 4120 8084
rect 4068 8041 4077 8075
rect 4077 8041 4111 8075
rect 4111 8041 4120 8075
rect 4068 8032 4120 8041
rect 7564 8032 7616 8084
rect 7748 8032 7800 8084
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 8576 8032 8628 8084
rect 2412 7939 2464 7948
rect 2412 7905 2421 7939
rect 2421 7905 2455 7939
rect 2455 7905 2464 7939
rect 2412 7896 2464 7905
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 10048 7964 10100 8016
rect 12532 8032 12584 8084
rect 20904 8032 20956 8084
rect 20996 8032 21048 8084
rect 6736 7896 6788 7948
rect 7288 7939 7340 7948
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 7380 7939 7432 7948
rect 7380 7905 7389 7939
rect 7389 7905 7423 7939
rect 7423 7905 7432 7939
rect 7380 7896 7432 7905
rect 6276 7828 6328 7880
rect 9036 7896 9088 7948
rect 9312 7896 9364 7948
rect 9496 7939 9548 7948
rect 9496 7905 9506 7939
rect 9506 7905 9540 7939
rect 9540 7905 9548 7939
rect 9496 7896 9548 7905
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 9864 7939 9916 7948
rect 9864 7905 9878 7939
rect 9878 7905 9912 7939
rect 9912 7905 9916 7939
rect 9864 7896 9916 7905
rect 10324 7939 10376 7948
rect 10324 7905 10333 7939
rect 10333 7905 10367 7939
rect 10367 7905 10376 7939
rect 10324 7896 10376 7905
rect 10416 7939 10468 7948
rect 10416 7905 10425 7939
rect 10425 7905 10459 7939
rect 10459 7905 10468 7939
rect 10416 7896 10468 7905
rect 13268 7964 13320 8016
rect 21732 8075 21784 8084
rect 21732 8041 21741 8075
rect 21741 8041 21775 8075
rect 21775 8041 21784 8075
rect 21732 8032 21784 8041
rect 21824 8032 21876 8084
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 8760 7871 8812 7880
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 11244 7828 11296 7880
rect 12164 7828 12216 7880
rect 5908 7760 5960 7812
rect 6828 7735 6880 7744
rect 6828 7701 6837 7735
rect 6837 7701 6871 7735
rect 6871 7701 6880 7735
rect 6828 7692 6880 7701
rect 7840 7760 7892 7812
rect 8576 7760 8628 7812
rect 9864 7760 9916 7812
rect 12348 7939 12400 7948
rect 12348 7905 12360 7939
rect 12360 7905 12394 7939
rect 12394 7905 12400 7939
rect 12348 7896 12400 7905
rect 12716 7896 12768 7948
rect 21180 7896 21232 7948
rect 21364 7939 21416 7948
rect 21364 7905 21373 7939
rect 21373 7905 21407 7939
rect 21407 7905 21416 7939
rect 21364 7896 21416 7905
rect 21824 7896 21876 7948
rect 12348 7760 12400 7812
rect 13820 7828 13872 7880
rect 21456 7828 21508 7880
rect 22376 7964 22428 8016
rect 22652 7964 22704 8016
rect 23756 7964 23808 8016
rect 22836 7896 22888 7948
rect 23020 7939 23072 7948
rect 23020 7905 23029 7939
rect 23029 7905 23063 7939
rect 23063 7905 23072 7939
rect 23020 7896 23072 7905
rect 23204 7939 23256 7948
rect 23204 7905 23213 7939
rect 23213 7905 23247 7939
rect 23247 7905 23256 7939
rect 23204 7896 23256 7905
rect 23296 7939 23348 7948
rect 23296 7905 23305 7939
rect 23305 7905 23339 7939
rect 23339 7905 23348 7939
rect 23296 7896 23348 7905
rect 23480 7939 23532 7948
rect 23480 7905 23489 7939
rect 23489 7905 23523 7939
rect 23523 7905 23532 7939
rect 23480 7896 23532 7905
rect 24124 7939 24176 7948
rect 24124 7905 24133 7939
rect 24133 7905 24167 7939
rect 24167 7905 24176 7939
rect 24124 7896 24176 7905
rect 23572 7828 23624 7880
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 24952 8032 25004 8084
rect 26424 8075 26476 8084
rect 26424 8041 26433 8075
rect 26433 8041 26467 8075
rect 26467 8041 26476 8075
rect 26424 8032 26476 8041
rect 25412 7964 25464 8016
rect 25504 7896 25556 7948
rect 26516 7896 26568 7948
rect 17408 7760 17460 7812
rect 8944 7692 8996 7744
rect 11336 7692 11388 7744
rect 13820 7692 13872 7744
rect 14280 7692 14332 7744
rect 15384 7692 15436 7744
rect 19340 7692 19392 7744
rect 19892 7735 19944 7744
rect 19892 7701 19901 7735
rect 19901 7701 19935 7735
rect 19935 7701 19944 7735
rect 19892 7692 19944 7701
rect 20076 7803 20128 7812
rect 20076 7769 20085 7803
rect 20085 7769 20119 7803
rect 20119 7769 20128 7803
rect 20076 7760 20128 7769
rect 22284 7760 22336 7812
rect 22192 7735 22244 7744
rect 22192 7701 22201 7735
rect 22201 7701 22235 7735
rect 22235 7701 22244 7735
rect 22192 7692 22244 7701
rect 22376 7692 22428 7744
rect 24584 7735 24636 7744
rect 24584 7701 24593 7735
rect 24593 7701 24627 7735
rect 24627 7701 24636 7735
rect 24584 7692 24636 7701
rect 25320 7692 25372 7744
rect 3756 7590 3808 7642
rect 3820 7590 3872 7642
rect 3884 7590 3936 7642
rect 3948 7590 4000 7642
rect 4012 7590 4064 7642
rect 10472 7590 10524 7642
rect 10536 7590 10588 7642
rect 10600 7590 10652 7642
rect 10664 7590 10716 7642
rect 10728 7590 10780 7642
rect 17188 7590 17240 7642
rect 17252 7590 17304 7642
rect 17316 7590 17368 7642
rect 17380 7590 17432 7642
rect 17444 7590 17496 7642
rect 23904 7590 23956 7642
rect 23968 7590 24020 7642
rect 24032 7590 24084 7642
rect 24096 7590 24148 7642
rect 24160 7590 24212 7642
rect 2412 7488 2464 7540
rect 3516 7488 3568 7540
rect 5908 7531 5960 7540
rect 5908 7497 5917 7531
rect 5917 7497 5951 7531
rect 5951 7497 5960 7531
rect 5908 7488 5960 7497
rect 6736 7488 6788 7540
rect 3332 7420 3384 7472
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 11244 7488 11296 7540
rect 3608 7352 3660 7404
rect 3516 7284 3568 7336
rect 5448 7352 5500 7404
rect 4160 7327 4212 7336
rect 4160 7293 4169 7327
rect 4169 7293 4203 7327
rect 4203 7293 4212 7327
rect 4160 7284 4212 7293
rect 3424 7259 3476 7268
rect 3424 7225 3433 7259
rect 3433 7225 3467 7259
rect 3467 7225 3476 7259
rect 3424 7216 3476 7225
rect 4436 7327 4488 7336
rect 4436 7293 4445 7327
rect 4445 7293 4479 7327
rect 4479 7293 4488 7327
rect 4436 7284 4488 7293
rect 4528 7327 4580 7336
rect 4528 7293 4537 7327
rect 4537 7293 4571 7327
rect 4571 7293 4580 7327
rect 4528 7284 4580 7293
rect 5356 7284 5408 7336
rect 5724 7327 5776 7336
rect 5724 7293 5733 7327
rect 5733 7293 5767 7327
rect 5767 7293 5776 7327
rect 6184 7327 6236 7336
rect 5724 7284 5776 7293
rect 6184 7293 6193 7327
rect 6193 7293 6227 7327
rect 6227 7293 6236 7327
rect 6184 7284 6236 7293
rect 6552 7327 6604 7336
rect 6552 7293 6561 7327
rect 6561 7293 6595 7327
rect 6595 7293 6604 7327
rect 6552 7284 6604 7293
rect 6828 7327 6880 7336
rect 6828 7293 6862 7327
rect 6862 7293 6880 7327
rect 6828 7284 6880 7293
rect 8392 7352 8444 7404
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 10968 7284 11020 7336
rect 12348 7284 12400 7336
rect 13820 7327 13872 7336
rect 13820 7293 13854 7327
rect 13854 7293 13872 7327
rect 13820 7284 13872 7293
rect 15200 7488 15252 7540
rect 15936 7531 15988 7540
rect 15936 7497 15945 7531
rect 15945 7497 15979 7531
rect 15979 7497 15988 7531
rect 15936 7488 15988 7497
rect 18788 7488 18840 7540
rect 19892 7488 19944 7540
rect 23020 7488 23072 7540
rect 23480 7488 23532 7540
rect 10876 7216 10928 7268
rect 11336 7259 11388 7268
rect 11336 7225 11370 7259
rect 11370 7225 11388 7259
rect 11336 7216 11388 7225
rect 16028 7284 16080 7336
rect 16304 7352 16356 7404
rect 20260 7352 20312 7404
rect 25504 7488 25556 7540
rect 25780 7420 25832 7472
rect 18696 7284 18748 7336
rect 4344 7191 4396 7200
rect 4344 7157 4353 7191
rect 4353 7157 4387 7191
rect 4387 7157 4396 7191
rect 4344 7148 4396 7157
rect 4804 7148 4856 7200
rect 5264 7148 5316 7200
rect 8300 7148 8352 7200
rect 11428 7148 11480 7200
rect 12164 7148 12216 7200
rect 12808 7148 12860 7200
rect 18880 7327 18932 7336
rect 18880 7293 18889 7327
rect 18889 7293 18923 7327
rect 18923 7293 18932 7327
rect 18880 7284 18932 7293
rect 19340 7284 19392 7336
rect 21456 7327 21508 7336
rect 21456 7293 21465 7327
rect 21465 7293 21499 7327
rect 21499 7293 21508 7327
rect 21456 7284 21508 7293
rect 21732 7327 21784 7336
rect 21732 7293 21741 7327
rect 21741 7293 21775 7327
rect 21775 7293 21784 7327
rect 21732 7284 21784 7293
rect 24584 7284 24636 7336
rect 25320 7327 25372 7336
rect 25320 7293 25329 7327
rect 25329 7293 25363 7327
rect 25363 7293 25372 7327
rect 25320 7284 25372 7293
rect 18604 7148 18656 7200
rect 23388 7259 23440 7268
rect 23388 7225 23397 7259
rect 23397 7225 23431 7259
rect 23431 7225 23440 7259
rect 23388 7216 23440 7225
rect 23756 7216 23808 7268
rect 25780 7327 25832 7336
rect 25780 7293 25789 7327
rect 25789 7293 25823 7327
rect 25823 7293 25832 7327
rect 25780 7284 25832 7293
rect 19524 7148 19576 7200
rect 19708 7148 19760 7200
rect 22100 7148 22152 7200
rect 25688 7191 25740 7200
rect 25688 7157 25697 7191
rect 25697 7157 25731 7191
rect 25731 7157 25740 7191
rect 25688 7148 25740 7157
rect 7114 7046 7166 7098
rect 7178 7046 7230 7098
rect 7242 7046 7294 7098
rect 7306 7046 7358 7098
rect 7370 7046 7422 7098
rect 13830 7046 13882 7098
rect 13894 7046 13946 7098
rect 13958 7046 14010 7098
rect 14022 7046 14074 7098
rect 14086 7046 14138 7098
rect 20546 7046 20598 7098
rect 20610 7046 20662 7098
rect 20674 7046 20726 7098
rect 20738 7046 20790 7098
rect 20802 7046 20854 7098
rect 27262 7046 27314 7098
rect 27326 7046 27378 7098
rect 27390 7046 27442 7098
rect 27454 7046 27506 7098
rect 27518 7046 27570 7098
rect 3608 6944 3660 6996
rect 4252 6944 4304 6996
rect 5356 6987 5408 6996
rect 5356 6953 5365 6987
rect 5365 6953 5399 6987
rect 5399 6953 5408 6987
rect 5356 6944 5408 6953
rect 5448 6987 5500 6996
rect 5448 6953 5457 6987
rect 5457 6953 5491 6987
rect 5491 6953 5500 6987
rect 5448 6944 5500 6953
rect 8760 6944 8812 6996
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 2044 6808 2096 6860
rect 2320 6808 2372 6860
rect 3516 6808 3568 6860
rect 4804 6808 4856 6860
rect 8116 6876 8168 6928
rect 9496 6876 9548 6928
rect 8300 6808 8352 6860
rect 2596 6672 2648 6724
rect 6552 6740 6604 6792
rect 7472 6783 7524 6792
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 8484 6740 8536 6792
rect 3056 6604 3108 6656
rect 5356 6672 5408 6724
rect 6276 6672 6328 6724
rect 4252 6647 4304 6656
rect 4252 6613 4261 6647
rect 4261 6613 4295 6647
rect 4295 6613 4304 6647
rect 4252 6604 4304 6613
rect 4436 6604 4488 6656
rect 5724 6604 5776 6656
rect 6184 6604 6236 6656
rect 11428 6851 11480 6860
rect 11428 6817 11437 6851
rect 11437 6817 11471 6851
rect 11471 6817 11480 6851
rect 11428 6808 11480 6817
rect 11060 6740 11112 6792
rect 12072 6851 12124 6860
rect 12072 6817 12081 6851
rect 12081 6817 12115 6851
rect 12115 6817 12124 6851
rect 12072 6808 12124 6817
rect 12256 6808 12308 6860
rect 14096 6808 14148 6860
rect 14556 6808 14608 6860
rect 14740 6851 14792 6860
rect 14740 6817 14749 6851
rect 14749 6817 14783 6851
rect 14783 6817 14792 6851
rect 14740 6808 14792 6817
rect 18880 6944 18932 6996
rect 23204 6987 23256 6996
rect 23204 6953 23213 6987
rect 23213 6953 23247 6987
rect 23247 6953 23256 6987
rect 23204 6944 23256 6953
rect 23756 6944 23808 6996
rect 15568 6851 15620 6860
rect 15568 6817 15577 6851
rect 15577 6817 15611 6851
rect 15611 6817 15620 6851
rect 15568 6808 15620 6817
rect 10232 6672 10284 6724
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 18788 6876 18840 6928
rect 20720 6876 20772 6928
rect 21732 6876 21784 6928
rect 22100 6919 22152 6928
rect 22100 6885 22134 6919
rect 22134 6885 22152 6919
rect 22100 6876 22152 6885
rect 23664 6876 23716 6928
rect 24400 6944 24452 6996
rect 25780 6987 25832 6996
rect 25780 6953 25789 6987
rect 25789 6953 25823 6987
rect 25823 6953 25832 6987
rect 25780 6944 25832 6953
rect 18512 6808 18564 6860
rect 25228 6876 25280 6928
rect 20260 6808 20312 6860
rect 18604 6783 18656 6792
rect 18604 6749 18613 6783
rect 18613 6749 18647 6783
rect 18647 6749 18656 6783
rect 18604 6740 18656 6749
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 20444 6851 20496 6860
rect 20444 6817 20453 6851
rect 20453 6817 20487 6851
rect 20487 6817 20496 6851
rect 20444 6808 20496 6817
rect 20536 6808 20588 6860
rect 20720 6740 20772 6792
rect 23020 6808 23072 6860
rect 24492 6808 24544 6860
rect 24768 6808 24820 6860
rect 25596 6808 25648 6860
rect 11336 6604 11388 6656
rect 11428 6604 11480 6656
rect 14280 6604 14332 6656
rect 15568 6604 15620 6656
rect 16028 6604 16080 6656
rect 17960 6604 18012 6656
rect 19340 6672 19392 6724
rect 19708 6604 19760 6656
rect 20076 6647 20128 6656
rect 20076 6613 20085 6647
rect 20085 6613 20119 6647
rect 20119 6613 20128 6647
rect 20076 6604 20128 6613
rect 20444 6604 20496 6656
rect 24676 6740 24728 6792
rect 25136 6783 25188 6792
rect 25136 6749 25145 6783
rect 25145 6749 25179 6783
rect 25179 6749 25188 6783
rect 25136 6740 25188 6749
rect 25872 6740 25924 6792
rect 23388 6672 23440 6724
rect 24952 6604 25004 6656
rect 3756 6502 3808 6554
rect 3820 6502 3872 6554
rect 3884 6502 3936 6554
rect 3948 6502 4000 6554
rect 4012 6502 4064 6554
rect 10472 6502 10524 6554
rect 10536 6502 10588 6554
rect 10600 6502 10652 6554
rect 10664 6502 10716 6554
rect 10728 6502 10780 6554
rect 17188 6502 17240 6554
rect 17252 6502 17304 6554
rect 17316 6502 17368 6554
rect 17380 6502 17432 6554
rect 17444 6502 17496 6554
rect 23904 6502 23956 6554
rect 23968 6502 24020 6554
rect 24032 6502 24084 6554
rect 24096 6502 24148 6554
rect 24160 6502 24212 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 2872 6400 2924 6452
rect 3608 6400 3660 6452
rect 4804 6443 4856 6452
rect 4804 6409 4813 6443
rect 4813 6409 4847 6443
rect 4847 6409 4856 6443
rect 4804 6400 4856 6409
rect 6276 6443 6328 6452
rect 6276 6409 6285 6443
rect 6285 6409 6319 6443
rect 6319 6409 6328 6443
rect 6276 6400 6328 6409
rect 9036 6400 9088 6452
rect 10232 6332 10284 6384
rect 11336 6375 11388 6384
rect 11336 6341 11345 6375
rect 11345 6341 11379 6375
rect 11379 6341 11388 6375
rect 11336 6332 11388 6341
rect 11612 6400 11664 6452
rect 14464 6400 14516 6452
rect 18696 6400 18748 6452
rect 21456 6400 21508 6452
rect 22192 6443 22244 6452
rect 22192 6409 22201 6443
rect 22201 6409 22235 6443
rect 22235 6409 22244 6443
rect 22192 6400 22244 6409
rect 24676 6400 24728 6452
rect 24952 6443 25004 6452
rect 24952 6409 24961 6443
rect 24961 6409 24995 6443
rect 24995 6409 25004 6443
rect 24952 6400 25004 6409
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 2688 6264 2740 6316
rect 2596 6239 2648 6248
rect 2596 6205 2605 6239
rect 2605 6205 2639 6239
rect 2639 6205 2648 6239
rect 2596 6196 2648 6205
rect 2872 6239 2924 6248
rect 2872 6205 2881 6239
rect 2881 6205 2915 6239
rect 2915 6205 2924 6239
rect 2872 6196 2924 6205
rect 3056 6239 3108 6248
rect 3056 6205 3065 6239
rect 3065 6205 3099 6239
rect 3099 6205 3108 6239
rect 3056 6196 3108 6205
rect 10876 6264 10928 6316
rect 11060 6264 11112 6316
rect 5540 6196 5592 6248
rect 6552 6196 6604 6248
rect 7472 6196 7524 6248
rect 10232 6239 10284 6248
rect 10232 6205 10241 6239
rect 10241 6205 10275 6239
rect 10275 6205 10284 6239
rect 10232 6196 10284 6205
rect 3332 6128 3384 6180
rect 4344 6128 4396 6180
rect 5172 6171 5224 6180
rect 5172 6137 5206 6171
rect 5206 6137 5224 6171
rect 5172 6128 5224 6137
rect 6368 6171 6420 6180
rect 6368 6137 6377 6171
rect 6377 6137 6411 6171
rect 6411 6137 6420 6171
rect 6368 6128 6420 6137
rect 8668 6171 8720 6180
rect 8668 6137 8702 6171
rect 8702 6137 8720 6171
rect 8668 6128 8720 6137
rect 4528 6060 4580 6112
rect 9036 6060 9088 6112
rect 9128 6060 9180 6112
rect 10232 6060 10284 6112
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 10600 6239 10652 6248
rect 10600 6205 10609 6239
rect 10609 6205 10643 6239
rect 10643 6205 10652 6239
rect 10600 6196 10652 6205
rect 10876 6171 10928 6180
rect 10876 6137 10885 6171
rect 10885 6137 10919 6171
rect 10919 6137 10928 6171
rect 10876 6128 10928 6137
rect 11428 6239 11480 6248
rect 11428 6205 11436 6239
rect 11436 6205 11470 6239
rect 11470 6205 11480 6239
rect 13084 6332 13136 6384
rect 15844 6375 15896 6384
rect 15844 6341 15853 6375
rect 15853 6341 15887 6375
rect 15887 6341 15896 6375
rect 15844 6332 15896 6341
rect 19524 6332 19576 6384
rect 19708 6332 19760 6384
rect 23020 6375 23072 6384
rect 23020 6341 23029 6375
rect 23029 6341 23063 6375
rect 23063 6341 23072 6375
rect 23020 6332 23072 6341
rect 23388 6332 23440 6384
rect 25412 6400 25464 6452
rect 25872 6400 25924 6452
rect 16304 6264 16356 6316
rect 11428 6196 11480 6205
rect 11888 6196 11940 6248
rect 12992 6196 13044 6248
rect 14096 6196 14148 6248
rect 16396 6196 16448 6248
rect 11244 6060 11296 6112
rect 14924 6128 14976 6180
rect 11980 6060 12032 6112
rect 13544 6060 13596 6112
rect 15292 6060 15344 6112
rect 16028 6103 16080 6112
rect 16028 6069 16037 6103
rect 16037 6069 16071 6103
rect 16071 6069 16080 6103
rect 16028 6060 16080 6069
rect 16488 6060 16540 6112
rect 17040 6239 17092 6248
rect 17040 6205 17049 6239
rect 17049 6205 17083 6239
rect 17083 6205 17092 6239
rect 17040 6196 17092 6205
rect 18512 6264 18564 6316
rect 19340 6264 19392 6316
rect 17960 6196 18012 6248
rect 19248 6196 19300 6248
rect 20628 6196 20680 6248
rect 20720 6239 20772 6248
rect 20720 6205 20729 6239
rect 20729 6205 20763 6239
rect 20763 6205 20772 6239
rect 20720 6196 20772 6205
rect 18880 6128 18932 6180
rect 20536 6171 20588 6180
rect 20536 6137 20545 6171
rect 20545 6137 20579 6171
rect 20579 6137 20588 6171
rect 20536 6128 20588 6137
rect 18052 6060 18104 6112
rect 20352 6060 20404 6112
rect 21088 6128 21140 6180
rect 23572 6264 23624 6316
rect 24400 6307 24452 6316
rect 24400 6273 24409 6307
rect 24409 6273 24443 6307
rect 24443 6273 24452 6307
rect 24400 6264 24452 6273
rect 22284 6128 22336 6180
rect 22376 6171 22428 6180
rect 22376 6137 22385 6171
rect 22385 6137 22419 6171
rect 22419 6137 22428 6171
rect 22376 6128 22428 6137
rect 25688 6196 25740 6248
rect 24768 6171 24820 6180
rect 24768 6137 24793 6171
rect 24793 6137 24820 6171
rect 24768 6128 24820 6137
rect 21456 6060 21508 6112
rect 22560 6060 22612 6112
rect 7114 5958 7166 6010
rect 7178 5958 7230 6010
rect 7242 5958 7294 6010
rect 7306 5958 7358 6010
rect 7370 5958 7422 6010
rect 13830 5958 13882 6010
rect 13894 5958 13946 6010
rect 13958 5958 14010 6010
rect 14022 5958 14074 6010
rect 14086 5958 14138 6010
rect 20546 5958 20598 6010
rect 20610 5958 20662 6010
rect 20674 5958 20726 6010
rect 20738 5958 20790 6010
rect 20802 5958 20854 6010
rect 27262 5958 27314 6010
rect 27326 5958 27378 6010
rect 27390 5958 27442 6010
rect 27454 5958 27506 6010
rect 27518 5958 27570 6010
rect 4252 5720 4304 5772
rect 3516 5652 3568 5704
rect 8484 5856 8536 5908
rect 8668 5899 8720 5908
rect 8668 5865 8677 5899
rect 8677 5865 8711 5899
rect 8711 5865 8720 5899
rect 8668 5856 8720 5865
rect 10416 5856 10468 5908
rect 5724 5788 5776 5840
rect 14004 5856 14056 5908
rect 14464 5856 14516 5908
rect 14924 5899 14976 5908
rect 14924 5865 14933 5899
rect 14933 5865 14967 5899
rect 14967 5865 14976 5899
rect 14924 5856 14976 5865
rect 17040 5856 17092 5908
rect 18052 5856 18104 5908
rect 18880 5856 18932 5908
rect 20352 5856 20404 5908
rect 6276 5720 6328 5772
rect 8576 5720 8628 5772
rect 8852 5720 8904 5772
rect 9128 5763 9180 5772
rect 9128 5729 9137 5763
rect 9137 5729 9171 5763
rect 9171 5729 9180 5763
rect 9128 5720 9180 5729
rect 10968 5763 11020 5772
rect 10968 5729 10977 5763
rect 10977 5729 11011 5763
rect 11011 5729 11020 5763
rect 10968 5720 11020 5729
rect 11060 5720 11112 5772
rect 11612 5720 11664 5772
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 10876 5652 10928 5704
rect 10784 5584 10836 5636
rect 12532 5652 12584 5704
rect 14556 5788 14608 5840
rect 14004 5763 14056 5772
rect 14004 5729 14013 5763
rect 14013 5729 14047 5763
rect 14047 5729 14056 5763
rect 14004 5720 14056 5729
rect 14188 5763 14240 5772
rect 14188 5729 14197 5763
rect 14197 5729 14231 5763
rect 14231 5729 14240 5763
rect 14188 5720 14240 5729
rect 14280 5720 14332 5772
rect 14464 5720 14516 5772
rect 16580 5788 16632 5840
rect 17500 5788 17552 5840
rect 15844 5720 15896 5772
rect 20076 5788 20128 5840
rect 20628 5788 20680 5840
rect 22100 5856 22152 5908
rect 22376 5856 22428 5908
rect 23296 5856 23348 5908
rect 23664 5856 23716 5908
rect 24400 5856 24452 5908
rect 25136 5856 25188 5908
rect 23388 5788 23440 5840
rect 25412 5788 25464 5840
rect 18696 5763 18748 5772
rect 12440 5627 12492 5636
rect 12440 5593 12449 5627
rect 12449 5593 12483 5627
rect 12483 5593 12492 5627
rect 12440 5584 12492 5593
rect 17316 5695 17368 5704
rect 17316 5661 17325 5695
rect 17325 5661 17359 5695
rect 17359 5661 17368 5695
rect 17316 5652 17368 5661
rect 18696 5729 18705 5763
rect 18705 5729 18739 5763
rect 18739 5729 18748 5763
rect 18696 5720 18748 5729
rect 19248 5720 19300 5772
rect 18512 5652 18564 5704
rect 17592 5584 17644 5636
rect 18788 5584 18840 5636
rect 5172 5516 5224 5568
rect 9036 5516 9088 5568
rect 14464 5516 14516 5568
rect 15936 5516 15988 5568
rect 17316 5516 17368 5568
rect 21088 5584 21140 5636
rect 22376 5763 22428 5772
rect 22376 5729 22385 5763
rect 22385 5729 22419 5763
rect 22419 5729 22428 5763
rect 22376 5720 22428 5729
rect 22560 5763 22612 5772
rect 22560 5729 22569 5763
rect 22569 5729 22603 5763
rect 22603 5729 22612 5763
rect 22560 5720 22612 5729
rect 22652 5763 22704 5772
rect 22652 5729 22661 5763
rect 22661 5729 22695 5763
rect 22695 5729 22704 5763
rect 22652 5720 22704 5729
rect 24492 5763 24544 5772
rect 24492 5729 24501 5763
rect 24501 5729 24535 5763
rect 24535 5729 24544 5763
rect 24492 5720 24544 5729
rect 25688 5763 25740 5772
rect 25688 5729 25706 5763
rect 25706 5729 25740 5763
rect 25688 5720 25740 5729
rect 20996 5516 21048 5568
rect 21456 5559 21508 5568
rect 21456 5525 21465 5559
rect 21465 5525 21499 5559
rect 21499 5525 21508 5559
rect 21456 5516 21508 5525
rect 24308 5516 24360 5568
rect 3756 5414 3808 5466
rect 3820 5414 3872 5466
rect 3884 5414 3936 5466
rect 3948 5414 4000 5466
rect 4012 5414 4064 5466
rect 10472 5414 10524 5466
rect 10536 5414 10588 5466
rect 10600 5414 10652 5466
rect 10664 5414 10716 5466
rect 10728 5414 10780 5466
rect 17188 5414 17240 5466
rect 17252 5414 17304 5466
rect 17316 5414 17368 5466
rect 17380 5414 17432 5466
rect 17444 5414 17496 5466
rect 23904 5414 23956 5466
rect 23968 5414 24020 5466
rect 24032 5414 24084 5466
rect 24096 5414 24148 5466
rect 24160 5414 24212 5466
rect 4068 5312 4120 5364
rect 5632 5312 5684 5364
rect 7196 5312 7248 5364
rect 7472 5312 7524 5364
rect 9956 5312 10008 5364
rect 10968 5312 11020 5364
rect 11796 5312 11848 5364
rect 13544 5355 13596 5364
rect 13544 5321 13553 5355
rect 13553 5321 13587 5355
rect 13587 5321 13596 5355
rect 13544 5312 13596 5321
rect 14648 5312 14700 5364
rect 15108 5312 15160 5364
rect 7656 5244 7708 5296
rect 5356 5176 5408 5228
rect 9128 5176 9180 5228
rect 5540 5108 5592 5160
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 5908 5108 5960 5117
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 7196 5151 7248 5160
rect 7196 5117 7205 5151
rect 7205 5117 7239 5151
rect 7239 5117 7248 5151
rect 7196 5108 7248 5117
rect 8024 5108 8076 5160
rect 8300 5108 8352 5160
rect 8760 5108 8812 5160
rect 8852 5151 8904 5160
rect 8852 5117 8861 5151
rect 8861 5117 8895 5151
rect 8895 5117 8904 5151
rect 8852 5108 8904 5117
rect 9036 5040 9088 5092
rect 9312 5151 9364 5160
rect 9312 5117 9321 5151
rect 9321 5117 9355 5151
rect 9355 5117 9364 5151
rect 9312 5108 9364 5117
rect 9404 5108 9456 5160
rect 10876 5244 10928 5296
rect 11152 5244 11204 5296
rect 15384 5244 15436 5296
rect 15568 5244 15620 5296
rect 10600 5176 10652 5228
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 14648 5176 14700 5228
rect 9680 5040 9732 5092
rect 11428 5151 11480 5160
rect 11428 5117 11437 5151
rect 11437 5117 11471 5151
rect 11471 5117 11480 5151
rect 11428 5108 11480 5117
rect 11520 5108 11572 5160
rect 12164 5108 12216 5160
rect 12808 5108 12860 5160
rect 15384 5108 15436 5160
rect 15476 5151 15528 5160
rect 15476 5117 15485 5151
rect 15485 5117 15519 5151
rect 15519 5117 15528 5151
rect 15476 5108 15528 5117
rect 14832 5083 14884 5092
rect 14832 5049 14841 5083
rect 14841 5049 14875 5083
rect 14875 5049 14884 5083
rect 14832 5040 14884 5049
rect 15936 5108 15988 5160
rect 16120 5151 16172 5160
rect 16120 5117 16129 5151
rect 16129 5117 16163 5151
rect 16163 5117 16172 5151
rect 16120 5108 16172 5117
rect 20260 5312 20312 5364
rect 16856 5244 16908 5296
rect 18788 5244 18840 5296
rect 22468 5312 22520 5364
rect 24952 5312 25004 5364
rect 25688 5312 25740 5364
rect 5908 4972 5960 5024
rect 6920 4972 6972 5024
rect 8208 4972 8260 5024
rect 9404 4972 9456 5024
rect 10324 4972 10376 5024
rect 12624 4972 12676 5024
rect 12992 5015 13044 5024
rect 12992 4981 13001 5015
rect 13001 4981 13035 5015
rect 13035 4981 13044 5015
rect 12992 4972 13044 4981
rect 13084 4972 13136 5024
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 19432 5176 19484 5228
rect 22652 5176 22704 5228
rect 18788 5151 18840 5160
rect 18788 5117 18797 5151
rect 18797 5117 18831 5151
rect 18831 5117 18840 5151
rect 18788 5108 18840 5117
rect 18880 5151 18932 5160
rect 18880 5117 18889 5151
rect 18889 5117 18923 5151
rect 18923 5117 18932 5151
rect 18880 5108 18932 5117
rect 20628 5108 20680 5160
rect 20996 5151 21048 5160
rect 20996 5117 21014 5151
rect 21014 5117 21048 5151
rect 20996 5108 21048 5117
rect 22376 5151 22428 5160
rect 22376 5117 22385 5151
rect 22385 5117 22419 5151
rect 22419 5117 22428 5151
rect 22376 5108 22428 5117
rect 23020 5151 23072 5160
rect 23020 5117 23029 5151
rect 23029 5117 23063 5151
rect 23063 5117 23072 5151
rect 23020 5108 23072 5117
rect 18604 5040 18656 5092
rect 19340 5040 19392 5092
rect 17132 5015 17184 5024
rect 17132 4981 17141 5015
rect 17141 4981 17175 5015
rect 17175 4981 17184 5015
rect 17132 4972 17184 4981
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 23388 5176 23440 5228
rect 23664 5108 23716 5160
rect 25228 5176 25280 5228
rect 24032 5151 24084 5160
rect 24032 5117 24041 5151
rect 24041 5117 24075 5151
rect 24075 5117 24084 5151
rect 24032 5108 24084 5117
rect 24308 5151 24360 5160
rect 24308 5117 24317 5151
rect 24317 5117 24351 5151
rect 24351 5117 24360 5151
rect 24308 5108 24360 5117
rect 24492 5151 24544 5160
rect 24492 5117 24501 5151
rect 24501 5117 24535 5151
rect 24535 5117 24544 5151
rect 24492 5108 24544 5117
rect 23296 5083 23348 5092
rect 23296 5049 23305 5083
rect 23305 5049 23339 5083
rect 23339 5049 23348 5083
rect 23296 5040 23348 5049
rect 23388 4972 23440 5024
rect 23664 5015 23716 5024
rect 23664 4981 23673 5015
rect 23673 4981 23707 5015
rect 23707 4981 23716 5015
rect 23664 4972 23716 4981
rect 7114 4870 7166 4922
rect 7178 4870 7230 4922
rect 7242 4870 7294 4922
rect 7306 4870 7358 4922
rect 7370 4870 7422 4922
rect 13830 4870 13882 4922
rect 13894 4870 13946 4922
rect 13958 4870 14010 4922
rect 14022 4870 14074 4922
rect 14086 4870 14138 4922
rect 20546 4870 20598 4922
rect 20610 4870 20662 4922
rect 20674 4870 20726 4922
rect 20738 4870 20790 4922
rect 20802 4870 20854 4922
rect 27262 4870 27314 4922
rect 27326 4870 27378 4922
rect 27390 4870 27442 4922
rect 27454 4870 27506 4922
rect 27518 4870 27570 4922
rect 6920 4768 6972 4820
rect 3424 4471 3476 4480
rect 3424 4437 3433 4471
rect 3433 4437 3467 4471
rect 3467 4437 3476 4471
rect 3424 4428 3476 4437
rect 4068 4675 4120 4684
rect 4068 4641 4077 4675
rect 4077 4641 4111 4675
rect 4111 4641 4120 4675
rect 4068 4632 4120 4641
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 5908 4700 5960 4752
rect 7656 4700 7708 4752
rect 5356 4675 5408 4684
rect 5356 4641 5365 4675
rect 5365 4641 5399 4675
rect 5399 4641 5408 4675
rect 5356 4632 5408 4641
rect 5632 4632 5684 4684
rect 5448 4564 5500 4616
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 7104 4675 7156 4684
rect 7104 4641 7113 4675
rect 7113 4641 7147 4675
rect 7147 4641 7156 4675
rect 7104 4632 7156 4641
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 7564 4675 7616 4684
rect 7564 4641 7573 4675
rect 7573 4641 7607 4675
rect 7607 4641 7616 4675
rect 7564 4632 7616 4641
rect 8300 4768 8352 4820
rect 8024 4700 8076 4752
rect 8208 4675 8260 4684
rect 8208 4641 8217 4675
rect 8217 4641 8251 4675
rect 8251 4641 8260 4675
rect 8208 4632 8260 4641
rect 8300 4632 8352 4684
rect 8576 4675 8628 4684
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 8576 4632 8628 4641
rect 8760 4768 8812 4820
rect 9220 4768 9272 4820
rect 9588 4768 9640 4820
rect 10140 4768 10192 4820
rect 10784 4768 10836 4820
rect 11520 4768 11572 4820
rect 11612 4811 11664 4820
rect 11612 4777 11621 4811
rect 11621 4777 11655 4811
rect 11655 4777 11664 4811
rect 11612 4768 11664 4777
rect 12440 4768 12492 4820
rect 15292 4811 15344 4820
rect 15292 4777 15301 4811
rect 15301 4777 15335 4811
rect 15335 4777 15344 4811
rect 15292 4768 15344 4777
rect 15476 4768 15528 4820
rect 19800 4768 19852 4820
rect 24032 4768 24084 4820
rect 9036 4632 9088 4684
rect 9128 4632 9180 4684
rect 9312 4675 9364 4684
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 8576 4496 8628 4548
rect 10232 4675 10284 4684
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 10324 4675 10376 4684
rect 10324 4641 10333 4675
rect 10333 4641 10367 4675
rect 10367 4641 10376 4675
rect 10324 4632 10376 4641
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 10876 4632 10928 4684
rect 11060 4632 11112 4684
rect 11244 4675 11296 4684
rect 11244 4641 11253 4675
rect 11253 4641 11287 4675
rect 11287 4641 11296 4675
rect 11244 4632 11296 4641
rect 14648 4700 14700 4752
rect 16672 4700 16724 4752
rect 17316 4700 17368 4752
rect 9680 4564 9732 4616
rect 12256 4632 12308 4684
rect 12440 4675 12492 4684
rect 12440 4641 12449 4675
rect 12449 4641 12483 4675
rect 12483 4641 12492 4675
rect 12440 4632 12492 4641
rect 12808 4632 12860 4684
rect 15200 4632 15252 4684
rect 15568 4632 15620 4684
rect 15844 4632 15896 4684
rect 17132 4675 17184 4684
rect 17132 4641 17141 4675
rect 17141 4641 17175 4675
rect 17175 4641 17184 4675
rect 17132 4632 17184 4641
rect 17960 4700 18012 4752
rect 18236 4700 18288 4752
rect 22468 4700 22520 4752
rect 24492 4700 24544 4752
rect 13084 4564 13136 4616
rect 14924 4564 14976 4616
rect 16396 4564 16448 4616
rect 18972 4632 19024 4684
rect 22652 4632 22704 4684
rect 22836 4675 22888 4684
rect 22836 4641 22870 4675
rect 22870 4641 22888 4675
rect 22836 4632 22888 4641
rect 9496 4496 9548 4548
rect 4896 4471 4948 4480
rect 4896 4437 4905 4471
rect 4905 4437 4939 4471
rect 4939 4437 4948 4471
rect 4896 4428 4948 4437
rect 4988 4428 5040 4480
rect 7380 4428 7432 4480
rect 9036 4428 9088 4480
rect 9772 4471 9824 4480
rect 9772 4437 9781 4471
rect 9781 4437 9815 4471
rect 9815 4437 9824 4471
rect 9772 4428 9824 4437
rect 11152 4428 11204 4480
rect 12256 4428 12308 4480
rect 15292 4496 15344 4548
rect 12716 4471 12768 4480
rect 12716 4437 12725 4471
rect 12725 4437 12759 4471
rect 12759 4437 12768 4471
rect 12716 4428 12768 4437
rect 14832 4428 14884 4480
rect 16120 4428 16172 4480
rect 19248 4428 19300 4480
rect 19800 4428 19852 4480
rect 3756 4326 3808 4378
rect 3820 4326 3872 4378
rect 3884 4326 3936 4378
rect 3948 4326 4000 4378
rect 4012 4326 4064 4378
rect 10472 4326 10524 4378
rect 10536 4326 10588 4378
rect 10600 4326 10652 4378
rect 10664 4326 10716 4378
rect 10728 4326 10780 4378
rect 17188 4326 17240 4378
rect 17252 4326 17304 4378
rect 17316 4326 17368 4378
rect 17380 4326 17432 4378
rect 17444 4326 17496 4378
rect 23904 4326 23956 4378
rect 23968 4326 24020 4378
rect 24032 4326 24084 4378
rect 24096 4326 24148 4378
rect 24160 4326 24212 4378
rect 5632 4224 5684 4276
rect 6368 4224 6420 4276
rect 12624 4267 12676 4276
rect 12624 4233 12633 4267
rect 12633 4233 12667 4267
rect 12667 4233 12676 4267
rect 12624 4224 12676 4233
rect 12992 4224 13044 4276
rect 14832 4224 14884 4276
rect 15292 4224 15344 4276
rect 6184 4088 6236 4140
rect 7104 4156 7156 4208
rect 7012 4088 7064 4140
rect 3700 3884 3752 3936
rect 3976 4063 4028 4072
rect 3976 4029 3985 4063
rect 3985 4029 4019 4063
rect 4019 4029 4028 4063
rect 3976 4020 4028 4029
rect 3884 3952 3936 4004
rect 5540 4020 5592 4072
rect 4896 3952 4948 4004
rect 7380 4020 7432 4072
rect 7472 4063 7524 4072
rect 7472 4029 7481 4063
rect 7481 4029 7515 4063
rect 7515 4029 7524 4063
rect 7472 4020 7524 4029
rect 7840 4020 7892 4072
rect 4988 3884 5040 3936
rect 6828 3927 6880 3936
rect 6828 3893 6837 3927
rect 6837 3893 6871 3927
rect 6871 3893 6880 3927
rect 6828 3884 6880 3893
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 8576 3884 8628 3893
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 9956 4156 10008 4208
rect 9772 4088 9824 4140
rect 9864 4063 9916 4072
rect 9864 4029 9873 4063
rect 9873 4029 9907 4063
rect 9907 4029 9916 4063
rect 9864 4020 9916 4029
rect 10324 4063 10376 4072
rect 10324 4029 10333 4063
rect 10333 4029 10367 4063
rect 10367 4029 10376 4063
rect 10324 4020 10376 4029
rect 14648 4156 14700 4208
rect 15016 4156 15068 4208
rect 15936 4224 15988 4276
rect 16304 4224 16356 4276
rect 11152 4063 11204 4072
rect 11152 4029 11161 4063
rect 11161 4029 11195 4063
rect 11195 4029 11204 4063
rect 11152 4020 11204 4029
rect 11244 4063 11296 4072
rect 11244 4029 11253 4063
rect 11253 4029 11287 4063
rect 11287 4029 11296 4063
rect 11244 4020 11296 4029
rect 12440 4063 12492 4072
rect 12440 4029 12449 4063
rect 12449 4029 12483 4063
rect 12483 4029 12492 4063
rect 12440 4020 12492 4029
rect 14648 4063 14700 4072
rect 14648 4029 14657 4063
rect 14657 4029 14691 4063
rect 14691 4029 14700 4063
rect 14648 4020 14700 4029
rect 15200 4088 15252 4140
rect 15016 4063 15068 4072
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15016 4020 15068 4029
rect 12072 3952 12124 4004
rect 14188 3952 14240 4004
rect 14280 3952 14332 4004
rect 17776 4156 17828 4208
rect 22100 4224 22152 4276
rect 22836 4267 22888 4276
rect 22836 4233 22845 4267
rect 22845 4233 22879 4267
rect 22879 4233 22888 4267
rect 22836 4224 22888 4233
rect 15936 4063 15988 4072
rect 15936 4029 15945 4063
rect 15945 4029 15979 4063
rect 15979 4029 15988 4063
rect 15936 4020 15988 4029
rect 16304 4063 16356 4072
rect 16304 4029 16313 4063
rect 16313 4029 16347 4063
rect 16347 4029 16356 4063
rect 16304 4020 16356 4029
rect 16580 4020 16632 4072
rect 16856 4020 16908 4072
rect 17776 4020 17828 4072
rect 19156 4088 19208 4140
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 11612 3927 11664 3936
rect 11612 3893 11621 3927
rect 11621 3893 11655 3927
rect 11655 3893 11664 3927
rect 11612 3884 11664 3893
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 15568 3995 15620 4004
rect 15568 3961 15577 3995
rect 15577 3961 15611 3995
rect 15611 3961 15620 3995
rect 15568 3952 15620 3961
rect 15844 3952 15896 4004
rect 16028 3884 16080 3936
rect 16212 3995 16264 4004
rect 16212 3961 16221 3995
rect 16221 3961 16255 3995
rect 16255 3961 16264 3995
rect 16212 3952 16264 3961
rect 23664 4020 23716 4072
rect 16304 3884 16356 3936
rect 18328 3927 18380 3936
rect 18328 3893 18337 3927
rect 18337 3893 18371 3927
rect 18371 3893 18380 3927
rect 18328 3884 18380 3893
rect 18512 3884 18564 3936
rect 18788 3884 18840 3936
rect 21456 3884 21508 3936
rect 7114 3782 7166 3834
rect 7178 3782 7230 3834
rect 7242 3782 7294 3834
rect 7306 3782 7358 3834
rect 7370 3782 7422 3834
rect 13830 3782 13882 3834
rect 13894 3782 13946 3834
rect 13958 3782 14010 3834
rect 14022 3782 14074 3834
rect 14086 3782 14138 3834
rect 20546 3782 20598 3834
rect 20610 3782 20662 3834
rect 20674 3782 20726 3834
rect 20738 3782 20790 3834
rect 20802 3782 20854 3834
rect 27262 3782 27314 3834
rect 27326 3782 27378 3834
rect 27390 3782 27442 3834
rect 27454 3782 27506 3834
rect 27518 3782 27570 3834
rect 4804 3680 4856 3732
rect 7840 3723 7892 3732
rect 7840 3689 7849 3723
rect 7849 3689 7883 3723
rect 7883 3689 7892 3723
rect 7840 3680 7892 3689
rect 10324 3680 10376 3732
rect 12440 3723 12492 3732
rect 12440 3689 12449 3723
rect 12449 3689 12483 3723
rect 12483 3689 12492 3723
rect 12440 3680 12492 3689
rect 13728 3680 13780 3732
rect 14372 3680 14424 3732
rect 3424 3612 3476 3664
rect 4160 3612 4212 3664
rect 5264 3612 5316 3664
rect 6828 3612 6880 3664
rect 3700 3587 3752 3596
rect 3700 3553 3709 3587
rect 3709 3553 3743 3587
rect 3743 3553 3752 3587
rect 3700 3544 3752 3553
rect 3332 3476 3384 3528
rect 3884 3544 3936 3596
rect 5540 3544 5592 3596
rect 6368 3544 6420 3596
rect 11612 3612 11664 3664
rect 8576 3587 8628 3596
rect 8576 3553 8610 3587
rect 8610 3553 8628 3587
rect 8576 3544 8628 3553
rect 9956 3544 10008 3596
rect 10968 3544 11020 3596
rect 15936 3680 15988 3732
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 12164 3544 12216 3596
rect 5172 3408 5224 3460
rect 5448 3408 5500 3460
rect 12716 3587 12768 3596
rect 12716 3553 12725 3587
rect 12725 3553 12759 3587
rect 12759 3553 12768 3587
rect 12716 3544 12768 3553
rect 15200 3612 15252 3664
rect 15108 3587 15160 3596
rect 15108 3553 15117 3587
rect 15117 3553 15151 3587
rect 15151 3553 15160 3587
rect 15108 3544 15160 3553
rect 3608 3340 3660 3392
rect 5540 3340 5592 3392
rect 6184 3340 6236 3392
rect 12900 3476 12952 3528
rect 14280 3476 14332 3528
rect 14556 3519 14608 3528
rect 14556 3485 14565 3519
rect 14565 3485 14599 3519
rect 14599 3485 14608 3519
rect 14556 3476 14608 3485
rect 16304 3587 16356 3596
rect 16304 3553 16313 3587
rect 16313 3553 16347 3587
rect 16347 3553 16356 3587
rect 16304 3544 16356 3553
rect 16396 3587 16448 3596
rect 16396 3553 16405 3587
rect 16405 3553 16439 3587
rect 16439 3553 16448 3587
rect 16396 3544 16448 3553
rect 16580 3544 16632 3596
rect 17776 3587 17828 3596
rect 17776 3553 17785 3587
rect 17785 3553 17819 3587
rect 17819 3553 17828 3587
rect 17776 3544 17828 3553
rect 18788 3680 18840 3732
rect 18328 3612 18380 3664
rect 18512 3587 18564 3596
rect 18512 3553 18521 3587
rect 18521 3553 18555 3587
rect 18555 3553 18564 3587
rect 18512 3544 18564 3553
rect 19064 3587 19116 3596
rect 19064 3553 19073 3587
rect 19073 3553 19107 3587
rect 19107 3553 19116 3587
rect 19064 3544 19116 3553
rect 21456 3544 21508 3596
rect 7472 3340 7524 3392
rect 8208 3340 8260 3392
rect 8300 3340 8352 3392
rect 18052 3408 18104 3460
rect 9864 3340 9916 3392
rect 12808 3340 12860 3392
rect 12900 3383 12952 3392
rect 12900 3349 12909 3383
rect 12909 3349 12943 3383
rect 12943 3349 12952 3383
rect 12900 3340 12952 3349
rect 13360 3340 13412 3392
rect 16212 3340 16264 3392
rect 16396 3340 16448 3392
rect 16580 3340 16632 3392
rect 17040 3340 17092 3392
rect 18328 3340 18380 3392
rect 18604 3340 18656 3392
rect 19984 3340 20036 3392
rect 3756 3238 3808 3290
rect 3820 3238 3872 3290
rect 3884 3238 3936 3290
rect 3948 3238 4000 3290
rect 4012 3238 4064 3290
rect 10472 3238 10524 3290
rect 10536 3238 10588 3290
rect 10600 3238 10652 3290
rect 10664 3238 10716 3290
rect 10728 3238 10780 3290
rect 17188 3238 17240 3290
rect 17252 3238 17304 3290
rect 17316 3238 17368 3290
rect 17380 3238 17432 3290
rect 17444 3238 17496 3290
rect 23904 3238 23956 3290
rect 23968 3238 24020 3290
rect 24032 3238 24084 3290
rect 24096 3238 24148 3290
rect 24160 3238 24212 3290
rect 5540 3136 5592 3188
rect 5724 3136 5776 3188
rect 4804 3068 4856 3120
rect 3332 3043 3384 3052
rect 3332 3009 3341 3043
rect 3341 3009 3375 3043
rect 3375 3009 3384 3043
rect 3332 3000 3384 3009
rect 3608 2975 3660 2984
rect 3608 2941 3642 2975
rect 3642 2941 3660 2975
rect 3608 2932 3660 2941
rect 5172 2932 5224 2984
rect 5540 2932 5592 2984
rect 5448 2907 5500 2916
rect 5448 2873 5457 2907
rect 5457 2873 5491 2907
rect 5491 2873 5500 2907
rect 5448 2864 5500 2873
rect 5724 2975 5776 2984
rect 5724 2941 5733 2975
rect 5733 2941 5767 2975
rect 5767 2941 5776 2975
rect 5724 2932 5776 2941
rect 5908 2975 5960 2984
rect 5908 2941 5917 2975
rect 5917 2941 5951 2975
rect 5951 2941 5960 2975
rect 5908 2932 5960 2941
rect 7840 3068 7892 3120
rect 10140 3179 10192 3188
rect 10140 3145 10149 3179
rect 10149 3145 10183 3179
rect 10183 3145 10192 3179
rect 10140 3136 10192 3145
rect 15108 3136 15160 3188
rect 15660 3136 15712 3188
rect 16028 3136 16080 3188
rect 18604 3136 18656 3188
rect 7472 2975 7524 2984
rect 7472 2941 7481 2975
rect 7481 2941 7515 2975
rect 7515 2941 7524 2975
rect 7472 2932 7524 2941
rect 8300 2932 8352 2984
rect 9956 2932 10008 2984
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 12440 3068 12492 3120
rect 14648 3068 14700 3120
rect 13728 3000 13780 3052
rect 15016 3000 15068 3052
rect 12716 2932 12768 2984
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 14556 2932 14608 2984
rect 16028 2975 16080 2984
rect 16028 2941 16037 2975
rect 16037 2941 16071 2975
rect 16071 2941 16080 2975
rect 16028 2932 16080 2941
rect 16304 3000 16356 3052
rect 16396 2975 16448 2984
rect 16396 2941 16405 2975
rect 16405 2941 16439 2975
rect 16439 2941 16448 2975
rect 16396 2932 16448 2941
rect 5080 2839 5132 2848
rect 5080 2805 5089 2839
rect 5089 2805 5123 2839
rect 5123 2805 5132 2839
rect 5080 2796 5132 2805
rect 5632 2796 5684 2848
rect 6276 2839 6328 2848
rect 6276 2805 6285 2839
rect 6285 2805 6319 2839
rect 6319 2805 6328 2839
rect 6276 2796 6328 2805
rect 7472 2796 7524 2848
rect 8024 2864 8076 2916
rect 10048 2864 10100 2916
rect 12256 2907 12308 2916
rect 12256 2873 12265 2907
rect 12265 2873 12299 2907
rect 12299 2873 12308 2907
rect 12256 2864 12308 2873
rect 16120 2864 16172 2916
rect 12440 2796 12492 2848
rect 12716 2839 12768 2848
rect 12716 2805 12725 2839
rect 12725 2805 12759 2839
rect 12759 2805 12768 2839
rect 12716 2796 12768 2805
rect 17040 2932 17092 2984
rect 17776 3000 17828 3052
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 19064 3136 19116 3188
rect 19892 3068 19944 3120
rect 16764 2796 16816 2848
rect 17224 2796 17276 2848
rect 7114 2694 7166 2746
rect 7178 2694 7230 2746
rect 7242 2694 7294 2746
rect 7306 2694 7358 2746
rect 7370 2694 7422 2746
rect 13830 2694 13882 2746
rect 13894 2694 13946 2746
rect 13958 2694 14010 2746
rect 14022 2694 14074 2746
rect 14086 2694 14138 2746
rect 20546 2694 20598 2746
rect 20610 2694 20662 2746
rect 20674 2694 20726 2746
rect 20738 2694 20790 2746
rect 20802 2694 20854 2746
rect 27262 2694 27314 2746
rect 27326 2694 27378 2746
rect 27390 2694 27442 2746
rect 27454 2694 27506 2746
rect 27518 2694 27570 2746
rect 5724 2592 5776 2644
rect 3608 2456 3660 2508
rect 4344 2456 4396 2508
rect 5080 2456 5132 2508
rect 6276 2456 6328 2508
rect 7472 2456 7524 2508
rect 8208 2456 8260 2508
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 9864 2524 9916 2576
rect 9772 2456 9824 2508
rect 10140 2592 10192 2644
rect 12256 2592 12308 2644
rect 12808 2592 12860 2644
rect 13084 2592 13136 2644
rect 14648 2635 14700 2644
rect 14648 2601 14657 2635
rect 14657 2601 14691 2635
rect 14691 2601 14700 2635
rect 14648 2592 14700 2601
rect 12716 2524 12768 2576
rect 13728 2524 13780 2576
rect 5448 2320 5500 2372
rect 5908 2320 5960 2372
rect 6920 2320 6972 2372
rect 8024 2320 8076 2372
rect 10324 2499 10376 2508
rect 10324 2465 10333 2499
rect 10333 2465 10367 2499
rect 10367 2465 10376 2499
rect 10324 2456 10376 2465
rect 10968 2456 11020 2508
rect 14924 2524 14976 2576
rect 16580 2567 16632 2576
rect 16580 2533 16589 2567
rect 16589 2533 16623 2567
rect 16623 2533 16632 2567
rect 16580 2524 16632 2533
rect 10232 2388 10284 2440
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 14464 2456 14516 2508
rect 15016 2499 15068 2508
rect 15016 2465 15025 2499
rect 15025 2465 15059 2499
rect 15059 2465 15068 2499
rect 15016 2456 15068 2465
rect 16764 2499 16816 2508
rect 16764 2465 16773 2499
rect 16773 2465 16807 2499
rect 16807 2465 16816 2499
rect 16764 2456 16816 2465
rect 17224 2499 17276 2508
rect 17224 2465 17233 2499
rect 17233 2465 17267 2499
rect 17267 2465 17276 2499
rect 17224 2456 17276 2465
rect 15384 2388 15436 2440
rect 16304 2431 16356 2440
rect 16304 2397 16313 2431
rect 16313 2397 16347 2431
rect 16347 2397 16356 2431
rect 16304 2388 16356 2397
rect 5816 2295 5868 2304
rect 5816 2261 5825 2295
rect 5825 2261 5859 2295
rect 5859 2261 5868 2295
rect 5816 2252 5868 2261
rect 6276 2295 6328 2304
rect 6276 2261 6285 2295
rect 6285 2261 6319 2295
rect 6319 2261 6328 2295
rect 6276 2252 6328 2261
rect 7656 2252 7708 2304
rect 8944 2252 8996 2304
rect 9680 2252 9732 2304
rect 9864 2252 9916 2304
rect 10876 2252 10928 2304
rect 14188 2320 14240 2372
rect 13912 2252 13964 2304
rect 16948 2295 17000 2304
rect 16948 2261 16957 2295
rect 16957 2261 16991 2295
rect 16991 2261 17000 2295
rect 16948 2252 17000 2261
rect 17040 2295 17092 2304
rect 17040 2261 17049 2295
rect 17049 2261 17083 2295
rect 17083 2261 17092 2295
rect 17040 2252 17092 2261
rect 3756 2150 3808 2202
rect 3820 2150 3872 2202
rect 3884 2150 3936 2202
rect 3948 2150 4000 2202
rect 4012 2150 4064 2202
rect 10472 2150 10524 2202
rect 10536 2150 10588 2202
rect 10600 2150 10652 2202
rect 10664 2150 10716 2202
rect 10728 2150 10780 2202
rect 17188 2150 17240 2202
rect 17252 2150 17304 2202
rect 17316 2150 17368 2202
rect 17380 2150 17432 2202
rect 17444 2150 17496 2202
rect 23904 2150 23956 2202
rect 23968 2150 24020 2202
rect 24032 2150 24084 2202
rect 24096 2150 24148 2202
rect 24160 2150 24212 2202
rect 4344 2091 4396 2100
rect 4344 2057 4353 2091
rect 4353 2057 4387 2091
rect 4387 2057 4396 2091
rect 4344 2048 4396 2057
rect 10324 2048 10376 2100
rect 6368 1955 6420 1964
rect 6368 1921 6377 1955
rect 6377 1921 6411 1955
rect 6411 1921 6420 1955
rect 6368 1912 6420 1921
rect 8668 1912 8720 1964
rect 9956 1955 10008 1964
rect 5816 1844 5868 1896
rect 6276 1844 6328 1896
rect 7656 1887 7708 1896
rect 7656 1853 7665 1887
rect 7665 1853 7699 1887
rect 7699 1853 7708 1887
rect 7656 1844 7708 1853
rect 8944 1887 8996 1896
rect 8944 1853 8953 1887
rect 8953 1853 8987 1887
rect 8987 1853 8996 1887
rect 8944 1844 8996 1853
rect 9680 1887 9732 1896
rect 9680 1853 9689 1887
rect 9689 1853 9723 1887
rect 9723 1853 9732 1887
rect 9680 1844 9732 1853
rect 9956 1921 9988 1955
rect 9988 1921 10008 1955
rect 15016 1980 15068 2032
rect 15292 2023 15344 2032
rect 15292 1989 15301 2023
rect 15301 1989 15335 2023
rect 15335 1989 15344 2023
rect 15292 1980 15344 1989
rect 9956 1912 10008 1921
rect 18512 1912 18564 1964
rect 20260 1955 20312 1964
rect 20260 1921 20269 1955
rect 20269 1921 20303 1955
rect 20303 1921 20312 1955
rect 20260 1912 20312 1921
rect 4896 1776 4948 1828
rect 6000 1776 6052 1828
rect 5632 1708 5684 1760
rect 6828 1708 6880 1760
rect 7564 1708 7616 1760
rect 9128 1751 9180 1760
rect 9128 1717 9137 1751
rect 9137 1717 9171 1751
rect 9171 1717 9180 1751
rect 9128 1708 9180 1717
rect 11520 1776 11572 1828
rect 12072 1776 12124 1828
rect 12440 1887 12492 1896
rect 12440 1853 12449 1887
rect 12449 1853 12483 1887
rect 12483 1853 12492 1887
rect 12440 1844 12492 1853
rect 12900 1844 12952 1896
rect 13912 1887 13964 1896
rect 13912 1853 13921 1887
rect 13921 1853 13955 1887
rect 13955 1853 13964 1887
rect 13912 1844 13964 1853
rect 14372 1887 14424 1896
rect 12992 1776 13044 1828
rect 14372 1853 14381 1887
rect 14381 1853 14415 1887
rect 14415 1853 14424 1887
rect 14372 1844 14424 1853
rect 14556 1844 14608 1896
rect 15016 1844 15068 1896
rect 15384 1844 15436 1896
rect 16764 1844 16816 1896
rect 17868 1844 17920 1896
rect 18420 1844 18472 1896
rect 18880 1844 18932 1896
rect 19800 1887 19852 1896
rect 19800 1853 19809 1887
rect 19809 1853 19843 1887
rect 19843 1853 19852 1887
rect 19800 1844 19852 1853
rect 19984 1887 20036 1896
rect 19984 1853 19993 1887
rect 19993 1853 20027 1887
rect 20027 1853 20036 1887
rect 19984 1844 20036 1853
rect 20352 1887 20404 1896
rect 20352 1853 20361 1887
rect 20361 1853 20395 1887
rect 20395 1853 20404 1887
rect 20352 1844 20404 1853
rect 21732 1844 21784 1896
rect 16948 1776 17000 1828
rect 17960 1776 18012 1828
rect 12900 1751 12952 1760
rect 12900 1717 12909 1751
rect 12909 1717 12943 1751
rect 12943 1717 12952 1751
rect 12900 1708 12952 1717
rect 15660 1751 15712 1760
rect 15660 1717 15669 1751
rect 15669 1717 15703 1751
rect 15703 1717 15712 1751
rect 15660 1708 15712 1717
rect 16028 1751 16080 1760
rect 16028 1717 16037 1751
rect 16037 1717 16071 1751
rect 16071 1717 16080 1751
rect 16028 1708 16080 1717
rect 16396 1708 16448 1760
rect 16488 1708 16540 1760
rect 18420 1708 18472 1760
rect 23572 1776 23624 1828
rect 21548 1708 21600 1760
rect 7114 1606 7166 1658
rect 7178 1606 7230 1658
rect 7242 1606 7294 1658
rect 7306 1606 7358 1658
rect 7370 1606 7422 1658
rect 13830 1606 13882 1658
rect 13894 1606 13946 1658
rect 13958 1606 14010 1658
rect 14022 1606 14074 1658
rect 14086 1606 14138 1658
rect 20546 1606 20598 1658
rect 20610 1606 20662 1658
rect 20674 1606 20726 1658
rect 20738 1606 20790 1658
rect 20802 1606 20854 1658
rect 27262 1606 27314 1658
rect 27326 1606 27378 1658
rect 27390 1606 27442 1658
rect 27454 1606 27506 1658
rect 27518 1606 27570 1658
rect 2596 1504 2648 1556
rect 6460 1504 6512 1556
rect 8300 1504 8352 1556
rect 10876 1504 10928 1556
rect 4344 1368 4396 1420
rect 4896 1411 4948 1420
rect 4896 1377 4905 1411
rect 4905 1377 4939 1411
rect 4939 1377 4948 1411
rect 4896 1368 4948 1377
rect 5724 1368 5776 1420
rect 7748 1436 7800 1488
rect 9128 1436 9180 1488
rect 6460 1411 6512 1420
rect 6460 1377 6469 1411
rect 6469 1377 6503 1411
rect 6503 1377 6512 1411
rect 6460 1368 6512 1377
rect 6828 1411 6880 1420
rect 6828 1377 6837 1411
rect 6837 1377 6871 1411
rect 6871 1377 6880 1411
rect 6828 1368 6880 1377
rect 7564 1411 7616 1420
rect 7564 1377 7598 1411
rect 7598 1377 7616 1411
rect 7564 1368 7616 1377
rect 8392 1368 8444 1420
rect 11520 1479 11572 1488
rect 11520 1445 11529 1479
rect 11529 1445 11563 1479
rect 11563 1445 11572 1479
rect 11520 1436 11572 1445
rect 11428 1411 11480 1420
rect 11428 1377 11432 1411
rect 11432 1377 11466 1411
rect 11466 1377 11480 1411
rect 11428 1368 11480 1377
rect 11612 1411 11664 1420
rect 11612 1377 11621 1411
rect 11621 1377 11655 1411
rect 11655 1377 11664 1411
rect 11612 1368 11664 1377
rect 12072 1547 12124 1556
rect 12072 1513 12081 1547
rect 12081 1513 12115 1547
rect 12115 1513 12124 1547
rect 12072 1504 12124 1513
rect 17960 1504 18012 1556
rect 18052 1504 18104 1556
rect 12900 1436 12952 1488
rect 15384 1436 15436 1488
rect 17040 1479 17092 1488
rect 17040 1445 17074 1479
rect 17074 1445 17092 1479
rect 17040 1436 17092 1445
rect 6736 1343 6788 1352
rect 6736 1309 6745 1343
rect 6745 1309 6779 1343
rect 6779 1309 6788 1343
rect 6736 1300 6788 1309
rect 6368 1232 6420 1284
rect 9956 1164 10008 1216
rect 11336 1164 11388 1216
rect 11888 1164 11940 1216
rect 14556 1411 14608 1420
rect 14556 1377 14565 1411
rect 14565 1377 14599 1411
rect 14599 1377 14608 1411
rect 14556 1368 14608 1377
rect 14096 1300 14148 1352
rect 14464 1300 14516 1352
rect 15200 1368 15252 1420
rect 15844 1368 15896 1420
rect 16304 1368 16356 1420
rect 16764 1343 16816 1352
rect 16764 1309 16773 1343
rect 16773 1309 16807 1343
rect 16807 1309 16816 1343
rect 16764 1300 16816 1309
rect 18420 1411 18472 1420
rect 18420 1377 18469 1411
rect 18469 1377 18472 1411
rect 18420 1368 18472 1377
rect 18880 1411 18932 1420
rect 18880 1377 18889 1411
rect 18889 1377 18923 1411
rect 18923 1377 18932 1411
rect 18880 1368 18932 1377
rect 18972 1411 19024 1420
rect 18972 1377 18981 1411
rect 18981 1377 19015 1411
rect 19015 1377 19024 1411
rect 18972 1368 19024 1377
rect 20076 1436 20128 1488
rect 19248 1411 19300 1420
rect 19248 1377 19257 1411
rect 19257 1377 19291 1411
rect 19291 1377 19300 1411
rect 19248 1368 19300 1377
rect 19800 1411 19852 1420
rect 19800 1377 19809 1411
rect 19809 1377 19843 1411
rect 19843 1377 19852 1411
rect 19800 1368 19852 1377
rect 19892 1411 19944 1420
rect 19892 1377 19901 1411
rect 19901 1377 19935 1411
rect 19935 1377 19944 1411
rect 19892 1368 19944 1377
rect 20352 1504 20404 1556
rect 21548 1504 21600 1556
rect 21824 1504 21876 1556
rect 25320 1436 25372 1488
rect 21456 1411 21508 1420
rect 21456 1377 21465 1411
rect 21465 1377 21499 1411
rect 21499 1377 21508 1411
rect 21456 1368 21508 1377
rect 21732 1368 21784 1420
rect 22008 1411 22060 1420
rect 22008 1377 22017 1411
rect 22017 1377 22051 1411
rect 22051 1377 22060 1411
rect 22008 1368 22060 1377
rect 22928 1368 22980 1420
rect 19800 1232 19852 1284
rect 14832 1164 14884 1216
rect 18328 1207 18380 1216
rect 18328 1173 18337 1207
rect 18337 1173 18371 1207
rect 18371 1173 18380 1207
rect 18328 1164 18380 1173
rect 3756 1062 3808 1114
rect 3820 1062 3872 1114
rect 3884 1062 3936 1114
rect 3948 1062 4000 1114
rect 4012 1062 4064 1114
rect 10472 1062 10524 1114
rect 10536 1062 10588 1114
rect 10600 1062 10652 1114
rect 10664 1062 10716 1114
rect 10728 1062 10780 1114
rect 17188 1062 17240 1114
rect 17252 1062 17304 1114
rect 17316 1062 17368 1114
rect 17380 1062 17432 1114
rect 17444 1062 17496 1114
rect 23904 1062 23956 1114
rect 23968 1062 24020 1114
rect 24032 1062 24084 1114
rect 24096 1062 24148 1114
rect 24160 1062 24212 1114
rect 11428 960 11480 1012
rect 12992 960 13044 1012
rect 14096 1003 14148 1012
rect 14096 969 14105 1003
rect 14105 969 14139 1003
rect 14139 969 14148 1003
rect 14096 960 14148 969
rect 6092 892 6144 944
rect 7840 892 7892 944
rect 9588 935 9640 944
rect 9588 901 9597 935
rect 9597 901 9631 935
rect 9631 901 9640 935
rect 9588 892 9640 901
rect 13084 935 13136 944
rect 13084 901 13093 935
rect 13093 901 13127 935
rect 13127 901 13136 935
rect 13084 892 13136 901
rect 6736 824 6788 876
rect 16580 892 16632 944
rect 19616 892 19668 944
rect 6184 799 6236 808
rect 6184 765 6193 799
rect 6193 765 6227 799
rect 6227 765 6236 799
rect 6184 756 6236 765
rect 6368 756 6420 808
rect 6552 756 6604 808
rect 7472 799 7524 808
rect 7472 765 7481 799
rect 7481 765 7515 799
rect 7515 765 7524 799
rect 7472 756 7524 765
rect 8300 688 8352 740
rect 9036 799 9088 808
rect 9036 765 9045 799
rect 9045 765 9079 799
rect 9079 765 9088 799
rect 9036 756 9088 765
rect 11428 756 11480 808
rect 11980 756 12032 808
rect 16764 824 16816 876
rect 19708 824 19760 876
rect 12808 799 12860 808
rect 12808 765 12817 799
rect 12817 765 12851 799
rect 12851 765 12860 799
rect 12808 756 12860 765
rect 12992 799 13044 808
rect 12992 765 12995 799
rect 12995 765 13044 799
rect 12992 756 13044 765
rect 15660 756 15712 808
rect 16120 799 16172 808
rect 16120 765 16129 799
rect 16129 765 16163 799
rect 16163 765 16172 799
rect 16120 756 16172 765
rect 16304 799 16356 808
rect 16304 765 16313 799
rect 16313 765 16347 799
rect 16347 765 16356 799
rect 16304 756 16356 765
rect 16396 799 16448 808
rect 16396 765 16405 799
rect 16405 765 16439 799
rect 16439 765 16448 799
rect 16396 756 16448 765
rect 16488 799 16540 808
rect 16488 765 16502 799
rect 16502 765 16536 799
rect 16536 765 16540 799
rect 16488 756 16540 765
rect 19800 799 19852 808
rect 19800 765 19809 799
rect 19809 765 19843 799
rect 19843 765 19852 799
rect 19800 756 19852 765
rect 20352 756 20404 808
rect 9864 688 9916 740
rect 11612 620 11664 672
rect 27068 688 27120 740
rect 7114 518 7166 570
rect 7178 518 7230 570
rect 7242 518 7294 570
rect 7306 518 7358 570
rect 7370 518 7422 570
rect 13830 518 13882 570
rect 13894 518 13946 570
rect 13958 518 14010 570
rect 14022 518 14074 570
rect 14086 518 14138 570
rect 20546 518 20598 570
rect 20610 518 20662 570
rect 20674 518 20726 570
rect 20738 518 20790 570
rect 20802 518 20854 570
rect 27262 518 27314 570
rect 27326 518 27378 570
rect 27390 518 27442 570
rect 27454 518 27506 570
rect 27518 518 27570 570
<< metal2 >>
rect 754 17762 810 18000
rect 1398 17762 1454 18000
rect 754 17734 888 17762
rect 754 17600 810 17734
rect 860 17338 888 17734
rect 1398 17734 1532 17762
rect 1398 17600 1454 17734
rect 1504 17338 1532 17734
rect 2042 17600 2098 18000
rect 2686 17600 2742 18000
rect 3330 17762 3386 18000
rect 3330 17734 3464 17762
rect 3330 17600 3386 17734
rect 848 17332 900 17338
rect 848 17274 900 17280
rect 1492 17332 1544 17338
rect 1492 17274 1544 17280
rect 2056 14890 2084 17600
rect 2700 17202 2728 17600
rect 3436 17202 3464 17734
rect 3974 17600 4030 18000
rect 4618 17762 4674 18000
rect 4618 17734 4752 17762
rect 4618 17600 4674 17734
rect 3988 17542 4016 17600
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3620 17338 3648 17478
rect 3756 17436 4064 17445
rect 3756 17434 3762 17436
rect 3818 17434 3842 17436
rect 3898 17434 3922 17436
rect 3978 17434 4002 17436
rect 4058 17434 4064 17436
rect 3818 17382 3820 17434
rect 4000 17382 4002 17434
rect 3756 17380 3762 17382
rect 3818 17380 3842 17382
rect 3898 17380 3922 17382
rect 3978 17380 4002 17382
rect 4058 17380 4064 17382
rect 3756 17371 4064 17380
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 4724 17202 4752 17734
rect 5262 17600 5318 18000
rect 5906 17600 5962 18000
rect 6550 17600 6606 18000
rect 7194 17762 7250 18000
rect 7194 17734 7512 17762
rect 7194 17600 7250 17734
rect 5276 17202 5304 17600
rect 5920 17338 5948 17600
rect 6564 17338 6592 17600
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 7114 16892 7422 16901
rect 7114 16890 7120 16892
rect 7176 16890 7200 16892
rect 7256 16890 7280 16892
rect 7336 16890 7360 16892
rect 7416 16890 7422 16892
rect 7176 16838 7178 16890
rect 7358 16838 7360 16890
rect 7114 16836 7120 16838
rect 7176 16836 7200 16838
rect 7256 16836 7280 16838
rect 7336 16836 7360 16838
rect 7416 16836 7422 16838
rect 7114 16827 7422 16836
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 3756 16348 4064 16357
rect 3756 16346 3762 16348
rect 3818 16346 3842 16348
rect 3898 16346 3922 16348
rect 3978 16346 4002 16348
rect 4058 16346 4064 16348
rect 3818 16294 3820 16346
rect 4000 16294 4002 16346
rect 3756 16292 3762 16294
rect 3818 16292 3842 16294
rect 3898 16292 3922 16294
rect 3978 16292 4002 16294
rect 4058 16292 4064 16294
rect 3756 16283 4064 16292
rect 5828 15570 5856 16526
rect 7484 16250 7512 17734
rect 7838 17600 7894 18000
rect 8482 17600 8538 18000
rect 9126 17600 9182 18000
rect 9770 17600 9826 18000
rect 10232 17604 10284 17610
rect 7852 17218 7880 17600
rect 8496 17338 8524 17600
rect 9140 17338 9168 17600
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 7852 17190 7972 17218
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7852 16454 7880 17070
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 6460 16176 6512 16182
rect 6460 16118 6512 16124
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 3756 15260 4064 15269
rect 3756 15258 3762 15260
rect 3818 15258 3842 15260
rect 3898 15258 3922 15260
rect 3978 15258 4002 15260
rect 4058 15258 4064 15260
rect 3818 15206 3820 15258
rect 4000 15206 4002 15258
rect 3756 15204 3762 15206
rect 3818 15204 3842 15206
rect 3898 15204 3922 15206
rect 3978 15204 4002 15206
rect 4058 15204 4064 15206
rect 3756 15195 4064 15204
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 2044 14884 2096 14890
rect 2044 14826 2096 14832
rect 2320 14816 2372 14822
rect 2320 14758 2372 14764
rect 2332 14482 2360 14758
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 1780 13802 1808 14214
rect 1768 13796 1820 13802
rect 1768 13738 1820 13744
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 13462 1992 13670
rect 1952 13456 2004 13462
rect 1952 13398 2004 13404
rect 2240 13326 2268 14214
rect 2424 13802 2452 14350
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2700 13870 2728 14214
rect 3252 14074 3280 14418
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3436 13870 3464 14350
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 3528 13870 3556 14282
rect 3620 14278 3648 14962
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 3804 14618 3832 14894
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 2412 13796 2464 13802
rect 2412 13738 2464 13744
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 2056 12714 2084 13126
rect 2424 12782 2452 13738
rect 2700 13394 2728 13806
rect 3620 13734 3648 14214
rect 3756 14172 4064 14181
rect 3756 14170 3762 14172
rect 3818 14170 3842 14172
rect 3898 14170 3922 14172
rect 3978 14170 4002 14172
rect 4058 14170 4064 14172
rect 3818 14118 3820 14170
rect 4000 14118 4002 14170
rect 3756 14116 3762 14118
rect 3818 14116 3842 14118
rect 3898 14116 3922 14118
rect 3978 14116 4002 14118
rect 4058 14116 4064 14118
rect 3756 14107 4064 14116
rect 4172 14074 4200 14894
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4172 13870 4200 14010
rect 4264 13870 4292 14418
rect 4632 14414 4660 15506
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5184 14890 5212 15302
rect 5828 14958 5856 15506
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5172 14884 5224 14890
rect 5172 14826 5224 14832
rect 6380 14618 6408 15506
rect 6472 15162 6500 16118
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4632 13938 4660 14214
rect 4816 14090 4844 14350
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4724 14074 4844 14090
rect 4712 14068 4844 14074
rect 4764 14062 4844 14068
rect 4712 14010 4764 14016
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 4160 13728 4212 13734
rect 4160 13670 4212 13676
rect 3620 13462 3648 13670
rect 4172 13530 4200 13670
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 3608 13456 3660 13462
rect 3608 13398 3660 13404
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 2976 12986 3004 13330
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2332 11626 2360 12038
rect 2424 11694 2452 12718
rect 3344 12714 3372 13126
rect 3436 12986 3464 13262
rect 3424 12980 3476 12986
rect 3620 12968 3648 13398
rect 4172 13190 4200 13466
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 3756 13084 4064 13093
rect 3756 13082 3762 13084
rect 3818 13082 3842 13084
rect 3898 13082 3922 13084
rect 3978 13082 4002 13084
rect 4058 13082 4064 13084
rect 3818 13030 3820 13082
rect 4000 13030 4002 13082
rect 3756 13028 3762 13030
rect 3818 13028 3842 13030
rect 3898 13028 3922 13030
rect 3978 13028 4002 13030
rect 4058 13028 4064 13030
rect 3756 13019 4064 13028
rect 3620 12940 3740 12968
rect 3424 12922 3476 12928
rect 3422 12880 3478 12889
rect 3422 12815 3478 12824
rect 3608 12844 3660 12850
rect 3436 12782 3464 12815
rect 3608 12786 3660 12792
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 3332 12708 3384 12714
rect 3332 12650 3384 12656
rect 2700 12306 2728 12650
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3252 12374 3280 12582
rect 3436 12442 3464 12582
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2424 10606 2452 11630
rect 3528 11354 3556 12242
rect 3620 12238 3648 12786
rect 3712 12782 3740 12940
rect 4172 12782 4200 13126
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 3712 12646 3740 12718
rect 4356 12714 4384 13806
rect 4816 13326 4844 14062
rect 4908 13870 4936 14214
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 5092 13258 5120 13670
rect 5184 13394 5212 13942
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5276 13462 5304 13670
rect 5552 13462 5580 13670
rect 5920 13530 5948 14282
rect 6182 13968 6238 13977
rect 6182 13903 6238 13912
rect 6196 13870 6224 13903
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4712 12912 4764 12918
rect 4710 12880 4712 12889
rect 4764 12880 4766 12889
rect 4710 12815 4766 12824
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 5000 12306 5028 13126
rect 5092 12986 5120 13194
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 5276 12442 5304 12650
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5644 12374 5672 13262
rect 6472 12918 6500 14554
rect 6564 14482 6592 14758
rect 6656 14550 6684 14758
rect 6644 14544 6696 14550
rect 6644 14486 6696 14492
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6644 14408 6696 14414
rect 6748 14396 6776 15914
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7114 15804 7422 15813
rect 7114 15802 7120 15804
rect 7176 15802 7200 15804
rect 7256 15802 7280 15804
rect 7336 15802 7360 15804
rect 7416 15802 7422 15804
rect 7176 15750 7178 15802
rect 7358 15750 7360 15802
rect 7114 15748 7120 15750
rect 7176 15748 7200 15750
rect 7256 15748 7280 15750
rect 7336 15748 7360 15750
rect 7416 15748 7422 15750
rect 7114 15739 7422 15748
rect 7484 15638 7512 15846
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6696 14368 6776 14396
rect 6644 14350 6696 14356
rect 6748 14074 6776 14368
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6840 13394 6868 14894
rect 6932 13870 6960 15370
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 7024 14958 7052 15302
rect 7484 15162 7512 15574
rect 7576 15450 7604 15982
rect 7852 15978 7880 16390
rect 7656 15972 7708 15978
rect 7656 15914 7708 15920
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 7668 15638 7696 15914
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 7576 15422 7696 15450
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 7024 14346 7052 14894
rect 7668 14890 7696 15422
rect 7656 14884 7708 14890
rect 7656 14826 7708 14832
rect 7114 14716 7422 14725
rect 7114 14714 7120 14716
rect 7176 14714 7200 14716
rect 7256 14714 7280 14716
rect 7336 14714 7360 14716
rect 7416 14714 7422 14716
rect 7176 14662 7178 14714
rect 7358 14662 7360 14714
rect 7114 14660 7120 14662
rect 7176 14660 7200 14662
rect 7256 14660 7280 14662
rect 7336 14660 7360 14662
rect 7416 14660 7422 14662
rect 7114 14651 7422 14660
rect 7012 14340 7064 14346
rect 7012 14282 7064 14288
rect 7564 14000 7616 14006
rect 7564 13942 7616 13948
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6932 13530 6960 13806
rect 7114 13628 7422 13637
rect 7114 13626 7120 13628
rect 7176 13626 7200 13628
rect 7256 13626 7280 13628
rect 7336 13626 7360 13628
rect 7416 13626 7422 13628
rect 7176 13574 7178 13626
rect 7358 13574 7360 13626
rect 7114 13572 7120 13574
rect 7176 13572 7200 13574
rect 7256 13572 7280 13574
rect 7336 13572 7360 13574
rect 7416 13572 7422 13574
rect 7114 13563 7422 13572
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7576 13462 7604 13942
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 6828 13388 6880 13394
rect 6748 13348 6828 13376
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6748 12782 6776 13348
rect 6828 13330 6880 13336
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7208 12986 7236 13330
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 5632 12368 5684 12374
rect 5632 12310 5684 12316
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 3620 12102 3648 12174
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11898 3648 12038
rect 3756 11996 4064 12005
rect 3756 11994 3762 11996
rect 3818 11994 3842 11996
rect 3898 11994 3922 11996
rect 3978 11994 4002 11996
rect 4058 11994 4064 11996
rect 3818 11942 3820 11994
rect 4000 11942 4002 11994
rect 3756 11940 3762 11942
rect 3818 11940 3842 11942
rect 3898 11940 3922 11942
rect 3978 11940 4002 11942
rect 4058 11940 4064 11942
rect 3756 11931 4064 11940
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 4816 11830 4844 12174
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 6104 11626 6132 12718
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6288 12374 6316 12582
rect 6840 12434 6868 12854
rect 7576 12782 7604 13126
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7114 12540 7422 12549
rect 7114 12538 7120 12540
rect 7176 12538 7200 12540
rect 7256 12538 7280 12540
rect 7336 12538 7360 12540
rect 7416 12538 7422 12540
rect 7176 12486 7178 12538
rect 7358 12486 7360 12538
rect 7114 12484 7120 12486
rect 7176 12484 7200 12486
rect 7256 12484 7280 12486
rect 7336 12484 7360 12486
rect 7416 12484 7422 12486
rect 7114 12475 7422 12484
rect 6656 12406 6868 12434
rect 7196 12436 7248 12442
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6656 12170 6684 12406
rect 7668 12434 7696 14826
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7760 14074 7788 14418
rect 7852 14278 7880 15914
rect 7944 15065 7972 17190
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8496 16250 8524 16594
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 9416 16046 9444 16934
rect 9784 16794 9812 17600
rect 10414 17604 10470 18000
rect 10414 17600 10416 17604
rect 10232 17546 10284 17552
rect 10468 17600 10470 17604
rect 11058 17600 11114 18000
rect 11702 17600 11758 18000
rect 12346 17600 12402 18000
rect 12990 17600 13046 18000
rect 13634 17600 13690 18000
rect 14278 17600 14334 18000
rect 14922 17600 14978 18000
rect 15566 17762 15622 18000
rect 16210 17762 16266 18000
rect 15566 17734 15884 17762
rect 15566 17600 15622 17734
rect 10416 17546 10468 17552
rect 10244 17338 10272 17546
rect 10472 17436 10780 17445
rect 10472 17434 10478 17436
rect 10534 17434 10558 17436
rect 10614 17434 10638 17436
rect 10694 17434 10718 17436
rect 10774 17434 10780 17436
rect 10534 17382 10536 17434
rect 10716 17382 10718 17434
rect 10472 17380 10478 17382
rect 10534 17380 10558 17382
rect 10614 17380 10638 17382
rect 10694 17380 10718 17382
rect 10774 17380 10780 17382
rect 10472 17371 10780 17380
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9692 16250 9720 16730
rect 9968 16658 9996 17070
rect 10796 16794 10824 17070
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10796 16658 10824 16730
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 10152 16046 10180 16390
rect 10472 16348 10780 16357
rect 10472 16346 10478 16348
rect 10534 16346 10558 16348
rect 10614 16346 10638 16348
rect 10694 16346 10718 16348
rect 10774 16346 10780 16348
rect 10534 16294 10536 16346
rect 10716 16294 10718 16346
rect 10472 16292 10478 16294
rect 10534 16292 10558 16294
rect 10614 16292 10638 16294
rect 10694 16292 10718 16294
rect 10774 16292 10780 16294
rect 10472 16283 10780 16292
rect 11072 16250 11100 17600
rect 11716 17338 11744 17600
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9680 16040 9732 16046
rect 10140 16040 10192 16046
rect 9732 16000 9904 16028
rect 9680 15982 9732 15988
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8680 15706 8708 15914
rect 8772 15706 8800 15982
rect 8864 15706 8892 15982
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 7930 15056 7986 15065
rect 7930 14991 7986 15000
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 8220 14006 8248 15506
rect 8680 15366 8708 15642
rect 9692 15638 9720 15846
rect 9680 15632 9732 15638
rect 9680 15574 9732 15580
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8300 14544 8352 14550
rect 8352 14492 8432 14498
rect 8300 14486 8432 14492
rect 8312 14470 8432 14486
rect 8496 14482 8524 14894
rect 8208 14000 8260 14006
rect 8206 13968 8208 13977
rect 8260 13968 8262 13977
rect 8206 13903 8262 13912
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7760 12918 7788 13670
rect 8312 13530 8340 13806
rect 8404 13802 8432 14470
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8392 13796 8444 13802
rect 8392 13738 8444 13744
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8404 13190 8432 13738
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 7748 12912 7800 12918
rect 7748 12854 7800 12860
rect 8392 12912 8444 12918
rect 8392 12854 8444 12860
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8128 12442 8156 12718
rect 8116 12436 8168 12442
rect 7668 12406 7788 12434
rect 7196 12378 7248 12384
rect 7208 12306 7236 12378
rect 7470 12336 7526 12345
rect 7196 12300 7248 12306
rect 7470 12271 7472 12280
rect 7196 12242 7248 12248
rect 7524 12271 7526 12280
rect 7472 12242 7524 12248
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2424 10130 2452 10542
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 1688 9178 1716 9386
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1872 9042 1900 9930
rect 2424 9518 2452 10066
rect 2884 9654 2912 10134
rect 3436 10130 3464 11154
rect 4816 11082 4844 11494
rect 5828 11150 5856 11562
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 3756 10908 4064 10917
rect 3756 10906 3762 10908
rect 3818 10906 3842 10908
rect 3898 10906 3922 10908
rect 3978 10906 4002 10908
rect 4058 10906 4064 10908
rect 3818 10854 3820 10906
rect 4000 10854 4002 10906
rect 3756 10852 3762 10854
rect 3818 10852 3842 10854
rect 3898 10852 3922 10854
rect 3978 10852 4002 10854
rect 4058 10852 4064 10854
rect 3756 10843 4064 10852
rect 5828 10606 5856 11086
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5632 10532 5684 10538
rect 5632 10474 5684 10480
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 3068 9518 3096 9862
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 1860 9036 1912 9042
rect 2056 9024 2084 9114
rect 2884 9042 2912 9318
rect 1912 8996 2084 9024
rect 1860 8978 1912 8984
rect 2056 8906 2084 8996
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 3160 8974 3188 9386
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 2044 8900 2096 8906
rect 2044 8842 2096 8848
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 1504 6866 1532 8366
rect 2240 8362 2268 8774
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2332 6866 2360 8910
rect 3160 8634 3188 8910
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 3436 8378 3464 10066
rect 3620 9654 3648 10202
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 3756 9820 4064 9829
rect 3756 9818 3762 9820
rect 3818 9818 3842 9820
rect 3898 9818 3922 9820
rect 3978 9818 4002 9820
rect 4058 9818 4064 9820
rect 3818 9766 3820 9818
rect 4000 9766 4002 9818
rect 3756 9764 3762 9766
rect 3818 9764 3842 9766
rect 3898 9764 3922 9766
rect 3978 9764 4002 9766
rect 4058 9764 4064 9766
rect 3756 9755 4064 9764
rect 3608 9648 3660 9654
rect 3608 9590 3660 9596
rect 4172 9518 4200 9862
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 3620 8514 3648 9454
rect 4448 8838 4476 9454
rect 5000 9450 5028 9930
rect 5460 9518 5488 10066
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 9654 5580 9862
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5644 9586 5672 10474
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10198 5764 10406
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 9042 4660 9318
rect 5000 9178 5028 9386
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5172 9104 5224 9110
rect 5170 9072 5172 9081
rect 5224 9072 5226 9081
rect 4620 9036 4672 9042
rect 5170 9007 5226 9016
rect 4620 8978 4672 8984
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 3756 8732 4064 8741
rect 3756 8730 3762 8732
rect 3818 8730 3842 8732
rect 3898 8730 3922 8732
rect 3978 8730 4002 8732
rect 4058 8730 4064 8732
rect 3818 8678 3820 8730
rect 4000 8678 4002 8730
rect 3756 8676 3762 8678
rect 3818 8676 3842 8678
rect 3898 8676 3922 8678
rect 3978 8676 4002 8678
rect 4058 8676 4064 8678
rect 3756 8667 4064 8676
rect 4344 8560 4396 8566
rect 3620 8498 3832 8514
rect 4344 8502 4396 8508
rect 3620 8492 3844 8498
rect 3620 8486 3792 8492
rect 3792 8434 3844 8440
rect 4068 8424 4120 8430
rect 3514 8392 3570 8401
rect 2700 7954 2728 8366
rect 3436 8350 3514 8378
rect 4068 8366 4120 8372
rect 3514 8327 3570 8336
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2424 7546 2452 7890
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2056 6458 2084 6802
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2332 6322 2360 6802
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2608 6254 2636 6666
rect 2700 6322 2728 7890
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2884 6254 2912 6394
rect 3068 6254 3096 6598
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3344 6186 3372 7414
rect 3436 7274 3464 8230
rect 3528 7546 3556 8327
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3620 7410 3648 8230
rect 4080 8090 4108 8366
rect 4356 8294 4384 8502
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4448 8294 4476 8434
rect 4528 8356 4580 8362
rect 4632 8344 4660 8978
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4816 8838 4844 8910
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4580 8316 4660 8344
rect 4528 8298 4580 8304
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3756 7644 4064 7653
rect 3756 7642 3762 7644
rect 3818 7642 3842 7644
rect 3898 7642 3922 7644
rect 3978 7642 4002 7644
rect 4058 7642 4064 7644
rect 3818 7590 3820 7642
rect 4000 7590 4002 7642
rect 3756 7588 3762 7590
rect 3818 7588 3842 7590
rect 3898 7588 3922 7590
rect 3978 7588 4002 7590
rect 4058 7588 4064 7590
rect 3756 7579 4064 7588
rect 4356 7426 4384 8230
rect 3608 7404 3660 7410
rect 4356 7398 4568 7426
rect 3608 7346 3660 7352
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3528 6866 3556 7278
rect 3620 7002 3648 7346
rect 4540 7342 4568 7398
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4172 7018 4200 7278
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4172 7002 4292 7018
rect 3608 6996 3660 7002
rect 4172 6996 4304 7002
rect 4172 6990 4252 6996
rect 3608 6938 3660 6944
rect 4252 6938 4304 6944
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 3528 5710 3556 6802
rect 3620 6458 3648 6938
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 3756 6556 4064 6565
rect 3756 6554 3762 6556
rect 3818 6554 3842 6556
rect 3898 6554 3922 6556
rect 3978 6554 4002 6556
rect 4058 6554 4064 6556
rect 3818 6502 3820 6554
rect 4000 6502 4002 6554
rect 3756 6500 3762 6502
rect 3818 6500 3842 6502
rect 3898 6500 3922 6502
rect 3978 6500 4002 6502
rect 4058 6500 4064 6502
rect 3756 6491 4064 6500
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 4264 5778 4292 6598
rect 4356 6186 4384 7142
rect 4448 6662 4476 7278
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4540 6118 4568 7278
rect 4816 7206 4844 8774
rect 5736 8430 5764 9386
rect 5828 9042 5856 10542
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 6104 10266 6132 10474
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6656 10130 6684 12106
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6932 11286 6960 12038
rect 7114 11452 7422 11461
rect 7114 11450 7120 11452
rect 7176 11450 7200 11452
rect 7256 11450 7280 11452
rect 7336 11450 7360 11452
rect 7416 11450 7422 11452
rect 7176 11398 7178 11450
rect 7358 11398 7360 11450
rect 7114 11396 7120 11398
rect 7176 11396 7200 11398
rect 7256 11396 7280 11398
rect 7336 11396 7360 11398
rect 7416 11396 7422 11398
rect 7114 11387 7422 11396
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4816 6458 4844 6802
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 5184 5574 5212 6122
rect 5276 5794 5304 7142
rect 5368 7002 5396 7278
rect 5460 7002 5488 7346
rect 5736 7342 5764 8366
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5920 7546 5948 7754
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5368 6730 5396 6938
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5276 5766 5488 5794
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 3756 5468 4064 5477
rect 3756 5466 3762 5468
rect 3818 5466 3842 5468
rect 3898 5466 3922 5468
rect 3978 5466 4002 5468
rect 4058 5466 4064 5468
rect 3818 5414 3820 5466
rect 4000 5414 4002 5466
rect 3756 5412 3762 5414
rect 3818 5412 3842 5414
rect 3898 5412 3922 5414
rect 3978 5412 4002 5414
rect 4058 5412 4064 5414
rect 3756 5403 4064 5412
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4080 4690 4108 5306
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5368 4690 5396 5170
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5460 4622 5488 5766
rect 5552 5166 5580 6190
rect 5736 5846 5764 6598
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3436 3670 3464 4422
rect 3756 4380 4064 4389
rect 3756 4378 3762 4380
rect 3818 4378 3842 4380
rect 3898 4378 3922 4380
rect 3978 4378 4002 4380
rect 4058 4378 4064 4380
rect 3818 4326 3820 4378
rect 4000 4326 4002 4378
rect 3756 4324 3762 4326
rect 3818 4324 3842 4326
rect 3898 4324 3922 4326
rect 3978 4324 4002 4326
rect 4058 4324 4064 4326
rect 3756 4315 4064 4324
rect 3976 4072 4028 4078
rect 4028 4032 4200 4060
rect 3976 4014 4028 4020
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 3712 3602 3740 3878
rect 3896 3602 3924 3946
rect 4172 3670 4200 4032
rect 4816 3738 4844 4558
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4908 4010 4936 4422
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 5000 3942 5028 4422
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3344 3058 3372 3470
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3344 2774 3372 2994
rect 3620 2990 3648 3334
rect 3756 3292 4064 3301
rect 3756 3290 3762 3292
rect 3818 3290 3842 3292
rect 3898 3290 3922 3292
rect 3978 3290 4002 3292
rect 4058 3290 4064 3292
rect 3818 3238 3820 3290
rect 4000 3238 4002 3290
rect 3756 3236 3762 3238
rect 3818 3236 3842 3238
rect 3898 3236 3922 3238
rect 3978 3236 4002 3238
rect 4058 3236 4064 3238
rect 3756 3227 4064 3236
rect 4816 3126 4844 3674
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 5184 2990 5212 3402
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 3344 2746 3648 2774
rect 3620 2514 3648 2746
rect 5092 2514 5120 2790
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 4344 2508 4396 2514
rect 4344 2450 4396 2456
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 3756 2204 4064 2213
rect 3756 2202 3762 2204
rect 3818 2202 3842 2204
rect 3898 2202 3922 2204
rect 3978 2202 4002 2204
rect 4058 2202 4064 2204
rect 3818 2150 3820 2202
rect 4000 2150 4002 2202
rect 3756 2148 3762 2150
rect 3818 2148 3842 2150
rect 3898 2148 3922 2150
rect 3978 2148 4002 2150
rect 4058 2148 4064 2150
rect 3756 2139 4064 2148
rect 4356 2106 4384 2450
rect 5276 2446 5304 3606
rect 5460 3466 5488 4558
rect 5552 4078 5580 5102
rect 5644 4690 5672 5306
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5920 5030 5948 5102
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5920 4758 5948 4966
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5552 3602 5580 4014
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5552 3194 5580 3334
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5540 2984 5592 2990
rect 5644 2972 5672 4218
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5736 2990 5764 3130
rect 5592 2944 5672 2972
rect 5724 2984 5776 2990
rect 5540 2926 5592 2932
rect 5724 2926 5776 2932
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5460 2378 5488 2858
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 4344 2100 4396 2106
rect 4344 2042 4396 2048
rect 846 1864 902 1873
rect 846 1799 902 1808
rect 4896 1828 4948 1834
rect 860 400 888 1799
rect 4896 1770 4948 1776
rect 2596 1556 2648 1562
rect 2596 1498 2648 1504
rect 2608 400 2636 1498
rect 4908 1426 4936 1770
rect 5644 1766 5672 2790
rect 5736 2650 5764 2926
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5632 1760 5684 1766
rect 5632 1702 5684 1708
rect 5736 1426 5764 2586
rect 5920 2378 5948 2926
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5828 1902 5856 2246
rect 6012 2009 6040 9454
rect 6104 9450 6132 10066
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6380 9722 6408 9930
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6092 9444 6144 9450
rect 6092 9386 6144 9392
rect 6288 7886 6316 9454
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6196 6662 6224 7278
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6288 6458 6316 6666
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6288 5778 6316 6394
rect 6366 6216 6422 6225
rect 6366 6151 6368 6160
rect 6420 6151 6422 6160
rect 6368 6122 6420 6128
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6380 4282 6408 4558
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6196 3398 6224 4082
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 5998 2000 6054 2009
rect 5998 1935 6054 1944
rect 5816 1896 5868 1902
rect 5816 1838 5868 1844
rect 6012 1834 6040 1935
rect 6000 1828 6052 1834
rect 6000 1770 6052 1776
rect 4344 1420 4396 1426
rect 4344 1362 4396 1368
rect 4896 1420 4948 1426
rect 4896 1362 4948 1368
rect 5724 1420 5776 1426
rect 5724 1362 5776 1368
rect 3756 1116 4064 1125
rect 3756 1114 3762 1116
rect 3818 1114 3842 1116
rect 3898 1114 3922 1116
rect 3978 1114 4002 1116
rect 4058 1114 4064 1116
rect 3818 1062 3820 1114
rect 4000 1062 4002 1114
rect 3756 1060 3762 1062
rect 3818 1060 3842 1062
rect 3898 1060 3922 1062
rect 3978 1060 4002 1062
rect 4058 1060 4064 1062
rect 3756 1051 4064 1060
rect 4356 400 4384 1362
rect 6092 944 6144 950
rect 6092 886 6144 892
rect 6104 400 6132 886
rect 6196 814 6224 3334
rect 6276 2848 6328 2854
rect 6276 2790 6328 2796
rect 6288 2514 6316 2790
rect 6276 2508 6328 2514
rect 6276 2450 6328 2456
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6288 1902 6316 2246
rect 6380 1970 6408 3538
rect 6472 2553 6500 9862
rect 6656 9518 6684 10066
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6748 9450 6776 10950
rect 6840 9586 6868 11018
rect 7300 10810 7328 11086
rect 7484 11014 7512 12242
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7576 11898 7604 12106
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7114 10364 7422 10373
rect 7114 10362 7120 10364
rect 7176 10362 7200 10364
rect 7256 10362 7280 10364
rect 7336 10362 7360 10364
rect 7416 10362 7422 10364
rect 7176 10310 7178 10362
rect 7358 10310 7360 10362
rect 7114 10308 7120 10310
rect 7176 10308 7200 10310
rect 7256 10308 7280 10310
rect 7336 10308 7360 10310
rect 7416 10308 7422 10310
rect 7114 10299 7422 10308
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7208 9926 7236 10066
rect 7668 9994 7696 12106
rect 7760 11665 7788 12406
rect 8116 12378 8168 12384
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7746 11656 7802 11665
rect 7746 11591 7802 11600
rect 7852 11257 7880 11834
rect 8036 11354 8064 12174
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 8128 11286 8156 12378
rect 8116 11280 8168 11286
rect 7838 11248 7894 11257
rect 8116 11222 8168 11228
rect 7838 11183 7894 11192
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7196 9920 7248 9926
rect 7760 9874 7788 10542
rect 7196 9862 7248 9868
rect 7668 9846 7788 9874
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6748 7954 6776 9386
rect 7114 9276 7422 9285
rect 7114 9274 7120 9276
rect 7176 9274 7200 9276
rect 7256 9274 7280 9276
rect 7336 9274 7360 9276
rect 7416 9274 7422 9276
rect 7176 9222 7178 9274
rect 7358 9222 7360 9274
rect 7114 9220 7120 9222
rect 7176 9220 7200 9222
rect 7256 9220 7280 9222
rect 7336 9220 7360 9222
rect 7416 9220 7422 9222
rect 7114 9211 7422 9220
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7024 8634 7052 8978
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 7024 8072 7052 8298
rect 7114 8188 7422 8197
rect 7114 8186 7120 8188
rect 7176 8186 7200 8188
rect 7256 8186 7280 8188
rect 7336 8186 7360 8188
rect 7416 8186 7422 8188
rect 7176 8134 7178 8186
rect 7358 8134 7360 8186
rect 7114 8132 7120 8134
rect 7176 8132 7200 8134
rect 7256 8132 7280 8134
rect 7336 8132 7360 8134
rect 7416 8132 7422 8134
rect 7114 8123 7422 8132
rect 7024 8044 7328 8072
rect 7300 7954 7328 8044
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7380 7948 7432 7954
rect 7484 7936 7512 8774
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7576 8090 7604 8366
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7668 7970 7696 9846
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 8090 7788 8230
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7432 7908 7512 7936
rect 7576 7942 7696 7970
rect 7380 7890 7432 7896
rect 6748 7546 6776 7890
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6840 7342 6868 7686
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6564 6798 6592 7278
rect 7114 7100 7422 7109
rect 7114 7098 7120 7100
rect 7176 7098 7200 7100
rect 7256 7098 7280 7100
rect 7336 7098 7360 7100
rect 7416 7098 7422 7100
rect 7176 7046 7178 7098
rect 7358 7046 7360 7098
rect 7114 7044 7120 7046
rect 7176 7044 7200 7046
rect 7256 7044 7280 7046
rect 7336 7044 7360 7046
rect 7416 7044 7422 7046
rect 7114 7035 7422 7044
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 6564 6254 6592 6734
rect 7484 6254 7512 6734
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7114 6012 7422 6021
rect 7114 6010 7120 6012
rect 7176 6010 7200 6012
rect 7256 6010 7280 6012
rect 7336 6010 7360 6012
rect 7416 6010 7422 6012
rect 7176 5958 7178 6010
rect 7358 5958 7360 6010
rect 7114 5956 7120 5958
rect 7176 5956 7200 5958
rect 7256 5956 7280 5958
rect 7336 5956 7360 5958
rect 7416 5956 7422 5958
rect 7114 5947 7422 5956
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7208 5166 7236 5306
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 6932 5030 6960 5102
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 4826 6960 4966
rect 7114 4924 7422 4933
rect 7114 4922 7120 4924
rect 7176 4922 7200 4924
rect 7256 4922 7280 4924
rect 7336 4922 7360 4924
rect 7416 4922 7422 4924
rect 7176 4870 7178 4922
rect 7358 4870 7360 4922
rect 7114 4868 7120 4870
rect 7176 4868 7200 4870
rect 7256 4868 7280 4870
rect 7336 4868 7360 4870
rect 7416 4868 7422 4870
rect 7114 4859 7422 4868
rect 6920 4820 6972 4826
rect 6972 4780 7052 4808
rect 6920 4762 6972 4768
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6840 3670 6868 3878
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6458 2544 6514 2553
rect 6514 2502 6592 2530
rect 6458 2479 6514 2488
rect 6368 1964 6420 1970
rect 6368 1906 6420 1912
rect 6276 1896 6328 1902
rect 6276 1838 6328 1844
rect 6380 1290 6408 1906
rect 6460 1556 6512 1562
rect 6460 1498 6512 1504
rect 6472 1426 6500 1498
rect 6460 1420 6512 1426
rect 6460 1362 6512 1368
rect 6368 1284 6420 1290
rect 6368 1226 6420 1232
rect 6184 808 6236 814
rect 6184 750 6236 756
rect 6368 808 6420 814
rect 6472 796 6500 1362
rect 6564 814 6592 2502
rect 6932 2378 6960 4626
rect 7024 4146 7052 4780
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7116 4214 7144 4626
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7392 4078 7420 4422
rect 7484 4078 7512 5306
rect 7576 4690 7604 7942
rect 7852 7936 7880 11183
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7944 10606 7972 10950
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7944 10062 7972 10542
rect 8128 10146 8156 11222
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8220 10266 8248 11154
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8312 10606 8340 11086
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8128 10118 8248 10146
rect 8312 10130 8340 10406
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 8220 9926 8248 10118
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8128 9178 8156 9454
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8220 8974 8248 9862
rect 8312 9178 8340 10066
rect 8404 9466 8432 12854
rect 8496 11694 8524 13670
rect 8680 12850 8708 15302
rect 9692 14958 9720 15574
rect 9876 15502 9904 16000
rect 10140 15982 10192 15988
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 9048 14482 9076 14758
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9416 13734 9444 14350
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8680 12434 8708 12582
rect 8588 12406 8708 12434
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8588 11234 8616 12406
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8680 11694 8708 12310
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8496 11206 8616 11234
rect 8772 11218 8800 12106
rect 8864 11694 8892 13126
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8668 11212 8720 11218
rect 8496 10538 8524 11206
rect 8668 11154 8720 11160
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8588 10690 8616 11086
rect 8680 10810 8708 11154
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8588 10662 8708 10690
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 8496 10112 8524 10474
rect 8588 10266 8616 10542
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8576 10124 8628 10130
rect 8496 10084 8576 10112
rect 8576 10066 8628 10072
rect 8680 9926 8708 10662
rect 8772 10538 8800 11154
rect 8864 10742 8892 11630
rect 8956 11558 8984 12242
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9232 11898 9260 12174
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8760 10532 8812 10538
rect 8760 10474 8812 10480
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8404 9438 8524 9466
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8404 9110 8432 9318
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8220 8362 8248 8910
rect 8496 8514 8524 9438
rect 8680 8634 8708 9862
rect 8772 9518 8800 10202
rect 8864 10130 8892 10678
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8956 10266 8984 10542
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8864 9178 8892 10066
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8772 8906 8800 9114
rect 8956 9042 8984 9998
rect 9048 9994 9076 11290
rect 9324 11286 9352 11630
rect 9416 11354 9444 12242
rect 9600 12238 9628 14486
rect 9692 13954 9720 14894
rect 9876 14890 9904 15438
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9864 14884 9916 14890
rect 9864 14826 9916 14832
rect 9864 14544 9916 14550
rect 9862 14512 9864 14521
rect 9916 14512 9918 14521
rect 9862 14447 9918 14456
rect 9968 14362 9996 15098
rect 10060 14958 10088 15370
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 10060 14822 10088 14894
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10152 14480 10180 15846
rect 10336 15337 10364 16186
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 10322 15328 10378 15337
rect 10322 15263 10378 15272
rect 10472 15260 10780 15269
rect 10472 15258 10478 15260
rect 10534 15258 10558 15260
rect 10614 15258 10638 15260
rect 10694 15258 10718 15260
rect 10774 15258 10780 15260
rect 10534 15206 10536 15258
rect 10716 15206 10718 15258
rect 10472 15204 10478 15206
rect 10534 15204 10558 15206
rect 10614 15204 10638 15206
rect 10694 15204 10718 15206
rect 10774 15204 10780 15206
rect 10472 15195 10780 15204
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10140 14474 10192 14480
rect 10140 14416 10192 14422
rect 10244 14362 10272 15030
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 9876 14334 9996 14362
rect 10152 14334 10272 14362
rect 10336 14464 10364 14758
rect 10612 14618 10640 14758
rect 10888 14618 10916 15982
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 11072 15858 11100 15982
rect 11164 15978 11192 16594
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11152 15972 11204 15978
rect 11152 15914 11204 15920
rect 10980 15570 11008 15846
rect 11072 15830 11192 15858
rect 10968 15564 11020 15570
rect 11020 15524 11100 15552
rect 10968 15506 11020 15512
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10980 15094 11008 15370
rect 11072 15162 11100 15524
rect 11164 15366 11192 15830
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11164 14958 11192 15030
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 11164 14822 11192 14894
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 11164 14482 11192 14758
rect 10416 14476 10468 14482
rect 10336 14436 10416 14464
rect 9876 14074 9904 14334
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9692 13926 9812 13954
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9692 13394 9720 13806
rect 9784 13802 9812 13926
rect 9876 13870 9904 14010
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9784 13326 9812 13738
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9692 12850 9720 13194
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9680 12436 9732 12442
rect 9784 12434 9812 12582
rect 9732 12406 9812 12434
rect 9680 12378 9732 12384
rect 9876 12306 9904 12786
rect 9968 12782 9996 14214
rect 10152 13802 10180 14334
rect 10336 13818 10364 14436
rect 10416 14418 10468 14424
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 10472 14172 10780 14181
rect 10472 14170 10478 14172
rect 10534 14170 10558 14172
rect 10614 14170 10638 14172
rect 10694 14170 10718 14172
rect 10774 14170 10780 14172
rect 10534 14118 10536 14170
rect 10716 14118 10718 14170
rect 10472 14116 10478 14118
rect 10534 14116 10558 14118
rect 10614 14116 10638 14118
rect 10694 14116 10718 14118
rect 10774 14116 10780 14118
rect 10472 14107 10780 14116
rect 10888 13954 10916 14418
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10796 13926 10916 13954
rect 10140 13796 10192 13802
rect 10336 13790 10732 13818
rect 10140 13738 10192 13744
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9600 11393 9628 11562
rect 9586 11384 9642 11393
rect 9404 11348 9456 11354
rect 9586 11319 9642 11328
rect 9404 11290 9456 11296
rect 9692 11286 9720 12038
rect 9968 11762 9996 12718
rect 10060 12646 10088 13126
rect 10152 12782 10180 13738
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10520 13462 10548 13670
rect 10508 13456 10560 13462
rect 10508 13398 10560 13404
rect 10704 13326 10732 13790
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10796 13190 10824 13926
rect 10876 13796 10928 13802
rect 10876 13738 10928 13744
rect 10888 13530 10916 13738
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10472 13084 10780 13093
rect 10472 13082 10478 13084
rect 10534 13082 10558 13084
rect 10614 13082 10638 13084
rect 10694 13082 10718 13084
rect 10774 13082 10780 13084
rect 10534 13030 10536 13082
rect 10716 13030 10718 13082
rect 10472 13028 10478 13030
rect 10534 13028 10558 13030
rect 10614 13028 10638 13030
rect 10694 13028 10718 13030
rect 10774 13028 10780 13030
rect 10472 13019 10780 13028
rect 10888 12986 10916 13330
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10980 12918 11008 14214
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 13394 11100 13670
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10060 12345 10088 12582
rect 11256 12434 11284 16050
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11348 15162 11376 15506
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11440 15026 11468 15302
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11348 14482 11376 14758
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 11532 14226 11560 15982
rect 11796 15972 11848 15978
rect 11796 15914 11848 15920
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11624 14618 11652 15642
rect 11716 15026 11744 15846
rect 11808 15570 11836 15914
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11796 15428 11848 15434
rect 11796 15370 11848 15376
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11440 14198 11560 14226
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11348 13530 11376 13670
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11348 13394 11376 13466
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11164 12406 11284 12434
rect 10046 12336 10102 12345
rect 10046 12271 10102 12280
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9140 10130 9168 10950
rect 9600 10606 9628 10950
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 9048 9058 9076 9930
rect 9232 9518 9260 10406
rect 9600 10198 9628 10542
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 8944 9036 8996 9042
rect 9048 9030 9168 9058
rect 8944 8978 8996 8984
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8404 8486 8524 8514
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8404 7970 8432 8486
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8496 8090 8524 8366
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8588 8090 8616 8298
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8404 7942 8616 7970
rect 7760 7908 7880 7936
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 7668 4758 7696 5238
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7114 3836 7422 3845
rect 7114 3834 7120 3836
rect 7176 3834 7200 3836
rect 7256 3834 7280 3836
rect 7336 3834 7360 3836
rect 7416 3834 7422 3836
rect 7176 3782 7178 3834
rect 7358 3782 7360 3834
rect 7114 3780 7120 3782
rect 7176 3780 7200 3782
rect 7256 3780 7280 3782
rect 7336 3780 7360 3782
rect 7416 3780 7422 3782
rect 7114 3771 7422 3780
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7484 2990 7512 3334
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7114 2748 7422 2757
rect 7114 2746 7120 2748
rect 7176 2746 7200 2748
rect 7256 2746 7280 2748
rect 7336 2746 7360 2748
rect 7416 2746 7422 2748
rect 7176 2694 7178 2746
rect 7358 2694 7360 2746
rect 7114 2692 7120 2694
rect 7176 2692 7200 2694
rect 7256 2692 7280 2694
rect 7336 2692 7360 2694
rect 7416 2692 7422 2694
rect 7114 2683 7422 2692
rect 7484 2514 7512 2790
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7668 1902 7696 2246
rect 7656 1896 7708 1902
rect 7656 1838 7708 1844
rect 6828 1760 6880 1766
rect 6828 1702 6880 1708
rect 7564 1760 7616 1766
rect 7564 1702 7616 1708
rect 6840 1426 6868 1702
rect 7114 1660 7422 1669
rect 7114 1658 7120 1660
rect 7176 1658 7200 1660
rect 7256 1658 7280 1660
rect 7336 1658 7360 1660
rect 7416 1658 7422 1660
rect 7176 1606 7178 1658
rect 7358 1606 7360 1658
rect 7114 1604 7120 1606
rect 7176 1604 7200 1606
rect 7256 1604 7280 1606
rect 7336 1604 7360 1606
rect 7416 1604 7422 1606
rect 7114 1595 7422 1604
rect 7470 1456 7526 1465
rect 6828 1420 6880 1426
rect 7576 1426 7604 1702
rect 7760 1494 7788 7908
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 7852 5250 7880 7754
rect 7944 7546 7972 7822
rect 8588 7818 8616 7942
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 7852 5222 7972 5250
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7852 3738 7880 4014
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7852 3126 7880 3674
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7748 1488 7800 1494
rect 7944 1465 7972 5222
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 8036 4758 8064 5102
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 8128 4672 8156 6870
rect 8312 6866 8340 7142
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8220 5030 8248 5646
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8312 4826 8340 5102
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8312 4690 8340 4762
rect 8208 4684 8260 4690
rect 8128 4644 8208 4672
rect 8208 4626 8260 4632
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8024 2916 8076 2922
rect 8024 2858 8076 2864
rect 8036 2378 8064 2858
rect 8220 2514 8248 3334
rect 8312 2990 8340 3334
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8024 2372 8076 2378
rect 8024 2314 8076 2320
rect 8312 1562 8340 2926
rect 8300 1556 8352 1562
rect 8300 1498 8352 1504
rect 7748 1430 7800 1436
rect 7930 1456 7986 1465
rect 7470 1391 7526 1400
rect 7564 1420 7616 1426
rect 6828 1362 6880 1368
rect 6736 1352 6788 1358
rect 6736 1294 6788 1300
rect 6748 882 6776 1294
rect 6736 876 6788 882
rect 6736 818 6788 824
rect 7484 814 7512 1391
rect 7930 1391 7986 1400
rect 7564 1362 7616 1368
rect 7840 944 7892 950
rect 7840 886 7892 892
rect 6420 768 6500 796
rect 6552 808 6604 814
rect 6368 750 6420 756
rect 6552 750 6604 756
rect 7472 808 7524 814
rect 7472 750 7524 756
rect 7114 572 7422 581
rect 7114 570 7120 572
rect 7176 570 7200 572
rect 7256 570 7280 572
rect 7336 570 7360 572
rect 7416 570 7422 572
rect 7176 518 7178 570
rect 7358 518 7360 570
rect 7114 516 7120 518
rect 7176 516 7200 518
rect 7256 516 7280 518
rect 7336 516 7360 518
rect 7416 516 7422 518
rect 7114 507 7422 516
rect 7852 400 7880 886
rect 8312 746 8340 1498
rect 8404 1426 8432 7346
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8496 5914 8524 6734
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8588 5778 8616 7754
rect 8680 6882 8708 8570
rect 8772 8430 8800 8842
rect 8956 8566 8984 8978
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 9048 8634 9076 8842
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8944 8560 8996 8566
rect 8944 8502 8996 8508
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8772 7002 8800 7822
rect 8864 7342 8892 8230
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8680 6854 8800 6882
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8680 5914 8708 6122
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8772 5166 8800 6854
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8864 5166 8892 5714
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8760 4820 8812 4826
rect 8864 4808 8892 5102
rect 8812 4780 8892 4808
rect 8760 4762 8812 4768
rect 8864 4729 8892 4780
rect 8850 4720 8906 4729
rect 8576 4684 8628 4690
rect 8850 4655 8906 4664
rect 8576 4626 8628 4632
rect 8588 4554 8616 4626
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8588 3602 8616 3878
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8668 2440 8720 2446
rect 8956 2417 8984 7686
rect 9048 7342 9076 7890
rect 9140 7834 9168 9030
rect 9232 8498 9260 9454
rect 9324 9178 9352 9590
rect 9600 9518 9628 10134
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9324 8430 9352 8978
rect 9416 8906 9444 9386
rect 9508 9364 9536 9454
rect 9680 9376 9732 9382
rect 9508 9336 9680 9364
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9324 7954 9352 8366
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9140 7806 9352 7834
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 6458 9076 7278
rect 9218 6896 9274 6905
rect 9218 6831 9274 6840
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9048 5574 9076 6054
rect 9140 5778 9168 6054
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9140 5234 9168 5714
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 9048 4690 9076 5034
rect 9140 4690 9168 5170
rect 9232 4826 9260 6831
rect 9324 5166 9352 7806
rect 9416 6905 9444 8366
rect 9508 7954 9536 9336
rect 9680 9318 9732 9324
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9784 8566 9812 9046
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9600 8430 9628 8502
rect 9784 8430 9812 8502
rect 9588 8424 9640 8430
rect 9772 8424 9824 8430
rect 9640 8384 9720 8412
rect 9588 8366 9640 8372
rect 9692 7954 9720 8384
rect 9772 8366 9824 8372
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9680 7948 9732 7954
rect 9784 7936 9812 8366
rect 9864 7948 9916 7954
rect 9784 7908 9864 7936
rect 9680 7890 9732 7896
rect 9864 7890 9916 7896
rect 9508 6934 9536 7890
rect 9862 7848 9918 7857
rect 9862 7783 9864 7792
rect 9916 7783 9918 7792
rect 9864 7754 9916 7760
rect 9496 6928 9548 6934
rect 9402 6896 9458 6905
rect 9496 6870 9548 6876
rect 9402 6831 9458 6840
rect 9968 5370 9996 11494
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 10060 8022 10088 8842
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9416 5030 9444 5102
rect 9680 5092 9732 5098
rect 9680 5034 9732 5040
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9310 4720 9366 4729
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 9128 4684 9180 4690
rect 9416 4706 9444 4966
rect 9588 4820 9640 4826
rect 9366 4678 9444 4706
rect 9508 4780 9588 4808
rect 9310 4655 9312 4664
rect 9128 4626 9180 4632
rect 9364 4655 9366 4664
rect 9312 4626 9364 4632
rect 9508 4554 9536 4780
rect 9588 4762 9640 4768
rect 9692 4622 9720 5034
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9048 4078 9076 4422
rect 9784 4146 9812 4422
rect 9968 4214 9996 5306
rect 10152 4826 10180 12174
rect 10472 11996 10780 12005
rect 10472 11994 10478 11996
rect 10534 11994 10558 11996
rect 10614 11994 10638 11996
rect 10694 11994 10718 11996
rect 10774 11994 10780 11996
rect 10534 11942 10536 11994
rect 10716 11942 10718 11994
rect 10472 11940 10478 11942
rect 10534 11940 10558 11942
rect 10614 11940 10638 11942
rect 10694 11940 10718 11942
rect 10774 11940 10780 11942
rect 10472 11931 10780 11940
rect 10472 10908 10780 10917
rect 10472 10906 10478 10908
rect 10534 10906 10558 10908
rect 10614 10906 10638 10908
rect 10694 10906 10718 10908
rect 10774 10906 10780 10908
rect 10534 10854 10536 10906
rect 10716 10854 10718 10906
rect 10472 10852 10478 10854
rect 10534 10852 10558 10854
rect 10614 10852 10638 10854
rect 10694 10852 10718 10854
rect 10774 10852 10780 10854
rect 10472 10843 10780 10852
rect 10472 9820 10780 9829
rect 10472 9818 10478 9820
rect 10534 9818 10558 9820
rect 10614 9818 10638 9820
rect 10694 9818 10718 9820
rect 10774 9818 10780 9820
rect 10534 9766 10536 9818
rect 10716 9766 10718 9818
rect 10472 9764 10478 9766
rect 10534 9764 10558 9766
rect 10614 9764 10638 9766
rect 10694 9764 10718 9766
rect 10774 9764 10780 9766
rect 10472 9755 10780 9764
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10472 8732 10780 8741
rect 10472 8730 10478 8732
rect 10534 8730 10558 8732
rect 10614 8730 10638 8732
rect 10694 8730 10718 8732
rect 10774 8730 10780 8732
rect 10534 8678 10536 8730
rect 10716 8678 10718 8730
rect 10472 8676 10478 8678
rect 10534 8676 10558 8678
rect 10614 8676 10638 8678
rect 10694 8676 10718 8678
rect 10774 8676 10780 8678
rect 10472 8667 10780 8676
rect 10980 8634 11008 9046
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10428 8294 10456 8434
rect 10980 8362 11008 8570
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10336 7954 10364 8230
rect 10428 7954 10456 8230
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10472 7644 10780 7653
rect 10472 7642 10478 7644
rect 10534 7642 10558 7644
rect 10614 7642 10638 7644
rect 10694 7642 10718 7644
rect 10774 7642 10780 7644
rect 10534 7590 10536 7642
rect 10716 7590 10718 7642
rect 10472 7588 10478 7590
rect 10534 7588 10558 7590
rect 10614 7588 10638 7590
rect 10694 7588 10718 7590
rect 10774 7588 10780 7590
rect 10472 7579 10780 7588
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10244 6390 10272 6666
rect 10472 6556 10780 6565
rect 10472 6554 10478 6556
rect 10534 6554 10558 6556
rect 10614 6554 10638 6556
rect 10694 6554 10718 6556
rect 10774 6554 10780 6556
rect 10534 6502 10536 6554
rect 10716 6502 10718 6554
rect 10472 6500 10478 6502
rect 10534 6500 10558 6502
rect 10614 6500 10638 6502
rect 10694 6500 10718 6502
rect 10774 6500 10780 6502
rect 10472 6491 10780 6500
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10598 6352 10654 6361
rect 10244 6254 10272 6326
rect 10888 6322 10916 7210
rect 10598 6287 10654 6296
rect 10876 6316 10928 6322
rect 10612 6254 10640 6287
rect 10876 6258 10928 6264
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10244 4690 10272 6054
rect 10428 5914 10456 6190
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10428 5624 10456 5850
rect 10888 5710 10916 6122
rect 10980 5778 11008 7278
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11072 6322 11100 6734
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 10876 5704 10928 5710
rect 10336 5596 10456 5624
rect 10782 5672 10838 5681
rect 10876 5646 10928 5652
rect 10782 5607 10784 5616
rect 10336 5030 10364 5596
rect 10836 5607 10838 5616
rect 10784 5578 10836 5584
rect 10472 5468 10780 5477
rect 10472 5466 10478 5468
rect 10534 5466 10558 5468
rect 10614 5466 10638 5468
rect 10694 5466 10718 5468
rect 10774 5466 10780 5468
rect 10534 5414 10536 5466
rect 10716 5414 10718 5466
rect 10472 5412 10478 5414
rect 10534 5412 10558 5414
rect 10614 5412 10638 5414
rect 10694 5412 10718 5414
rect 10774 5412 10780 5414
rect 10472 5403 10780 5412
rect 10980 5370 11008 5714
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10336 4690 10364 4966
rect 10612 4690 10640 5170
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10796 4570 10824 4762
rect 10888 4690 10916 5238
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10796 4542 10916 4570
rect 10472 4380 10780 4389
rect 10472 4378 10478 4380
rect 10534 4378 10558 4380
rect 10614 4378 10638 4380
rect 10694 4378 10718 4380
rect 10774 4378 10780 4380
rect 10534 4326 10536 4378
rect 10716 4326 10718 4378
rect 10472 4324 10478 4326
rect 10534 4324 10558 4326
rect 10614 4324 10638 4326
rect 10694 4324 10718 4326
rect 10774 4324 10780 4326
rect 10472 4315 10780 4324
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 9876 3398 9904 4014
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9876 2582 9904 3334
rect 9968 2990 9996 3538
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 9968 2530 9996 2926
rect 10060 2922 10088 3878
rect 10336 3738 10364 4014
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10152 3194 10180 3470
rect 10472 3292 10780 3301
rect 10472 3290 10478 3292
rect 10534 3290 10558 3292
rect 10614 3290 10638 3292
rect 10694 3290 10718 3292
rect 10774 3290 10780 3292
rect 10534 3238 10536 3290
rect 10716 3238 10718 3290
rect 10472 3236 10478 3238
rect 10534 3236 10558 3238
rect 10614 3236 10638 3238
rect 10694 3236 10718 3238
rect 10774 3236 10780 3238
rect 10472 3227 10780 3236
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10048 2916 10100 2922
rect 10048 2858 10100 2864
rect 10152 2650 10180 3130
rect 10888 2774 10916 4542
rect 10980 3602 11008 5306
rect 11072 4690 11100 5714
rect 11164 5302 11192 12406
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11348 8498 11376 8978
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11256 7886 11284 8366
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11256 6118 11284 7482
rect 11348 7274 11376 7686
rect 11440 7290 11468 14198
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11532 12306 11560 13738
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11532 11762 11560 12242
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11532 11218 11560 11698
rect 11624 11694 11652 12038
rect 11716 11694 11744 13126
rect 11808 12986 11836 15370
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11900 12434 11928 17070
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 11992 13870 12020 14894
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 12084 14074 12112 14350
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 12084 12850 12112 13670
rect 12176 13394 12204 17206
rect 12360 16810 12388 17600
rect 12268 16782 12388 16810
rect 13004 16794 13032 17600
rect 13648 17338 13676 17600
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13830 16892 14138 16901
rect 13830 16890 13836 16892
rect 13892 16890 13916 16892
rect 13972 16890 13996 16892
rect 14052 16890 14076 16892
rect 14132 16890 14138 16892
rect 13892 16838 13894 16890
rect 14074 16838 14076 16890
rect 13830 16836 13836 16838
rect 13892 16836 13916 16838
rect 13972 16836 13996 16838
rect 14052 16836 14076 16838
rect 14132 16836 14138 16838
rect 13830 16827 14138 16836
rect 14292 16794 14320 17600
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 12992 16788 13044 16794
rect 12268 16250 12296 16782
rect 12992 16730 13044 16736
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 14002 16688 14058 16697
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12360 15570 12388 16594
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12452 15706 12480 15982
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12636 15638 12664 15982
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12360 14890 12388 15506
rect 12728 15065 12756 16662
rect 12992 16652 13044 16658
rect 14002 16623 14004 16632
rect 12992 16594 13044 16600
rect 14056 16623 14058 16632
rect 14280 16652 14332 16658
rect 14004 16594 14056 16600
rect 14280 16594 14332 16600
rect 12714 15056 12770 15065
rect 12714 14991 12770 15000
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11808 12406 11928 12434
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11532 9586 11560 11154
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11336 7268 11388 7274
rect 11440 7262 11652 7290
rect 11336 7210 11388 7216
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11440 6866 11468 7142
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11348 6390 11376 6598
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11440 6254 11468 6598
rect 11624 6458 11652 7262
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11426 5264 11482 5273
rect 11426 5199 11482 5208
rect 11440 5166 11468 5199
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11532 4826 11560 5102
rect 11624 4826 11652 5714
rect 11808 5370 11836 12406
rect 11992 11608 12020 12718
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12084 11898 12112 12242
rect 12176 12102 12204 12378
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12176 11694 12204 12038
rect 12728 11830 12756 12038
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12072 11620 12124 11626
rect 11992 11580 12072 11608
rect 12072 11562 12124 11568
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11900 9178 11928 9386
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11900 8498 11928 8910
rect 12084 8537 12112 11562
rect 12176 10266 12204 11630
rect 12452 11626 12480 11766
rect 12440 11620 12492 11626
rect 12440 11562 12492 11568
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12438 11384 12494 11393
rect 12438 11319 12494 11328
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12348 10192 12400 10198
rect 12348 10134 12400 10140
rect 12256 10124 12308 10130
rect 12176 10084 12256 10112
rect 12176 9178 12204 10084
rect 12256 10066 12308 10072
rect 12360 9450 12388 10134
rect 12452 9625 12480 11319
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12438 9616 12494 9625
rect 12438 9551 12494 9560
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12070 8528 12126 8537
rect 11888 8492 11940 8498
rect 12070 8463 12126 8472
rect 11888 8434 11940 8440
rect 12176 8430 12204 9114
rect 12360 9042 12388 9386
rect 12440 9376 12492 9382
rect 12438 9344 12440 9353
rect 12492 9344 12494 9353
rect 12438 9279 12494 9288
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 12084 6866 12112 8298
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12176 7206 12204 7822
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 11886 6352 11942 6361
rect 11886 6287 11942 6296
rect 11900 6254 11928 6287
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 4078 11192 4422
rect 11256 4078 11284 4626
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11624 3670 11652 3878
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10888 2746 11008 2774
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9968 2502 10272 2530
rect 10980 2514 11008 2746
rect 8668 2382 8720 2388
rect 8942 2408 8998 2417
rect 8680 1970 8708 2382
rect 9784 2394 9812 2450
rect 8998 2366 9076 2394
rect 9784 2366 9904 2394
rect 8942 2343 8998 2352
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8668 1964 8720 1970
rect 8668 1906 8720 1912
rect 8956 1902 8984 2246
rect 8944 1896 8996 1902
rect 8944 1838 8996 1844
rect 8392 1420 8444 1426
rect 8392 1362 8444 1368
rect 9048 814 9076 2366
rect 9876 2310 9904 2366
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 9692 1902 9720 2246
rect 9680 1896 9732 1902
rect 9680 1838 9732 1844
rect 9128 1760 9180 1766
rect 9128 1702 9180 1708
rect 9140 1494 9168 1702
rect 9128 1488 9180 1494
rect 9128 1430 9180 1436
rect 9588 944 9640 950
rect 9588 886 9640 892
rect 9036 808 9088 814
rect 9036 750 9088 756
rect 8300 740 8352 746
rect 8300 682 8352 688
rect 9600 400 9628 886
rect 9876 746 9904 2246
rect 9968 1970 9996 2502
rect 10244 2446 10272 2502
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10336 2106 10364 2450
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10472 2204 10780 2213
rect 10472 2202 10478 2204
rect 10534 2202 10558 2204
rect 10614 2202 10638 2204
rect 10694 2202 10718 2204
rect 10774 2202 10780 2204
rect 10534 2150 10536 2202
rect 10716 2150 10718 2202
rect 10472 2148 10478 2150
rect 10534 2148 10558 2150
rect 10614 2148 10638 2150
rect 10694 2148 10718 2150
rect 10774 2148 10780 2150
rect 10472 2139 10780 2148
rect 10324 2100 10376 2106
rect 10324 2042 10376 2048
rect 9956 1964 10008 1970
rect 9956 1906 10008 1912
rect 9968 1222 9996 1906
rect 10888 1562 10916 2246
rect 11520 1828 11572 1834
rect 11520 1770 11572 1776
rect 10876 1556 10928 1562
rect 10876 1498 10928 1504
rect 11532 1494 11560 1770
rect 11520 1488 11572 1494
rect 11520 1430 11572 1436
rect 11428 1420 11480 1426
rect 11428 1362 11480 1368
rect 11612 1420 11664 1426
rect 11612 1362 11664 1368
rect 9956 1216 10008 1222
rect 9956 1158 10008 1164
rect 11336 1216 11388 1222
rect 11336 1158 11388 1164
rect 10472 1116 10780 1125
rect 10472 1114 10478 1116
rect 10534 1114 10558 1116
rect 10614 1114 10638 1116
rect 10694 1114 10718 1116
rect 10774 1114 10780 1116
rect 10534 1062 10536 1114
rect 10716 1062 10718 1114
rect 10472 1060 10478 1062
rect 10534 1060 10558 1062
rect 10614 1060 10638 1062
rect 10694 1060 10718 1062
rect 10774 1060 10780 1062
rect 10472 1051 10780 1060
rect 9864 740 9916 746
rect 9864 682 9916 688
rect 11348 400 11376 1158
rect 11440 1018 11468 1362
rect 11428 1012 11480 1018
rect 11428 954 11480 960
rect 11440 814 11468 954
rect 11428 808 11480 814
rect 11428 750 11480 756
rect 11624 678 11652 1362
rect 11900 1222 11928 2382
rect 11888 1216 11940 1222
rect 11888 1158 11940 1164
rect 11992 814 12020 6054
rect 12176 5166 12204 7142
rect 12268 6866 12296 8774
rect 12360 8430 12388 8842
rect 12544 8566 12572 10678
rect 12636 10606 12664 11494
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12728 10810 12756 11222
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12820 10146 12848 11562
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12912 10266 12940 10542
rect 13004 10266 13032 16594
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 16046 13400 16390
rect 14292 16046 14320 16594
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13096 15638 13124 15846
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 13372 15162 13400 15982
rect 13830 15804 14138 15813
rect 13830 15802 13836 15804
rect 13892 15802 13916 15804
rect 13972 15802 13996 15804
rect 14052 15802 14076 15804
rect 14132 15802 14138 15804
rect 13892 15750 13894 15802
rect 14074 15750 14076 15802
rect 13830 15748 13836 15750
rect 13892 15748 13916 15750
rect 13972 15748 13996 15750
rect 14052 15748 14076 15750
rect 14132 15748 14138 15750
rect 13830 15739 14138 15748
rect 14292 15434 14320 15982
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13372 14482 13400 15098
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13556 14482 13584 14758
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13096 10690 13124 14418
rect 13740 14346 13768 14758
rect 13830 14716 14138 14725
rect 13830 14714 13836 14716
rect 13892 14714 13916 14716
rect 13972 14714 13996 14716
rect 14052 14714 14076 14716
rect 14132 14714 14138 14716
rect 13892 14662 13894 14714
rect 14074 14662 14076 14714
rect 13830 14660 13836 14662
rect 13892 14660 13916 14662
rect 13972 14660 13996 14662
rect 14052 14660 14076 14662
rect 14132 14660 14138 14662
rect 13830 14651 14138 14660
rect 14002 14512 14058 14521
rect 14002 14447 14058 14456
rect 14016 14414 14044 14447
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 14096 13864 14148 13870
rect 14200 13818 14228 14894
rect 14292 14498 14320 15370
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14384 14618 14412 14826
rect 14476 14618 14504 15302
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14292 14470 14504 14498
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14384 14074 14412 14350
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14148 13812 14228 13818
rect 14096 13806 14228 13812
rect 14108 13790 14228 13806
rect 13830 13628 14138 13637
rect 13830 13626 13836 13628
rect 13892 13626 13916 13628
rect 13972 13626 13996 13628
rect 14052 13626 14076 13628
rect 14132 13626 14138 13628
rect 13892 13574 13894 13626
rect 14074 13574 14076 13626
rect 13830 13572 13836 13574
rect 13892 13572 13916 13574
rect 13972 13572 13996 13574
rect 14052 13572 14076 13574
rect 14132 13572 14138 13574
rect 13830 13563 14138 13572
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13372 13161 13400 13262
rect 13636 13184 13688 13190
rect 13358 13152 13414 13161
rect 13636 13126 13688 13132
rect 13358 13087 13414 13096
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13188 12714 13216 12922
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13188 11762 13216 12650
rect 13648 12306 13676 13126
rect 14200 12782 14228 13790
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 13830 12540 14138 12549
rect 13830 12538 13836 12540
rect 13892 12538 13916 12540
rect 13972 12538 13996 12540
rect 14052 12538 14076 12540
rect 14132 12538 14138 12540
rect 13892 12486 13894 12538
rect 14074 12486 14076 12538
rect 13830 12484 13836 12486
rect 13892 12484 13916 12486
rect 13972 12484 13996 12486
rect 14052 12484 14076 12486
rect 14132 12484 14138 12486
rect 13830 12475 14138 12484
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13832 11898 13860 12378
rect 14200 12374 14228 12718
rect 14292 12442 14320 13262
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14384 12782 14412 13126
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14280 12436 14332 12442
rect 14476 12434 14504 14470
rect 14280 12378 14332 12384
rect 14384 12406 14504 12434
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13740 11354 13768 11698
rect 13924 11694 13952 12242
rect 14384 12186 14412 12406
rect 14200 12158 14412 12186
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14094 11792 14150 11801
rect 14200 11778 14228 12158
rect 14200 11750 14320 11778
rect 14094 11727 14096 11736
rect 14148 11727 14150 11736
rect 14096 11698 14148 11704
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13830 11452 14138 11461
rect 13830 11450 13836 11452
rect 13892 11450 13916 11452
rect 13972 11450 13996 11452
rect 14052 11450 14076 11452
rect 14132 11450 14138 11452
rect 13892 11398 13894 11450
rect 14074 11398 14076 11450
rect 13830 11396 13836 11398
rect 13892 11396 13916 11398
rect 13972 11396 13996 11398
rect 14052 11396 14076 11398
rect 14132 11396 14138 11398
rect 13830 11387 14138 11396
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 13096 10662 13216 10690
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12624 10124 12676 10130
rect 12820 10118 12940 10146
rect 12624 10066 12676 10072
rect 12636 8634 12664 10066
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12532 8560 12584 8566
rect 12452 8508 12532 8514
rect 12452 8502 12584 8508
rect 12452 8486 12572 8502
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12452 8362 12480 8486
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12348 7948 12400 7954
rect 12452 7936 12480 8298
rect 12544 8090 12572 8366
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12400 7908 12480 7936
rect 12716 7948 12768 7954
rect 12348 7890 12400 7896
rect 12768 7908 12848 7936
rect 12716 7890 12768 7896
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12360 7342 12388 7754
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12820 7206 12848 7908
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12820 6905 12848 7142
rect 12806 6896 12862 6905
rect 12256 6860 12308 6866
rect 12806 6831 12862 6840
rect 12256 6802 12308 6808
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 12084 2990 12112 3946
rect 12176 3602 12204 5102
rect 12452 4826 12480 5578
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12440 4684 12492 4690
rect 12544 4672 12572 5646
rect 12820 5166 12848 6831
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12492 4644 12572 4672
rect 12440 4626 12492 4632
rect 12268 4486 12296 4626
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12084 1834 12112 2926
rect 12268 2922 12296 4422
rect 12636 4282 12664 4966
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12452 3738 12480 4014
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12452 3126 12480 3674
rect 12728 3602 12756 4422
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12820 3482 12848 4626
rect 12912 3534 12940 10118
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13004 8430 13032 9454
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 13004 6254 13032 8366
rect 13096 8362 13124 10542
rect 13188 9518 13216 10662
rect 13830 10364 14138 10373
rect 13830 10362 13836 10364
rect 13892 10362 13916 10364
rect 13972 10362 13996 10364
rect 14052 10362 14076 10364
rect 14132 10362 14138 10364
rect 13892 10310 13894 10362
rect 14074 10310 14076 10362
rect 13830 10308 13836 10310
rect 13892 10308 13916 10310
rect 13972 10308 13996 10310
rect 14052 10308 14076 10310
rect 14132 10308 14138 10310
rect 13830 10299 14138 10308
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13188 9042 13216 9318
rect 13280 9110 13308 9386
rect 13372 9353 13400 10066
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13464 9722 13492 9998
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13358 9344 13414 9353
rect 13358 9279 13414 9288
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13280 8022 13308 8230
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 13084 6384 13136 6390
rect 13084 6326 13136 6332
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13096 5234 13124 6326
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13004 4282 13032 4966
rect 13096 4622 13124 4966
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 12992 4276 13044 4282
rect 12992 4218 13044 4224
rect 12728 3454 12848 3482
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 12728 2990 12756 3454
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12256 2916 12308 2922
rect 12256 2858 12308 2864
rect 12268 2650 12296 2858
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12452 1902 12480 2790
rect 12728 2582 12756 2790
rect 12820 2774 12848 3334
rect 12912 2990 12940 3334
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12820 2746 12940 2774
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 12440 1896 12492 1902
rect 12440 1838 12492 1844
rect 12072 1828 12124 1834
rect 12072 1770 12124 1776
rect 12084 1562 12112 1770
rect 12072 1556 12124 1562
rect 12072 1498 12124 1504
rect 12820 814 12848 2586
rect 12912 1902 12940 2746
rect 13096 2650 13124 4558
rect 13372 3398 13400 9279
rect 13464 8974 13492 9658
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13556 8634 13584 8978
rect 13648 8634 13676 8978
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13556 5370 13584 6054
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13740 3738 13768 9930
rect 13830 9276 14138 9285
rect 13830 9274 13836 9276
rect 13892 9274 13916 9276
rect 13972 9274 13996 9276
rect 14052 9274 14076 9276
rect 14132 9274 14138 9276
rect 13892 9222 13894 9274
rect 14074 9222 14076 9274
rect 13830 9220 13836 9222
rect 13892 9220 13916 9222
rect 13972 9220 13996 9222
rect 14052 9220 14076 9222
rect 14132 9220 14138 9222
rect 13830 9211 14138 9220
rect 13830 8188 14138 8197
rect 13830 8186 13836 8188
rect 13892 8186 13916 8188
rect 13972 8186 13996 8188
rect 14052 8186 14076 8188
rect 14132 8186 14138 8188
rect 13892 8134 13894 8186
rect 14074 8134 14076 8186
rect 13830 8132 13836 8134
rect 13892 8132 13916 8134
rect 13972 8132 13996 8134
rect 14052 8132 14076 8134
rect 14132 8132 14138 8134
rect 13830 8123 14138 8132
rect 13820 7880 13872 7886
rect 13818 7848 13820 7857
rect 13872 7848 13874 7857
rect 13818 7783 13874 7792
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13832 7342 13860 7686
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13830 7100 14138 7109
rect 13830 7098 13836 7100
rect 13892 7098 13916 7100
rect 13972 7098 13996 7100
rect 14052 7098 14076 7100
rect 14132 7098 14138 7100
rect 13892 7046 13894 7098
rect 14074 7046 14076 7098
rect 13830 7044 13836 7046
rect 13892 7044 13916 7046
rect 13972 7044 13996 7046
rect 14052 7044 14076 7046
rect 14132 7044 14138 7046
rect 13830 7035 14138 7044
rect 14096 6860 14148 6866
rect 14200 6848 14228 11154
rect 14292 10554 14320 11750
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14384 11014 14412 11698
rect 14476 11150 14504 12174
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14384 10674 14412 10950
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14292 10526 14504 10554
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 14292 9178 14320 10134
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14292 8430 14320 8910
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14292 7750 14320 8366
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14148 6820 14228 6848
rect 14096 6802 14148 6808
rect 14108 6254 14136 6802
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14096 6248 14148 6254
rect 14148 6196 14228 6202
rect 14096 6190 14228 6196
rect 14108 6174 14228 6190
rect 13830 6012 14138 6021
rect 13830 6010 13836 6012
rect 13892 6010 13916 6012
rect 13972 6010 13996 6012
rect 14052 6010 14076 6012
rect 14132 6010 14138 6012
rect 13892 5958 13894 6010
rect 14074 5958 14076 6010
rect 13830 5956 13836 5958
rect 13892 5956 13916 5958
rect 13972 5956 13996 5958
rect 14052 5956 14076 5958
rect 14132 5956 14138 5958
rect 13830 5947 14138 5956
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14016 5778 14044 5850
rect 14200 5778 14228 6174
rect 14292 5778 14320 6598
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 13830 4924 14138 4933
rect 13830 4922 13836 4924
rect 13892 4922 13916 4924
rect 13972 4922 13996 4924
rect 14052 4922 14076 4924
rect 14132 4922 14138 4924
rect 13892 4870 13894 4922
rect 14074 4870 14076 4922
rect 13830 4868 13836 4870
rect 13892 4868 13916 4870
rect 13972 4868 13996 4870
rect 14052 4868 14076 4870
rect 14132 4868 14138 4870
rect 13830 4859 14138 4868
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 13830 3836 14138 3845
rect 13830 3834 13836 3836
rect 13892 3834 13916 3836
rect 13972 3834 13996 3836
rect 14052 3834 14076 3836
rect 14132 3834 14138 3836
rect 13892 3782 13894 3834
rect 14074 3782 14076 3834
rect 13830 3780 13836 3782
rect 13892 3780 13916 3782
rect 13972 3780 13996 3782
rect 14052 3780 14076 3782
rect 14132 3780 14138 3782
rect 13830 3771 14138 3780
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 13740 2582 13768 2994
rect 13830 2748 14138 2757
rect 13830 2746 13836 2748
rect 13892 2746 13916 2748
rect 13972 2746 13996 2748
rect 14052 2746 14076 2748
rect 14132 2746 14138 2748
rect 13892 2694 13894 2746
rect 14074 2694 14076 2746
rect 13830 2692 13836 2694
rect 13892 2692 13916 2694
rect 13972 2692 13996 2694
rect 14052 2692 14076 2694
rect 14132 2692 14138 2694
rect 13830 2683 14138 2692
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 14200 2378 14228 3946
rect 14292 3534 14320 3946
rect 14384 3738 14412 10406
rect 14476 9738 14504 10526
rect 14568 10266 14596 17070
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14844 16130 14872 16526
rect 14936 16250 14964 17600
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15120 16590 15148 16934
rect 15856 16794 15884 17734
rect 16210 17734 16528 17762
rect 16210 17600 16266 17734
rect 16500 17134 16528 17734
rect 16764 17604 16816 17610
rect 16854 17600 16910 18000
rect 17498 17762 17554 18000
rect 17498 17734 17816 17762
rect 17498 17600 17554 17734
rect 16764 17546 16816 17552
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 16776 16658 16804 17546
rect 16868 17134 16896 17600
rect 17188 17436 17496 17445
rect 17188 17434 17194 17436
rect 17250 17434 17274 17436
rect 17330 17434 17354 17436
rect 17410 17434 17434 17436
rect 17490 17434 17496 17436
rect 17250 17382 17252 17434
rect 17432 17382 17434 17434
rect 17188 17380 17194 17382
rect 17250 17380 17274 17382
rect 17330 17380 17354 17382
rect 17410 17380 17434 17382
rect 17490 17380 17496 17382
rect 17188 17371 17496 17380
rect 17788 17134 17816 17734
rect 18142 17600 18198 18000
rect 18786 17600 18842 18000
rect 19430 17600 19486 18000
rect 20074 17600 20130 18000
rect 20718 17600 20774 18000
rect 21362 17600 21418 18000
rect 22006 17600 22062 18000
rect 22650 17600 22706 18000
rect 23294 17600 23350 18000
rect 23938 17762 23994 18000
rect 23768 17734 23994 17762
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18984 17134 19012 17478
rect 19064 17264 19116 17270
rect 19064 17206 19116 17212
rect 19076 17134 19104 17206
rect 19444 17202 19472 17600
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 19522 17232 19578 17241
rect 19432 17196 19484 17202
rect 19522 17167 19578 17176
rect 19984 17196 20036 17202
rect 19432 17138 19484 17144
rect 19536 17134 19564 17167
rect 20168 17196 20220 17202
rect 20036 17156 20168 17184
rect 19984 17138 20036 17144
rect 20168 17138 20220 17144
rect 20364 17134 20392 17274
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20732 17134 20760 17206
rect 21376 17134 21404 17600
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 21364 17128 21416 17134
rect 22020 17116 22048 17600
rect 22664 17134 22692 17600
rect 23308 17134 23336 17600
rect 23768 17134 23796 17734
rect 23938 17600 23994 17734
rect 24582 17600 24638 18000
rect 25136 17604 25188 17610
rect 23904 17436 24212 17445
rect 23904 17434 23910 17436
rect 23966 17434 23990 17436
rect 24046 17434 24070 17436
rect 24126 17434 24150 17436
rect 24206 17434 24212 17436
rect 23966 17382 23968 17434
rect 24148 17382 24150 17434
rect 23904 17380 23910 17382
rect 23966 17380 23990 17382
rect 24046 17380 24070 17382
rect 24126 17380 24150 17382
rect 24206 17380 24212 17382
rect 23904 17371 24212 17380
rect 24032 17264 24084 17270
rect 24030 17232 24032 17241
rect 24084 17232 24086 17241
rect 24030 17167 24086 17176
rect 24596 17134 24624 17600
rect 25226 17600 25282 18000
rect 25870 17600 25926 18000
rect 26514 17762 26570 18000
rect 26252 17734 26570 17762
rect 25136 17546 25188 17552
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24688 17338 24716 17478
rect 25148 17338 25176 17546
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25240 17134 25268 17600
rect 25884 17202 25912 17600
rect 25872 17196 25924 17202
rect 25872 17138 25924 17144
rect 22284 17128 22336 17134
rect 22020 17088 22284 17116
rect 21364 17070 21416 17076
rect 22284 17070 22336 17076
rect 22652 17128 22704 17134
rect 22652 17070 22704 17076
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23756 17128 23808 17134
rect 23756 17070 23808 17076
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 25228 17128 25280 17134
rect 25228 17070 25280 17076
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 17592 16992 17644 16998
rect 17592 16934 17644 16940
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 17604 16726 17632 16934
rect 17592 16720 17644 16726
rect 17592 16662 17644 16668
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 14844 16102 14964 16130
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14660 11898 14688 15982
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14660 11121 14688 11494
rect 14646 11112 14702 11121
rect 14646 11047 14702 11056
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14476 9710 14596 9738
rect 14464 9648 14516 9654
rect 14462 9616 14464 9625
rect 14516 9616 14518 9625
rect 14462 9551 14518 9560
rect 14462 6896 14518 6905
rect 14568 6866 14596 9710
rect 14462 6831 14518 6840
rect 14556 6860 14608 6866
rect 14476 6798 14504 6831
rect 14556 6802 14608 6808
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14476 6458 14504 6734
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14476 5914 14504 6394
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14568 5846 14596 6802
rect 14556 5840 14608 5846
rect 14556 5782 14608 5788
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14476 5574 14504 5714
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14660 5370 14688 9998
rect 14752 6866 14780 15982
rect 14936 15910 14964 16102
rect 15120 16046 15148 16526
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14830 14512 14886 14521
rect 14830 14447 14832 14456
rect 14884 14447 14886 14456
rect 14832 14418 14884 14424
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14844 12782 14872 14214
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14936 12238 14964 15846
rect 15014 13424 15070 13433
rect 15014 13359 15016 13368
rect 15068 13359 15070 13368
rect 15016 13330 15068 13336
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 14922 11656 14978 11665
rect 14922 11591 14978 11600
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14844 10674 14872 11154
rect 14936 11150 14964 11591
rect 15028 11558 15056 12038
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14924 11144 14976 11150
rect 15120 11121 15148 13262
rect 14924 11086 14976 11092
rect 15106 11112 15162 11121
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14844 10062 14872 10610
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14936 6746 14964 11086
rect 15106 11047 15162 11056
rect 15120 10674 15148 11047
rect 15212 10810 15240 16594
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15488 15162 15516 15438
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15304 13870 15332 14214
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15488 13530 15516 14282
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15488 13161 15516 13262
rect 15474 13152 15530 13161
rect 15474 13087 15530 13096
rect 15488 12986 15516 13087
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15580 11898 15608 16594
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 16040 13870 16068 14418
rect 16132 14278 16160 14758
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16132 13870 16160 14214
rect 16408 14074 16436 14554
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 15752 13796 15804 13802
rect 15752 13738 15804 13744
rect 15764 13530 15792 13738
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 16210 13424 16266 13433
rect 16210 13359 16266 13368
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 15934 12336 15990 12345
rect 15934 12271 15936 12280
rect 15988 12271 15990 12280
rect 15936 12242 15988 12248
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15580 11614 15792 11642
rect 15580 11558 15608 11614
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 14752 6718 14964 6746
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14660 4758 14688 5170
rect 14648 4752 14700 4758
rect 14648 4694 14700 4700
rect 14660 4214 14688 4694
rect 14648 4208 14700 4214
rect 14568 4156 14648 4162
rect 14568 4150 14700 4156
rect 14568 4134 14688 4150
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14568 3534 14596 4134
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14568 2990 14596 3470
rect 14660 3126 14688 4014
rect 14648 3120 14700 3126
rect 14648 3062 14700 3068
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 14752 2774 14780 6718
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14936 5914 14964 6122
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 15028 5794 15056 10406
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 14936 5766 15056 5794
rect 14832 5092 14884 5098
rect 14832 5034 14884 5040
rect 14844 4486 14872 5034
rect 14936 4622 14964 5766
rect 15120 5370 15148 9998
rect 15212 7546 15240 10542
rect 15304 9586 15332 10542
rect 15396 10266 15424 10542
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15488 9110 15516 9862
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15304 4826 15332 6054
rect 15396 5302 15424 7686
rect 15580 6866 15608 11154
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15580 5302 15608 6598
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 15568 5296 15620 5302
rect 15568 5238 15620 5244
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14476 2746 14780 2774
rect 14844 2774 14872 4218
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 15028 4078 15056 4150
rect 15212 4146 15240 4626
rect 15304 4554 15332 4762
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 15304 4282 15332 4490
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 15028 3058 15056 4014
rect 15396 3992 15424 5102
rect 15488 4826 15516 5102
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15580 4690 15608 5238
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15568 4004 15620 4010
rect 15396 3964 15568 3992
rect 15568 3946 15620 3952
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15212 3670 15240 3878
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15120 3194 15148 3538
rect 15672 3194 15700 11494
rect 15764 11150 15792 11614
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 15764 9654 15792 10474
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15750 9480 15806 9489
rect 15750 9415 15752 9424
rect 15804 9415 15806 9424
rect 15752 9386 15804 9392
rect 15856 9058 15884 12038
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 15948 10266 15976 10474
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 16040 9722 16068 12038
rect 16132 11694 16160 12718
rect 16224 12442 16252 13359
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16394 12336 16450 12345
rect 16394 12271 16450 12280
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 15764 9030 15884 9058
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 15764 2774 15792 9030
rect 15948 7546 15976 9386
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16040 8430 16068 9318
rect 16132 8634 16160 9454
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16040 6662 16068 7278
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 15844 6384 15896 6390
rect 15844 6326 15896 6332
rect 15856 5778 15884 6326
rect 16040 6118 16068 6598
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15948 5166 15976 5510
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15856 4010 15884 4626
rect 15948 4282 15976 5102
rect 16132 4486 16160 5102
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 16224 4298 16252 11086
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16316 8498 16344 8910
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16316 7410 16344 8434
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16316 6322 16344 7346
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16408 6254 16436 12271
rect 16592 11257 16620 16594
rect 17188 16348 17496 16357
rect 17188 16346 17194 16348
rect 17250 16346 17274 16348
rect 17330 16346 17354 16348
rect 17410 16346 17434 16348
rect 17490 16346 17496 16348
rect 17250 16294 17252 16346
rect 17432 16294 17434 16346
rect 17188 16292 17194 16294
rect 17250 16292 17274 16294
rect 17330 16292 17354 16294
rect 17410 16292 17434 16294
rect 17490 16292 17496 16294
rect 17188 16283 17496 16292
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16684 14958 16712 15506
rect 17052 15162 17080 15982
rect 17188 15260 17496 15269
rect 17188 15258 17194 15260
rect 17250 15258 17274 15260
rect 17330 15258 17354 15260
rect 17410 15258 17434 15260
rect 17490 15258 17496 15260
rect 17250 15206 17252 15258
rect 17432 15206 17434 15258
rect 17188 15204 17194 15206
rect 17250 15204 17274 15206
rect 17330 15204 17354 15206
rect 17410 15204 17434 15206
rect 17490 15204 17496 15206
rect 17188 15195 17496 15204
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16684 14006 16712 14350
rect 16960 14278 16988 14894
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16672 13864 16724 13870
rect 16960 13818 16988 14214
rect 17052 14006 17080 15098
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17188 14172 17496 14181
rect 17188 14170 17194 14172
rect 17250 14170 17274 14172
rect 17330 14170 17354 14172
rect 17410 14170 17434 14172
rect 17490 14170 17496 14172
rect 17250 14118 17252 14170
rect 17432 14118 17434 14170
rect 17188 14116 17194 14118
rect 17250 14116 17274 14118
rect 17330 14116 17354 14118
rect 17410 14116 17434 14118
rect 17490 14116 17496 14118
rect 17188 14107 17496 14116
rect 17040 14000 17092 14006
rect 17040 13942 17092 13948
rect 17040 13864 17092 13870
rect 16724 13812 16896 13818
rect 16672 13806 16896 13812
rect 16684 13790 16896 13806
rect 16960 13812 17040 13818
rect 16960 13806 17092 13812
rect 16960 13790 17080 13806
rect 17604 13802 17632 14214
rect 16868 13716 16896 13790
rect 16868 13688 16988 13716
rect 16960 13326 16988 13688
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16684 12374 16712 13262
rect 16960 12986 16988 13262
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17052 12764 17080 13790
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17592 13796 17644 13802
rect 17592 13738 17644 13744
rect 17236 13326 17264 13738
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17188 13084 17496 13093
rect 17188 13082 17194 13084
rect 17250 13082 17274 13084
rect 17330 13082 17354 13084
rect 17410 13082 17434 13084
rect 17490 13082 17496 13084
rect 17250 13030 17252 13082
rect 17432 13030 17434 13082
rect 17188 13028 17194 13030
rect 17250 13028 17274 13030
rect 17330 13028 17354 13030
rect 17410 13028 17434 13030
rect 17490 13028 17496 13030
rect 17188 13019 17496 13028
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17132 12776 17184 12782
rect 17052 12736 17132 12764
rect 17132 12718 17184 12724
rect 16948 12708 17000 12714
rect 16948 12650 17000 12656
rect 16960 12442 16988 12650
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 17328 12306 17356 12922
rect 17604 12442 17632 13126
rect 17592 12436 17644 12442
rect 17788 12434 17816 16934
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18340 15638 18368 15982
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 17880 14618 17908 14826
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17972 12850 18000 13806
rect 18064 13530 18092 14350
rect 18156 13530 18184 14554
rect 18248 13938 18276 14826
rect 18340 14482 18368 15574
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18248 13462 18276 13874
rect 18340 13870 18368 14418
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 18328 13388 18380 13394
rect 18328 13330 18380 13336
rect 18064 12986 18092 13330
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17592 12378 17644 12384
rect 17696 12406 17816 12434
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17592 12164 17644 12170
rect 17592 12106 17644 12112
rect 17188 11996 17496 12005
rect 17188 11994 17194 11996
rect 17250 11994 17274 11996
rect 17330 11994 17354 11996
rect 17410 11994 17434 11996
rect 17490 11994 17496 11996
rect 17250 11942 17252 11994
rect 17432 11942 17434 11994
rect 17188 11940 17194 11942
rect 17250 11940 17274 11942
rect 17330 11940 17354 11942
rect 17410 11940 17434 11942
rect 17490 11940 17496 11942
rect 17188 11931 17496 11940
rect 17604 11898 17632 12106
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17144 11558 17172 11630
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 16578 11248 16634 11257
rect 16578 11183 16634 11192
rect 16960 11150 16988 11494
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16960 10810 16988 11086
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16684 10130 16712 10406
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16592 9654 16620 10066
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16868 9518 16896 10066
rect 17052 9926 17080 11494
rect 17144 11218 17172 11494
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17188 10908 17496 10917
rect 17188 10906 17194 10908
rect 17250 10906 17274 10908
rect 17330 10906 17354 10908
rect 17410 10906 17434 10908
rect 17490 10906 17496 10908
rect 17250 10854 17252 10906
rect 17432 10854 17434 10906
rect 17188 10852 17194 10854
rect 17250 10852 17274 10854
rect 17330 10852 17354 10854
rect 17410 10852 17434 10854
rect 17490 10852 17496 10854
rect 17188 10843 17496 10852
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17328 10266 17356 10406
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17604 10130 17632 10950
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17040 9920 17092 9926
rect 16960 9868 17040 9874
rect 16960 9862 17092 9868
rect 16960 9846 17080 9862
rect 16960 9586 16988 9846
rect 17188 9820 17496 9829
rect 17188 9818 17194 9820
rect 17250 9818 17274 9820
rect 17330 9818 17354 9820
rect 17410 9818 17434 9820
rect 17490 9818 17496 9820
rect 17250 9766 17252 9818
rect 17432 9766 17434 9818
rect 17188 9764 17194 9766
rect 17250 9764 17274 9766
rect 17330 9764 17354 9766
rect 17410 9764 17434 9766
rect 17490 9764 17496 9766
rect 17188 9755 17496 9764
rect 17604 9654 17632 10066
rect 17592 9648 17644 9654
rect 17052 9586 17264 9602
rect 17592 9590 17644 9596
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 17052 9580 17276 9586
rect 17052 9574 17224 9580
rect 16856 9512 16908 9518
rect 17052 9466 17080 9574
rect 17224 9522 17276 9528
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 16856 9454 16908 9460
rect 16960 9438 17080 9466
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 16578 9072 16634 9081
rect 16578 9007 16634 9016
rect 16764 9036 16816 9042
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 16132 4270 16252 4298
rect 16304 4276 16356 4282
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15844 4004 15896 4010
rect 15844 3946 15896 3952
rect 15948 3738 15976 4014
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 16040 3194 16068 3878
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 14844 2746 14964 2774
rect 15764 2746 15884 2774
rect 14476 2666 14504 2746
rect 14384 2638 14504 2666
rect 14646 2680 14702 2689
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 13912 2304 13964 2310
rect 13912 2246 13964 2252
rect 13924 1902 13952 2246
rect 14384 1902 14412 2638
rect 14646 2615 14648 2624
rect 14700 2615 14702 2624
rect 14648 2586 14700 2592
rect 14936 2582 14964 2746
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 12900 1896 12952 1902
rect 12900 1838 12952 1844
rect 13912 1896 13964 1902
rect 13912 1838 13964 1844
rect 14372 1896 14424 1902
rect 14372 1838 14424 1844
rect 12992 1828 13044 1834
rect 12992 1770 13044 1776
rect 12900 1760 12952 1766
rect 12900 1702 12952 1708
rect 12912 1494 12940 1702
rect 12900 1488 12952 1494
rect 12900 1430 12952 1436
rect 13004 1018 13032 1770
rect 13830 1660 14138 1669
rect 13830 1658 13836 1660
rect 13892 1658 13916 1660
rect 13972 1658 13996 1660
rect 14052 1658 14076 1660
rect 14132 1658 14138 1660
rect 13892 1606 13894 1658
rect 14074 1606 14076 1658
rect 13830 1604 13836 1606
rect 13892 1604 13916 1606
rect 13972 1604 13996 1606
rect 14052 1604 14076 1606
rect 14132 1604 14138 1606
rect 13830 1595 14138 1604
rect 14476 1358 14504 2450
rect 15028 2038 15056 2450
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 15016 2032 15068 2038
rect 15016 1974 15068 1980
rect 15292 2032 15344 2038
rect 15292 1974 15344 1980
rect 14556 1896 14608 1902
rect 14556 1838 14608 1844
rect 15016 1896 15068 1902
rect 15068 1856 15240 1884
rect 15304 1873 15332 1974
rect 15396 1902 15424 2382
rect 15384 1896 15436 1902
rect 15016 1838 15068 1844
rect 14568 1426 14596 1838
rect 15212 1426 15240 1856
rect 15290 1864 15346 1873
rect 15384 1838 15436 1844
rect 15290 1799 15346 1808
rect 15396 1494 15424 1838
rect 15660 1760 15712 1766
rect 15660 1702 15712 1708
rect 15384 1488 15436 1494
rect 15384 1430 15436 1436
rect 14556 1420 14608 1426
rect 14556 1362 14608 1368
rect 15200 1420 15252 1426
rect 15200 1362 15252 1368
rect 14096 1352 14148 1358
rect 14096 1294 14148 1300
rect 14464 1352 14516 1358
rect 14464 1294 14516 1300
rect 14108 1018 14136 1294
rect 14832 1216 14884 1222
rect 14832 1158 14884 1164
rect 12992 1012 13044 1018
rect 12992 954 13044 960
rect 14096 1012 14148 1018
rect 14096 954 14148 960
rect 13004 814 13032 954
rect 13084 944 13136 950
rect 13084 886 13136 892
rect 11980 808 12032 814
rect 11980 750 12032 756
rect 12808 808 12860 814
rect 12808 750 12860 756
rect 12992 808 13044 814
rect 12992 750 13044 756
rect 11612 672 11664 678
rect 11612 614 11664 620
rect 13096 400 13124 886
rect 13830 572 14138 581
rect 13830 570 13836 572
rect 13892 570 13916 572
rect 13972 570 13996 572
rect 14052 570 14076 572
rect 14132 570 14138 572
rect 13892 518 13894 570
rect 14074 518 14076 570
rect 13830 516 13836 518
rect 13892 516 13916 518
rect 13972 516 13996 518
rect 14052 516 14076 518
rect 14132 516 14138 518
rect 13830 507 14138 516
rect 14844 400 14872 1158
rect 15672 814 15700 1702
rect 15856 1426 15884 2746
rect 16040 1766 16068 2926
rect 16132 2922 16160 4270
rect 16304 4218 16356 4224
rect 16316 4078 16344 4218
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16212 4004 16264 4010
rect 16212 3946 16264 3952
rect 16224 3398 16252 3946
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16316 3602 16344 3878
rect 16408 3602 16436 4558
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 16316 3058 16344 3538
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16408 2990 16436 3334
rect 16396 2984 16448 2990
rect 16396 2926 16448 2932
rect 16120 2916 16172 2922
rect 16120 2858 16172 2864
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16028 1760 16080 1766
rect 16028 1702 16080 1708
rect 16316 1426 16344 2382
rect 16500 1766 16528 6054
rect 16592 5846 16620 9007
rect 16764 8978 16816 8984
rect 16776 8634 16804 8978
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 16960 5681 16988 9438
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17052 8430 17080 9318
rect 17144 9081 17172 9454
rect 17512 9450 17540 9522
rect 17500 9444 17552 9450
rect 17552 9404 17632 9432
rect 17500 9386 17552 9392
rect 17130 9072 17186 9081
rect 17130 9007 17186 9016
rect 17188 8732 17496 8741
rect 17188 8730 17194 8732
rect 17250 8730 17274 8732
rect 17330 8730 17354 8732
rect 17410 8730 17434 8732
rect 17490 8730 17496 8732
rect 17250 8678 17252 8730
rect 17432 8678 17434 8730
rect 17188 8676 17194 8678
rect 17250 8676 17274 8678
rect 17330 8676 17354 8678
rect 17410 8676 17434 8678
rect 17490 8676 17496 8678
rect 17188 8667 17496 8676
rect 17604 8616 17632 9404
rect 17420 8588 17632 8616
rect 17420 8430 17448 8588
rect 17590 8528 17646 8537
rect 17590 8463 17646 8472
rect 17604 8430 17632 8463
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17420 7818 17448 8366
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17188 7644 17496 7653
rect 17188 7642 17194 7644
rect 17250 7642 17274 7644
rect 17330 7642 17354 7644
rect 17410 7642 17434 7644
rect 17490 7642 17496 7644
rect 17250 7590 17252 7642
rect 17432 7590 17434 7642
rect 17188 7588 17194 7590
rect 17250 7588 17274 7590
rect 17330 7588 17354 7590
rect 17410 7588 17434 7590
rect 17490 7588 17496 7590
rect 17188 7579 17496 7588
rect 17188 6556 17496 6565
rect 17188 6554 17194 6556
rect 17250 6554 17274 6556
rect 17330 6554 17354 6556
rect 17410 6554 17434 6556
rect 17490 6554 17496 6556
rect 17250 6502 17252 6554
rect 17432 6502 17434 6554
rect 17188 6500 17194 6502
rect 17250 6500 17274 6502
rect 17330 6500 17354 6502
rect 17410 6500 17434 6502
rect 17490 6500 17496 6502
rect 17188 6491 17496 6500
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 17052 5914 17080 6190
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17500 5840 17552 5846
rect 17552 5800 17632 5828
rect 17500 5782 17552 5788
rect 17316 5704 17368 5710
rect 16946 5672 17002 5681
rect 16946 5607 17002 5616
rect 17314 5672 17316 5681
rect 17368 5672 17370 5681
rect 17604 5642 17632 5800
rect 17314 5607 17370 5616
rect 17592 5636 17644 5642
rect 17328 5574 17356 5607
rect 17592 5578 17644 5584
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 17188 5468 17496 5477
rect 17188 5466 17194 5468
rect 17250 5466 17274 5468
rect 17330 5466 17354 5468
rect 17410 5466 17434 5468
rect 17490 5466 17496 5468
rect 17250 5414 17252 5466
rect 17432 5414 17434 5466
rect 17188 5412 17194 5414
rect 17250 5412 17274 5414
rect 17330 5412 17354 5414
rect 17410 5412 17434 5414
rect 17490 5412 17496 5414
rect 17188 5403 17496 5412
rect 16856 5296 16908 5302
rect 16856 5238 16908 5244
rect 16868 5166 16896 5238
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16592 3602 16620 4014
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16592 3398 16620 3538
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16684 2774 16712 4694
rect 16868 4078 16896 5102
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17144 4690 17172 4966
rect 17696 4842 17724 12406
rect 18156 11898 18184 13330
rect 18340 12306 18368 13330
rect 18328 12300 18380 12306
rect 18328 12242 18380 12248
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18064 11354 18092 11630
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17788 9178 17816 9998
rect 17880 9994 17908 10542
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17972 8838 18000 9454
rect 18064 9382 18092 11018
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18248 9722 18276 9998
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 18064 9110 18092 9318
rect 18052 9104 18104 9110
rect 18052 9046 18104 9052
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17776 8560 17828 8566
rect 17776 8502 17828 8508
rect 17788 8401 17816 8502
rect 17774 8392 17830 8401
rect 17972 8362 18000 8774
rect 17960 8356 18012 8362
rect 17830 8336 17908 8344
rect 17774 8327 17908 8336
rect 17788 8316 17908 8327
rect 17880 8242 17908 8316
rect 17960 8298 18012 8304
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 18064 8242 18092 8298
rect 17880 8214 18092 8242
rect 17972 6662 18000 8214
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 17328 4814 17724 4842
rect 17328 4758 17356 4814
rect 17972 4758 18000 6190
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 18064 5914 18092 6054
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4758 18276 4966
rect 17316 4752 17368 4758
rect 17316 4694 17368 4700
rect 17960 4752 18012 4758
rect 17960 4694 18012 4700
rect 18236 4752 18288 4758
rect 18236 4694 18288 4700
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 17188 4380 17496 4389
rect 17188 4378 17194 4380
rect 17250 4378 17274 4380
rect 17330 4378 17354 4380
rect 17410 4378 17434 4380
rect 17490 4378 17496 4380
rect 17250 4326 17252 4378
rect 17432 4326 17434 4378
rect 17188 4324 17194 4326
rect 17250 4324 17274 4326
rect 17330 4324 17354 4326
rect 17410 4324 17434 4326
rect 17490 4324 17496 4326
rect 17188 4315 17496 4324
rect 17776 4208 17828 4214
rect 17776 4150 17828 4156
rect 17788 4078 17816 4150
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17788 3602 17816 4014
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17052 2990 17080 3334
rect 17188 3292 17496 3301
rect 17188 3290 17194 3292
rect 17250 3290 17274 3292
rect 17330 3290 17354 3292
rect 17410 3290 17434 3292
rect 17490 3290 17496 3292
rect 17250 3238 17252 3290
rect 17432 3238 17434 3290
rect 17188 3236 17194 3238
rect 17250 3236 17274 3238
rect 17330 3236 17354 3238
rect 17410 3236 17434 3238
rect 17490 3236 17496 3238
rect 17188 3227 17496 3236
rect 17788 3058 17816 3538
rect 17972 3482 18000 4694
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18340 3670 18368 3878
rect 18328 3664 18380 3670
rect 18328 3606 18380 3612
rect 17880 3454 18000 3482
rect 18052 3460 18104 3466
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 16592 2746 16712 2774
rect 16592 2582 16620 2746
rect 16580 2576 16632 2582
rect 16580 2518 16632 2524
rect 16776 2514 16804 2790
rect 17236 2514 17264 2790
rect 16764 2508 16816 2514
rect 16764 2450 16816 2456
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 16764 1896 16816 1902
rect 16764 1838 16816 1844
rect 16396 1760 16448 1766
rect 16396 1702 16448 1708
rect 16488 1760 16540 1766
rect 16488 1702 16540 1708
rect 15844 1420 15896 1426
rect 15844 1362 15896 1368
rect 16304 1420 16356 1426
rect 16304 1362 16356 1368
rect 16118 912 16174 921
rect 16118 847 16174 856
rect 16132 814 16160 847
rect 16316 814 16344 1362
rect 16408 814 16436 1702
rect 16500 814 16528 1702
rect 16776 1358 16804 1838
rect 16960 1834 16988 2246
rect 16948 1828 17000 1834
rect 16948 1770 17000 1776
rect 17052 1494 17080 2246
rect 17188 2204 17496 2213
rect 17188 2202 17194 2204
rect 17250 2202 17274 2204
rect 17330 2202 17354 2204
rect 17410 2202 17434 2204
rect 17490 2202 17496 2204
rect 17250 2150 17252 2202
rect 17432 2150 17434 2202
rect 17188 2148 17194 2150
rect 17250 2148 17274 2150
rect 17330 2148 17354 2150
rect 17410 2148 17434 2150
rect 17490 2148 17496 2150
rect 17188 2139 17496 2148
rect 17880 1902 17908 3454
rect 18052 3402 18104 3408
rect 17868 1896 17920 1902
rect 17868 1838 17920 1844
rect 17960 1828 18012 1834
rect 17960 1770 18012 1776
rect 17972 1562 18000 1770
rect 18064 1562 18092 3402
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18340 2990 18368 3334
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18432 2009 18460 16934
rect 19076 16658 19104 17070
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 24676 17060 24728 17066
rect 24676 17002 24728 17008
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 19352 16697 19380 16934
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19338 16688 19394 16697
rect 19064 16652 19116 16658
rect 19812 16658 19840 16730
rect 19904 16697 19932 16934
rect 19890 16688 19946 16697
rect 19338 16623 19394 16632
rect 19616 16652 19668 16658
rect 19064 16594 19116 16600
rect 19616 16594 19668 16600
rect 19800 16652 19852 16658
rect 19890 16623 19946 16632
rect 19800 16594 19852 16600
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18524 15706 18552 16526
rect 19628 16454 19656 16594
rect 19064 16448 19116 16454
rect 19064 16390 19116 16396
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18892 14958 18920 15846
rect 19076 15570 19104 16390
rect 19628 15570 19656 16390
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19076 15162 19104 15506
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 19064 14952 19116 14958
rect 19168 14940 19196 15438
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19260 14958 19288 15302
rect 19812 15026 19840 16594
rect 19892 15428 19944 15434
rect 19892 15370 19944 15376
rect 19904 15162 19932 15370
rect 19892 15156 19944 15162
rect 19892 15098 19944 15104
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19116 14912 19196 14940
rect 19248 14952 19300 14958
rect 19064 14894 19116 14900
rect 19248 14894 19300 14900
rect 18616 14278 18644 14894
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18800 14618 18828 14826
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 19076 14482 19104 14894
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18524 13954 18552 14214
rect 18616 14074 18644 14214
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18524 13926 18644 13954
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18524 11354 18552 13806
rect 18616 13802 18644 13926
rect 19260 13802 19288 14894
rect 19432 14816 19484 14822
rect 19996 14770 20024 16934
rect 20546 16892 20854 16901
rect 20546 16890 20552 16892
rect 20608 16890 20632 16892
rect 20688 16890 20712 16892
rect 20768 16890 20792 16892
rect 20848 16890 20854 16892
rect 20608 16838 20610 16890
rect 20790 16838 20792 16890
rect 20546 16836 20552 16838
rect 20608 16836 20632 16838
rect 20688 16836 20712 16838
rect 20768 16836 20792 16838
rect 20848 16836 20854 16838
rect 20546 16827 20854 16836
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20732 16114 20760 16662
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20916 15910 20944 16526
rect 21364 16448 21416 16454
rect 21364 16390 21416 16396
rect 21376 16046 21404 16390
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 21364 16040 21416 16046
rect 21364 15982 21416 15988
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20546 15804 20854 15813
rect 20546 15802 20552 15804
rect 20608 15802 20632 15804
rect 20688 15802 20712 15804
rect 20768 15802 20792 15804
rect 20848 15802 20854 15804
rect 20608 15750 20610 15802
rect 20790 15750 20792 15802
rect 20546 15748 20552 15750
rect 20608 15748 20632 15750
rect 20688 15748 20712 15750
rect 20768 15748 20792 15750
rect 20848 15748 20854 15750
rect 20546 15739 20854 15748
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 19432 14758 19484 14764
rect 19444 14550 19472 14758
rect 19628 14742 20024 14770
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19536 13870 19564 14214
rect 19524 13864 19576 13870
rect 19338 13832 19394 13841
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 19248 13796 19300 13802
rect 19524 13806 19576 13812
rect 19338 13767 19394 13776
rect 19248 13738 19300 13744
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18616 11218 18644 13738
rect 19352 13462 19380 13767
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19444 13394 19472 13670
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18708 12306 18736 12786
rect 18984 12374 19012 13126
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 18972 12368 19024 12374
rect 18972 12310 19024 12316
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18616 9654 18644 11154
rect 18708 10674 18736 12242
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18984 11830 19012 12038
rect 18972 11824 19024 11830
rect 18786 11792 18842 11801
rect 18972 11766 19024 11772
rect 18786 11727 18842 11736
rect 18800 11694 18828 11727
rect 19444 11694 19472 12582
rect 19536 11694 19564 13806
rect 18788 11688 18840 11694
rect 19340 11688 19392 11694
rect 18788 11630 18840 11636
rect 19338 11656 19340 11665
rect 19432 11688 19484 11694
rect 19392 11656 19394 11665
rect 19432 11630 19484 11636
rect 19524 11688 19576 11694
rect 19524 11630 19576 11636
rect 19338 11591 19394 11600
rect 18972 11552 19024 11558
rect 19024 11500 19564 11506
rect 18972 11494 19564 11500
rect 18984 11478 19564 11494
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18708 10130 18736 10610
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18800 9178 18828 11154
rect 18892 11121 18920 11154
rect 19260 11121 19288 11290
rect 19432 11280 19484 11286
rect 19432 11222 19484 11228
rect 18878 11112 18934 11121
rect 18878 11047 18934 11056
rect 19246 11112 19302 11121
rect 19246 11047 19302 11056
rect 19260 10418 19288 11047
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19352 10606 19380 10950
rect 19444 10606 19472 11222
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19260 10390 19380 10418
rect 19352 9518 19380 10390
rect 19536 10010 19564 11478
rect 19444 9982 19564 10010
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18800 7546 18828 8978
rect 19444 8634 19472 9982
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19536 9586 19564 9862
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19536 8430 19564 8774
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19524 8424 19576 8430
rect 19524 8366 19576 8372
rect 19352 7750 19380 8366
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18696 7336 18748 7342
rect 18696 7278 18748 7284
rect 18604 7200 18656 7206
rect 18708 7188 18736 7278
rect 18656 7160 18736 7188
rect 18604 7142 18656 7148
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18524 6322 18552 6802
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18708 6746 18736 7160
rect 18800 6934 18828 7482
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 18892 7002 18920 7278
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 18788 6928 18840 6934
rect 18788 6870 18840 6876
rect 18788 6792 18840 6798
rect 18708 6740 18788 6746
rect 18708 6734 18840 6740
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18524 5710 18552 6258
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18616 5098 18644 6734
rect 18708 6718 18828 6734
rect 19352 6730 19380 7278
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19340 6724 19392 6730
rect 18708 6458 18736 6718
rect 19340 6666 19392 6672
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18708 5778 18736 6394
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 18880 6180 18932 6186
rect 18880 6122 18932 6128
rect 18892 5914 18920 6122
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18788 5636 18840 5642
rect 18788 5578 18840 5584
rect 18800 5302 18828 5578
rect 18788 5296 18840 5302
rect 18788 5238 18840 5244
rect 18800 5166 18828 5238
rect 18892 5166 18920 5850
rect 19260 5778 19288 6190
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18880 5160 18932 5166
rect 18880 5102 18932 5108
rect 19352 5098 19380 6258
rect 19444 5234 19472 6734
rect 19536 6390 19564 7142
rect 19524 6384 19576 6390
rect 19524 6326 19576 6332
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18984 4162 19012 4626
rect 19248 4480 19300 4486
rect 19248 4422 19300 4428
rect 18984 4146 19196 4162
rect 18984 4140 19208 4146
rect 18984 4134 19156 4140
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18524 3602 18552 3878
rect 18800 3738 18828 3878
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 19076 3602 19104 4134
rect 19156 4082 19208 4088
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 3194 18644 3334
rect 19076 3194 19104 3538
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 18418 2000 18474 2009
rect 18418 1935 18474 1944
rect 18512 1964 18564 1970
rect 18432 1902 18460 1935
rect 18512 1906 18564 1912
rect 18420 1896 18472 1902
rect 18420 1838 18472 1844
rect 18420 1760 18472 1766
rect 18524 1748 18552 1906
rect 18880 1896 18932 1902
rect 18880 1838 18932 1844
rect 18472 1720 18552 1748
rect 18420 1702 18472 1708
rect 17960 1556 18012 1562
rect 17960 1498 18012 1504
rect 18052 1556 18104 1562
rect 18052 1498 18104 1504
rect 17040 1488 17092 1494
rect 17040 1430 17092 1436
rect 18432 1426 18460 1702
rect 18892 1426 18920 1838
rect 18970 1456 19026 1465
rect 18420 1420 18472 1426
rect 18420 1362 18472 1368
rect 18880 1420 18932 1426
rect 19260 1426 19288 4422
rect 18970 1391 18972 1400
rect 18880 1362 18932 1368
rect 19024 1391 19026 1400
rect 19248 1420 19300 1426
rect 18972 1362 19024 1368
rect 19248 1362 19300 1368
rect 16764 1352 16816 1358
rect 16764 1294 16816 1300
rect 16580 944 16632 950
rect 16580 886 16632 892
rect 15660 808 15712 814
rect 15660 750 15712 756
rect 16120 808 16172 814
rect 16120 750 16172 756
rect 16304 808 16356 814
rect 16304 750 16356 756
rect 16396 808 16448 814
rect 16396 750 16448 756
rect 16488 808 16540 814
rect 16488 750 16540 756
rect 16592 400 16620 886
rect 16776 882 16804 1294
rect 18328 1216 18380 1222
rect 18328 1158 18380 1164
rect 17188 1116 17496 1125
rect 17188 1114 17194 1116
rect 17250 1114 17274 1116
rect 17330 1114 17354 1116
rect 17410 1114 17434 1116
rect 17490 1114 17496 1116
rect 17250 1062 17252 1114
rect 17432 1062 17434 1114
rect 17188 1060 17194 1062
rect 17250 1060 17274 1062
rect 17330 1060 17354 1062
rect 17410 1060 17434 1062
rect 17490 1060 17496 1062
rect 17188 1051 17496 1060
rect 16764 876 16816 882
rect 16764 818 16816 824
rect 18340 400 18368 1158
rect 19628 950 19656 14742
rect 20088 14618 20116 15438
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20260 15020 20312 15026
rect 20260 14962 20312 14968
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19812 12374 19840 13806
rect 19800 12368 19852 12374
rect 19800 12310 19852 12316
rect 19904 11898 19932 13806
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19996 12442 20024 13330
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 19892 11688 19944 11694
rect 19890 11656 19892 11665
rect 19944 11656 19946 11665
rect 19800 11620 19852 11626
rect 19890 11591 19946 11600
rect 19800 11562 19852 11568
rect 19812 11354 19840 11562
rect 19708 11348 19760 11354
rect 19708 11290 19760 11296
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19720 11234 19748 11290
rect 19892 11280 19944 11286
rect 19720 11228 19892 11234
rect 19720 11222 19944 11228
rect 19720 11206 19932 11222
rect 19996 10810 20024 12242
rect 20088 12170 20116 14350
rect 20180 14074 20208 14894
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20272 13870 20300 14962
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 20628 14952 20680 14958
rect 20732 14940 20760 15302
rect 20916 15026 20944 15846
rect 21100 15026 21128 15982
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 20680 14912 20760 14940
rect 20628 14894 20680 14900
rect 20364 14550 20392 14894
rect 20732 14804 20760 14912
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20732 14776 20944 14804
rect 20546 14716 20854 14725
rect 20546 14714 20552 14716
rect 20608 14714 20632 14716
rect 20688 14714 20712 14716
rect 20768 14714 20792 14716
rect 20848 14714 20854 14716
rect 20608 14662 20610 14714
rect 20790 14662 20792 14714
rect 20546 14660 20552 14662
rect 20608 14660 20632 14662
rect 20688 14660 20712 14662
rect 20768 14660 20792 14662
rect 20848 14660 20854 14662
rect 20546 14651 20854 14660
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 20352 14544 20404 14550
rect 20352 14486 20404 14492
rect 20628 14476 20680 14482
rect 20548 14436 20628 14464
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 20272 12782 20300 13670
rect 20364 12866 20392 14214
rect 20548 13870 20576 14436
rect 20628 14418 20680 14424
rect 20536 13864 20588 13870
rect 20720 13864 20772 13870
rect 20536 13806 20588 13812
rect 20718 13832 20720 13841
rect 20772 13832 20774 13841
rect 20548 13716 20576 13806
rect 20718 13767 20774 13776
rect 20824 13734 20852 14554
rect 20916 14006 20944 14776
rect 21008 14618 21036 14894
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 21192 13870 21220 14758
rect 21284 14260 21312 15506
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21376 14618 21404 15438
rect 21468 14770 21496 16934
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22100 16516 22152 16522
rect 22100 16458 22152 16464
rect 22112 15706 22140 16458
rect 22664 16250 22692 16594
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 22284 16040 22336 16046
rect 22940 15994 22968 16050
rect 22284 15982 22336 15988
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22296 15570 22324 15982
rect 22756 15966 22968 15994
rect 22468 15632 22520 15638
rect 22468 15574 22520 15580
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22100 15360 22152 15366
rect 22100 15302 22152 15308
rect 21732 14952 21784 14958
rect 21652 14912 21732 14940
rect 21468 14742 21588 14770
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21364 14272 21416 14278
rect 21284 14232 21364 14260
rect 21364 14214 21416 14220
rect 21376 13870 21404 14214
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 20456 13688 20576 13716
rect 20812 13728 20864 13734
rect 20456 12986 20484 13688
rect 20812 13670 20864 13676
rect 20546 13628 20854 13637
rect 20546 13626 20552 13628
rect 20608 13626 20632 13628
rect 20688 13626 20712 13628
rect 20768 13626 20792 13628
rect 20848 13626 20854 13628
rect 20608 13574 20610 13626
rect 20790 13574 20792 13626
rect 20546 13572 20552 13574
rect 20608 13572 20632 13574
rect 20688 13572 20712 13574
rect 20768 13572 20792 13574
rect 20848 13572 20854 13574
rect 20546 13563 20854 13572
rect 21100 13530 21128 13806
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20364 12838 20484 12866
rect 21100 12850 21128 13466
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20272 12646 20300 12718
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20364 12306 20392 12582
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 20456 11694 20484 12838
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 20546 12540 20854 12549
rect 20546 12538 20552 12540
rect 20608 12538 20632 12540
rect 20688 12538 20712 12540
rect 20768 12538 20792 12540
rect 20848 12538 20854 12540
rect 20608 12486 20610 12538
rect 20790 12486 20792 12538
rect 20546 12484 20552 12486
rect 20608 12484 20632 12486
rect 20688 12484 20712 12486
rect 20768 12484 20792 12486
rect 20848 12484 20854 12486
rect 20546 12475 20854 12484
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 20548 11898 20576 12242
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 21192 11694 21220 13330
rect 21284 12434 21312 13806
rect 21284 12406 21496 12434
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 9518 19932 10406
rect 20272 10266 20300 11494
rect 20546 11452 20854 11461
rect 20546 11450 20552 11452
rect 20608 11450 20632 11452
rect 20688 11450 20712 11452
rect 20768 11450 20792 11452
rect 20848 11450 20854 11452
rect 20608 11398 20610 11450
rect 20790 11398 20792 11450
rect 20546 11396 20552 11398
rect 20608 11396 20632 11398
rect 20688 11396 20712 11398
rect 20768 11396 20792 11398
rect 20848 11396 20854 11398
rect 20546 11387 20854 11396
rect 21284 11354 21312 12174
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21376 11626 21404 12038
rect 21468 11898 21496 12406
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21364 11620 21416 11626
rect 21364 11562 21416 11568
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21468 11218 21496 11834
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 21456 11212 21508 11218
rect 21456 11154 21508 11160
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20180 9518 20208 9998
rect 20456 9654 20484 11154
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20732 10810 20760 11086
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20546 10364 20854 10373
rect 20546 10362 20552 10364
rect 20608 10362 20632 10364
rect 20688 10362 20712 10364
rect 20768 10362 20792 10364
rect 20848 10362 20854 10364
rect 20608 10310 20610 10362
rect 20790 10310 20792 10362
rect 20546 10308 20552 10310
rect 20608 10308 20632 10310
rect 20688 10308 20712 10310
rect 20768 10308 20792 10310
rect 20848 10308 20854 10310
rect 20546 10299 20854 10308
rect 21376 9654 21404 11018
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 21364 9648 21416 9654
rect 21364 9590 21416 9596
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 19904 9110 19932 9454
rect 21192 9382 21220 9454
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 19892 9104 19944 9110
rect 19892 9046 19944 9052
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 20088 7818 20116 8978
rect 20076 7812 20128 7818
rect 20076 7754 20128 7760
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19904 7546 19932 7686
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 19708 7200 19760 7206
rect 19708 7142 19760 7148
rect 19720 6662 19748 7142
rect 20272 6866 20300 7346
rect 20456 6866 20484 9318
rect 20546 9276 20854 9285
rect 20546 9274 20552 9276
rect 20608 9274 20632 9276
rect 20688 9274 20712 9276
rect 20768 9274 20792 9276
rect 20848 9274 20854 9276
rect 20608 9222 20610 9274
rect 20790 9222 20792 9274
rect 20546 9220 20552 9222
rect 20608 9220 20632 9222
rect 20688 9220 20712 9222
rect 20768 9220 20792 9222
rect 20848 9220 20854 9222
rect 20546 9211 20854 9220
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20916 8498 20944 8978
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20546 8188 20854 8197
rect 20546 8186 20552 8188
rect 20608 8186 20632 8188
rect 20688 8186 20712 8188
rect 20768 8186 20792 8188
rect 20848 8186 20854 8188
rect 20608 8134 20610 8186
rect 20790 8134 20792 8186
rect 20546 8132 20552 8134
rect 20608 8132 20632 8134
rect 20688 8132 20712 8134
rect 20768 8132 20792 8134
rect 20848 8132 20854 8134
rect 20546 8123 20854 8132
rect 20916 8090 20944 8230
rect 21008 8090 21036 8366
rect 21192 8362 21220 9318
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21192 7954 21220 8298
rect 21376 7954 21404 8434
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21468 7886 21496 8366
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21456 7336 21508 7342
rect 21456 7278 21508 7284
rect 20546 7100 20854 7109
rect 20546 7098 20552 7100
rect 20608 7098 20632 7100
rect 20688 7098 20712 7100
rect 20768 7098 20792 7100
rect 20848 7098 20854 7100
rect 20608 7046 20610 7098
rect 20790 7046 20792 7098
rect 20546 7044 20552 7046
rect 20608 7044 20632 7046
rect 20688 7044 20712 7046
rect 20768 7044 20792 7046
rect 20848 7044 20854 7046
rect 20546 7035 20854 7044
rect 20720 6928 20772 6934
rect 20640 6876 20720 6882
rect 20640 6870 20772 6876
rect 20260 6860 20312 6866
rect 20444 6860 20496 6866
rect 20260 6802 20312 6808
rect 20364 6820 20444 6848
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 19720 6390 19748 6598
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 20088 5846 20116 6598
rect 20076 5840 20128 5846
rect 20076 5782 20128 5788
rect 20272 5370 20300 6802
rect 20364 6118 20392 6820
rect 20444 6802 20496 6808
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 20640 6854 20760 6870
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 20364 5914 20392 6054
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20456 5828 20484 6598
rect 20548 6186 20576 6802
rect 20640 6254 20668 6854
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20732 6254 20760 6734
rect 21468 6458 21496 7278
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 21088 6180 21140 6186
rect 21088 6122 21140 6128
rect 20546 6012 20854 6021
rect 20546 6010 20552 6012
rect 20608 6010 20632 6012
rect 20688 6010 20712 6012
rect 20768 6010 20792 6012
rect 20848 6010 20854 6012
rect 20608 5958 20610 6010
rect 20790 5958 20792 6010
rect 20546 5956 20552 5958
rect 20608 5956 20632 5958
rect 20688 5956 20712 5958
rect 20768 5956 20792 5958
rect 20848 5956 20854 5958
rect 20546 5947 20854 5956
rect 20628 5840 20680 5846
rect 20456 5800 20628 5828
rect 20628 5782 20680 5788
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20640 5166 20668 5782
rect 21100 5642 21128 6122
rect 21456 6112 21508 6118
rect 21456 6054 21508 6060
rect 21088 5636 21140 5642
rect 21088 5578 21140 5584
rect 21468 5574 21496 6054
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21008 5166 21036 5510
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 20546 4924 20854 4933
rect 20546 4922 20552 4924
rect 20608 4922 20632 4924
rect 20688 4922 20712 4924
rect 20768 4922 20792 4924
rect 20848 4922 20854 4924
rect 20608 4870 20610 4922
rect 20790 4870 20792 4922
rect 20546 4868 20552 4870
rect 20608 4868 20632 4870
rect 20688 4868 20712 4870
rect 20768 4868 20792 4870
rect 20848 4868 20854 4870
rect 20546 4859 20854 4868
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19812 4486 19840 4762
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 19812 2774 19840 4422
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 20546 3836 20854 3845
rect 20546 3834 20552 3836
rect 20608 3834 20632 3836
rect 20688 3834 20712 3836
rect 20768 3834 20792 3836
rect 20848 3834 20854 3836
rect 20608 3782 20610 3834
rect 20790 3782 20792 3834
rect 20546 3780 20552 3782
rect 20608 3780 20632 3782
rect 20688 3780 20712 3782
rect 20768 3780 20792 3782
rect 20848 3780 20854 3782
rect 20546 3771 20854 3780
rect 21468 3602 21496 3878
rect 21456 3596 21508 3602
rect 21456 3538 21508 3544
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19892 3120 19944 3126
rect 19892 3062 19944 3068
rect 19720 2746 19840 2774
rect 19616 944 19668 950
rect 19616 886 19668 892
rect 19720 882 19748 2746
rect 19800 1896 19852 1902
rect 19800 1838 19852 1844
rect 19812 1426 19840 1838
rect 19904 1426 19932 3062
rect 19996 1902 20024 3334
rect 20546 2748 20854 2757
rect 20546 2746 20552 2748
rect 20608 2746 20632 2748
rect 20688 2746 20712 2748
rect 20768 2746 20792 2748
rect 20848 2746 20854 2748
rect 20608 2694 20610 2746
rect 20790 2694 20792 2746
rect 20546 2692 20552 2694
rect 20608 2692 20632 2694
rect 20688 2692 20712 2694
rect 20768 2692 20792 2694
rect 20848 2692 20854 2694
rect 20546 2683 20854 2692
rect 20258 2000 20314 2009
rect 20258 1935 20260 1944
rect 20312 1935 20314 1944
rect 20260 1906 20312 1912
rect 19984 1896 20036 1902
rect 19984 1838 20036 1844
rect 20352 1896 20404 1902
rect 20352 1838 20404 1844
rect 20364 1562 20392 1838
rect 20546 1660 20854 1669
rect 20546 1658 20552 1660
rect 20608 1658 20632 1660
rect 20688 1658 20712 1660
rect 20768 1658 20792 1660
rect 20848 1658 20854 1660
rect 20608 1606 20610 1658
rect 20790 1606 20792 1658
rect 20546 1604 20552 1606
rect 20608 1604 20632 1606
rect 20688 1604 20712 1606
rect 20768 1604 20792 1606
rect 20848 1604 20854 1606
rect 20546 1595 20854 1604
rect 20352 1556 20404 1562
rect 20352 1498 20404 1504
rect 20076 1488 20128 1494
rect 20076 1430 20128 1436
rect 19800 1420 19852 1426
rect 19800 1362 19852 1368
rect 19892 1420 19944 1426
rect 19892 1362 19944 1368
rect 19812 1290 19840 1362
rect 19800 1284 19852 1290
rect 19800 1226 19852 1232
rect 19708 876 19760 882
rect 19708 818 19760 824
rect 19812 814 19840 1226
rect 19800 808 19852 814
rect 19800 750 19852 756
rect 20088 400 20116 1430
rect 20364 814 20392 1498
rect 21468 1426 21496 3538
rect 21560 1766 21588 14742
rect 21652 13394 21680 14912
rect 21732 14894 21784 14900
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 22020 14074 22048 14418
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 22112 13870 22140 15302
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 22376 14884 22428 14890
rect 22376 14826 22428 14832
rect 22296 14618 22324 14826
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22388 14482 22416 14826
rect 22480 14822 22508 15574
rect 22756 15570 22784 15966
rect 22836 15904 22888 15910
rect 22836 15846 22888 15852
rect 22744 15564 22796 15570
rect 22744 15506 22796 15512
rect 22756 15162 22784 15506
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22744 14952 22796 14958
rect 22744 14894 22796 14900
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 22756 14414 22784 14894
rect 22848 14822 22876 15846
rect 23020 15564 23072 15570
rect 23020 15506 23072 15512
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22836 14816 22888 14822
rect 22836 14758 22888 14764
rect 22848 14550 22876 14758
rect 22836 14544 22888 14550
rect 22836 14486 22888 14492
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22940 14346 22968 15438
rect 22928 14340 22980 14346
rect 22928 14282 22980 14288
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 21732 13864 21784 13870
rect 21730 13832 21732 13841
rect 21824 13864 21876 13870
rect 21784 13832 21786 13841
rect 21824 13806 21876 13812
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 21730 13767 21786 13776
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21640 12708 21692 12714
rect 21640 12650 21692 12656
rect 21652 12617 21680 12650
rect 21638 12608 21694 12617
rect 21638 12543 21694 12552
rect 21744 12374 21772 13670
rect 21732 12368 21784 12374
rect 21732 12310 21784 12316
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 21744 10810 21772 11154
rect 21732 10804 21784 10810
rect 21732 10746 21784 10752
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21744 10130 21772 10406
rect 21836 10266 21864 13806
rect 22664 13802 22692 14214
rect 22940 14074 22968 14282
rect 22928 14068 22980 14074
rect 22928 14010 22980 14016
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22652 13796 22704 13802
rect 22652 13738 22704 13744
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22388 13462 22416 13670
rect 22376 13456 22428 13462
rect 22376 13398 22428 13404
rect 22756 12442 22784 13806
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 22848 12986 22876 13330
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22848 12220 22876 12922
rect 22940 12714 22968 14010
rect 22928 12708 22980 12714
rect 22928 12650 22980 12656
rect 22756 12192 22876 12220
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 22020 10169 22048 10474
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22006 10160 22062 10169
rect 21732 10124 21784 10130
rect 22006 10095 22008 10104
rect 21732 10066 21784 10072
rect 22060 10095 22062 10104
rect 22008 10066 22060 10072
rect 21640 9648 21692 9654
rect 21640 9590 21692 9596
rect 21652 8974 21680 9590
rect 22112 9518 22140 10202
rect 22204 10130 22232 10542
rect 22192 10124 22244 10130
rect 22192 10066 22244 10072
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 21652 8430 21680 8774
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 21744 8090 21772 9046
rect 22112 9042 22140 9454
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 21928 8430 21956 8774
rect 22204 8634 22232 9386
rect 22296 9382 22324 11154
rect 22756 11150 22784 12192
rect 22836 11688 22888 11694
rect 22836 11630 22888 11636
rect 22848 11218 22876 11630
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22652 11076 22704 11082
rect 22652 11018 22704 11024
rect 22664 10742 22692 11018
rect 22652 10736 22704 10742
rect 22652 10678 22704 10684
rect 22376 10192 22428 10198
rect 22376 10134 22428 10140
rect 22388 9722 22416 10134
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22296 8634 22324 9318
rect 22388 9178 22416 9658
rect 22756 9586 22784 11086
rect 22928 11008 22980 11014
rect 22928 10950 22980 10956
rect 22940 10606 22968 10950
rect 22928 10600 22980 10606
rect 22928 10542 22980 10548
rect 23032 10266 23060 15506
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22284 8628 22336 8634
rect 22284 8570 22336 8576
rect 21916 8424 21968 8430
rect 21916 8366 21968 8372
rect 22756 8362 22784 9318
rect 23124 8922 23152 16934
rect 24136 16794 24164 17002
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 24136 16658 24164 16730
rect 24124 16652 24176 16658
rect 24124 16594 24176 16600
rect 24308 16652 24360 16658
rect 24308 16594 24360 16600
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23492 16182 23520 16526
rect 23904 16348 24212 16357
rect 23904 16346 23910 16348
rect 23966 16346 23990 16348
rect 24046 16346 24070 16348
rect 24126 16346 24150 16348
rect 24206 16346 24212 16348
rect 23966 16294 23968 16346
rect 24148 16294 24150 16346
rect 23904 16292 23910 16294
rect 23966 16292 23990 16294
rect 24046 16292 24070 16294
rect 24126 16292 24150 16294
rect 24206 16292 24212 16294
rect 23904 16283 24212 16292
rect 23480 16176 23532 16182
rect 23480 16118 23532 16124
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23308 15706 23336 15846
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23204 14952 23256 14958
rect 23204 14894 23256 14900
rect 23216 13938 23244 14894
rect 23308 14822 23336 15642
rect 23492 15638 23520 16118
rect 23480 15632 23532 15638
rect 23480 15574 23532 15580
rect 23572 15428 23624 15434
rect 23572 15370 23624 15376
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23492 14890 23520 15302
rect 23480 14884 23532 14890
rect 23480 14826 23532 14832
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23584 14482 23612 15370
rect 23904 15260 24212 15269
rect 23904 15258 23910 15260
rect 23966 15258 23990 15260
rect 24046 15258 24070 15260
rect 24126 15258 24150 15260
rect 24206 15258 24212 15260
rect 23966 15206 23968 15258
rect 24148 15206 24150 15258
rect 23904 15204 23910 15206
rect 23966 15204 23990 15206
rect 24046 15204 24070 15206
rect 24126 15204 24150 15206
rect 24206 15204 24212 15206
rect 23904 15195 24212 15204
rect 23848 15020 23900 15026
rect 23848 14962 23900 14968
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23204 13932 23256 13938
rect 23204 13874 23256 13880
rect 23204 13728 23256 13734
rect 23204 13670 23256 13676
rect 23216 12782 23244 13670
rect 23204 12776 23256 12782
rect 23204 12718 23256 12724
rect 23308 10266 23336 14418
rect 23584 13841 23612 14418
rect 23860 14414 23888 14962
rect 23848 14408 23900 14414
rect 23848 14350 23900 14356
rect 23904 14172 24212 14181
rect 23904 14170 23910 14172
rect 23966 14170 23990 14172
rect 24046 14170 24070 14172
rect 24126 14170 24150 14172
rect 24206 14170 24212 14172
rect 23966 14118 23968 14170
rect 24148 14118 24150 14170
rect 23904 14116 23910 14118
rect 23966 14116 23990 14118
rect 24046 14116 24070 14118
rect 24126 14116 24150 14118
rect 24206 14116 24212 14118
rect 23904 14107 24212 14116
rect 24320 14074 24348 16594
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24492 15156 24544 15162
rect 24492 15098 24544 15104
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24412 14278 24440 14758
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24412 13870 24440 14214
rect 24504 13938 24532 15098
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 24216 13864 24268 13870
rect 23570 13832 23626 13841
rect 24400 13864 24452 13870
rect 24268 13841 24348 13852
rect 24268 13832 24362 13841
rect 24268 13824 24306 13832
rect 24216 13806 24268 13812
rect 23570 13767 23626 13776
rect 24400 13806 24452 13812
rect 24306 13767 24362 13776
rect 23480 13184 23532 13190
rect 23480 13126 23532 13132
rect 23492 12850 23520 13126
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23388 12708 23440 12714
rect 23388 12650 23440 12656
rect 23400 12374 23428 12650
rect 23388 12368 23440 12374
rect 23388 12310 23440 12316
rect 23492 12306 23520 12786
rect 23584 12646 23612 13767
rect 23904 13084 24212 13093
rect 23904 13082 23910 13084
rect 23966 13082 23990 13084
rect 24046 13082 24070 13084
rect 24126 13082 24150 13084
rect 24206 13082 24212 13084
rect 23966 13030 23968 13082
rect 24148 13030 24150 13082
rect 23904 13028 23910 13030
rect 23966 13028 23990 13030
rect 24046 13028 24070 13030
rect 24126 13028 24150 13030
rect 24206 13028 24212 13030
rect 23904 13019 24212 13028
rect 24320 12782 24348 13767
rect 24412 12918 24440 13806
rect 24400 12912 24452 12918
rect 24400 12854 24452 12860
rect 24308 12776 24360 12782
rect 24308 12718 24360 12724
rect 23572 12640 23624 12646
rect 23572 12582 23624 12588
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24320 12306 24348 12582
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 24308 12300 24360 12306
rect 24308 12242 24360 12248
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 23492 11898 23520 12106
rect 23904 11996 24212 12005
rect 23904 11994 23910 11996
rect 23966 11994 23990 11996
rect 24046 11994 24070 11996
rect 24126 11994 24150 11996
rect 24206 11994 24212 11996
rect 23966 11942 23968 11994
rect 24148 11942 24150 11994
rect 23904 11940 23910 11942
rect 23966 11940 23990 11942
rect 24046 11940 24070 11942
rect 24126 11940 24150 11942
rect 24206 11940 24212 11942
rect 23904 11931 24212 11940
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23386 10160 23442 10169
rect 23296 10124 23348 10130
rect 23386 10095 23388 10104
rect 23296 10066 23348 10072
rect 23440 10095 23442 10104
rect 23388 10066 23440 10072
rect 23308 9602 23336 10066
rect 23308 9574 23428 9602
rect 23400 9518 23428 9574
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23296 9444 23348 9450
rect 23296 9386 23348 9392
rect 23308 9042 23336 9386
rect 23400 9042 23428 9454
rect 23584 9058 23612 10746
rect 23676 10606 23704 11494
rect 23756 11212 23808 11218
rect 23756 11154 23808 11160
rect 23768 10810 23796 11154
rect 23904 10908 24212 10917
rect 23904 10906 23910 10908
rect 23966 10906 23990 10908
rect 24046 10906 24070 10908
rect 24126 10906 24150 10908
rect 24206 10906 24212 10908
rect 23966 10854 23968 10906
rect 24148 10854 24150 10906
rect 23904 10852 23910 10854
rect 23966 10852 23990 10854
rect 24046 10852 24070 10854
rect 24126 10852 24150 10854
rect 24206 10852 24212 10854
rect 23904 10843 24212 10852
rect 23756 10804 23808 10810
rect 23756 10746 23808 10752
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 24124 10464 24176 10470
rect 24320 10452 24348 12242
rect 24412 11762 24440 12582
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24412 11354 24440 11698
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24176 10424 24348 10452
rect 24124 10406 24176 10412
rect 24136 10198 24164 10406
rect 24124 10192 24176 10198
rect 24124 10134 24176 10140
rect 23756 10124 23808 10130
rect 23756 10066 23808 10072
rect 24308 10124 24360 10130
rect 24308 10066 24360 10072
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 23768 9518 23796 10066
rect 24320 9926 24348 10066
rect 24412 10033 24440 10066
rect 24398 10024 24454 10033
rect 24504 9994 24532 10542
rect 24398 9959 24454 9968
rect 24492 9988 24544 9994
rect 24492 9930 24544 9936
rect 24308 9920 24360 9926
rect 24308 9862 24360 9868
rect 23904 9820 24212 9829
rect 23904 9818 23910 9820
rect 23966 9818 23990 9820
rect 24046 9818 24070 9820
rect 24126 9818 24150 9820
rect 24206 9818 24212 9820
rect 23966 9766 23968 9818
rect 24148 9766 24150 9818
rect 23904 9764 23910 9766
rect 23966 9764 23990 9766
rect 24046 9764 24070 9766
rect 24126 9764 24150 9766
rect 24206 9764 24212 9766
rect 23904 9755 24212 9764
rect 24504 9518 24532 9930
rect 23756 9512 23808 9518
rect 23756 9454 23808 9460
rect 24492 9512 24544 9518
rect 24492 9454 24544 9460
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 23296 9036 23348 9042
rect 23296 8978 23348 8984
rect 23388 9036 23440 9042
rect 23584 9030 23704 9058
rect 23388 8978 23440 8984
rect 22940 8894 23152 8922
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 22744 8356 22796 8362
rect 22744 8298 22796 8304
rect 22836 8356 22888 8362
rect 22836 8298 22888 8304
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 21836 8090 21864 8230
rect 21732 8084 21784 8090
rect 21732 8026 21784 8032
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21836 7954 21864 8026
rect 22376 8016 22428 8022
rect 22652 8016 22704 8022
rect 22428 7976 22652 8004
rect 22376 7958 22428 7964
rect 22652 7958 22704 7964
rect 22848 7954 22876 8298
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 22836 7948 22888 7954
rect 22836 7890 22888 7896
rect 22284 7812 22336 7818
rect 22284 7754 22336 7760
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 21730 7440 21786 7449
rect 21730 7375 21786 7384
rect 21744 7342 21772 7375
rect 21732 7336 21784 7342
rect 21732 7278 21784 7284
rect 21744 6934 21772 7278
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22112 6934 22140 7142
rect 21732 6928 21784 6934
rect 21732 6870 21784 6876
rect 22100 6928 22152 6934
rect 22100 6870 22152 6876
rect 22204 6458 22232 7686
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22296 6186 22324 7754
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22388 6186 22416 7686
rect 22284 6180 22336 6186
rect 22284 6122 22336 6128
rect 22376 6180 22428 6186
rect 22376 6122 22428 6128
rect 22388 5914 22416 6122
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22112 4282 22140 5850
rect 22572 5778 22600 6054
rect 22376 5772 22428 5778
rect 22376 5714 22428 5720
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22388 5166 22416 5714
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 22480 4758 22508 5306
rect 22664 5234 22692 5714
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22468 4752 22520 4758
rect 22468 4694 22520 4700
rect 22664 4690 22692 5170
rect 22652 4684 22704 4690
rect 22652 4626 22704 4632
rect 22836 4684 22888 4690
rect 22836 4626 22888 4632
rect 22848 4282 22876 4626
rect 22100 4276 22152 4282
rect 22100 4218 22152 4224
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 21732 1896 21784 1902
rect 21732 1838 21784 1844
rect 21548 1760 21600 1766
rect 21548 1702 21600 1708
rect 21560 1562 21588 1702
rect 21548 1556 21600 1562
rect 21548 1498 21600 1504
rect 21744 1426 21772 1838
rect 21824 1556 21876 1562
rect 21824 1498 21876 1504
rect 21456 1420 21508 1426
rect 21456 1362 21508 1368
rect 21732 1420 21784 1426
rect 21732 1362 21784 1368
rect 20352 808 20404 814
rect 20352 750 20404 756
rect 20546 572 20854 581
rect 20546 570 20552 572
rect 20608 570 20632 572
rect 20688 570 20712 572
rect 20768 570 20792 572
rect 20848 570 20854 572
rect 20608 518 20610 570
rect 20790 518 20792 570
rect 20546 516 20552 518
rect 20608 516 20632 518
rect 20688 516 20712 518
rect 20768 516 20792 518
rect 20848 516 20854 518
rect 20546 507 20854 516
rect 21836 400 21864 1498
rect 22006 1456 22062 1465
rect 22940 1426 22968 8894
rect 23112 8832 23164 8838
rect 23112 8774 23164 8780
rect 23124 8566 23152 8774
rect 23112 8560 23164 8566
rect 23112 8502 23164 8508
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23032 7954 23060 8230
rect 23216 7954 23244 8910
rect 23308 8906 23336 8978
rect 23296 8900 23348 8906
rect 23296 8842 23348 8848
rect 23400 8650 23428 8978
rect 23572 8900 23624 8906
rect 23572 8842 23624 8848
rect 23308 8622 23428 8650
rect 23308 8362 23336 8622
rect 23584 8566 23612 8842
rect 23572 8560 23624 8566
rect 23572 8502 23624 8508
rect 23296 8356 23348 8362
rect 23296 8298 23348 8304
rect 23308 7954 23336 8298
rect 23584 7970 23612 8502
rect 23492 7954 23612 7970
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 23480 7948 23612 7954
rect 23532 7942 23612 7948
rect 23480 7890 23532 7896
rect 23032 7546 23060 7890
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 23216 7002 23244 7890
rect 23492 7546 23520 7890
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23388 7268 23440 7274
rect 23388 7210 23440 7216
rect 23204 6996 23256 7002
rect 23204 6938 23256 6944
rect 23020 6860 23072 6866
rect 23020 6802 23072 6808
rect 23032 6390 23060 6802
rect 23400 6730 23428 7210
rect 23388 6724 23440 6730
rect 23388 6666 23440 6672
rect 23400 6390 23428 6666
rect 23020 6384 23072 6390
rect 23020 6326 23072 6332
rect 23388 6384 23440 6390
rect 23388 6326 23440 6332
rect 23032 5166 23060 6326
rect 23296 5908 23348 5914
rect 23296 5850 23348 5856
rect 23020 5160 23072 5166
rect 23020 5102 23072 5108
rect 23308 5098 23336 5850
rect 23400 5846 23428 6326
rect 23584 6322 23612 7822
rect 23676 6934 23704 9030
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 24308 9036 24360 9042
rect 24308 8978 24360 8984
rect 23768 8634 23796 8978
rect 23904 8732 24212 8741
rect 23904 8730 23910 8732
rect 23966 8730 23990 8732
rect 24046 8730 24070 8732
rect 24126 8730 24150 8732
rect 24206 8730 24212 8732
rect 23966 8678 23968 8730
rect 24148 8678 24150 8730
rect 23904 8676 23910 8678
rect 23966 8676 23990 8678
rect 24046 8676 24070 8678
rect 24126 8676 24150 8678
rect 24206 8676 24212 8678
rect 23904 8667 24212 8676
rect 24320 8634 24348 8978
rect 24400 8832 24452 8838
rect 24400 8774 24452 8780
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 24308 8628 24360 8634
rect 24308 8570 24360 8576
rect 24412 8498 24440 8774
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 24400 8492 24452 8498
rect 24400 8434 24452 8440
rect 23756 8016 23808 8022
rect 23756 7958 23808 7964
rect 23768 7274 23796 7958
rect 23860 7886 23888 8434
rect 24124 8424 24176 8430
rect 24124 8366 24176 8372
rect 24136 7954 24164 8366
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23904 7644 24212 7653
rect 23904 7642 23910 7644
rect 23966 7642 23990 7644
rect 24046 7642 24070 7644
rect 24126 7642 24150 7644
rect 24206 7642 24212 7644
rect 23966 7590 23968 7642
rect 24148 7590 24150 7642
rect 23904 7588 23910 7590
rect 23966 7588 23990 7590
rect 24046 7588 24070 7590
rect 24126 7588 24150 7590
rect 24206 7588 24212 7590
rect 23904 7579 24212 7588
rect 23756 7268 23808 7274
rect 23756 7210 23808 7216
rect 23768 7002 23796 7210
rect 23756 6996 23808 7002
rect 23756 6938 23808 6944
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 23664 6928 23716 6934
rect 23664 6870 23716 6876
rect 23904 6556 24212 6565
rect 23904 6554 23910 6556
rect 23966 6554 23990 6556
rect 24046 6554 24070 6556
rect 24126 6554 24150 6556
rect 24206 6554 24212 6556
rect 23966 6502 23968 6554
rect 24148 6502 24150 6554
rect 23904 6500 23910 6502
rect 23966 6500 23990 6502
rect 24046 6500 24070 6502
rect 24126 6500 24150 6502
rect 24206 6500 24212 6502
rect 23904 6491 24212 6500
rect 24412 6322 24440 6938
rect 24504 6866 24532 9318
rect 24596 7834 24624 15982
rect 24688 14890 24716 17002
rect 25320 16652 25372 16658
rect 25320 16594 25372 16600
rect 24952 16448 25004 16454
rect 24952 16390 25004 16396
rect 24964 15978 24992 16390
rect 25332 16250 25360 16594
rect 25320 16244 25372 16250
rect 25320 16186 25372 16192
rect 24860 15972 24912 15978
rect 24860 15914 24912 15920
rect 24952 15972 25004 15978
rect 24952 15914 25004 15920
rect 24872 15502 24900 15914
rect 24768 15496 24820 15502
rect 24768 15438 24820 15444
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 24780 15162 24808 15438
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 24688 12782 24716 14826
rect 24872 14414 24900 15438
rect 25044 14884 25096 14890
rect 25044 14826 25096 14832
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24872 12918 24900 14350
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 24964 13530 24992 13806
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 24860 12912 24912 12918
rect 24860 12854 24912 12860
rect 24676 12776 24728 12782
rect 24676 12718 24728 12724
rect 24688 12102 24716 12718
rect 24768 12164 24820 12170
rect 24768 12106 24820 12112
rect 24676 12096 24728 12102
rect 24676 12038 24728 12044
rect 24688 11898 24716 12038
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24676 10532 24728 10538
rect 24676 10474 24728 10480
rect 24688 9994 24716 10474
rect 24676 9988 24728 9994
rect 24676 9930 24728 9936
rect 24780 9654 24808 12106
rect 24872 11762 24900 12854
rect 25056 12850 25084 14826
rect 25412 13728 25464 13734
rect 25412 13670 25464 13676
rect 25228 13320 25280 13326
rect 25228 13262 25280 13268
rect 25240 12986 25268 13262
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25044 12844 25096 12850
rect 25044 12786 25096 12792
rect 25056 12646 25084 12786
rect 25424 12782 25452 13670
rect 25412 12776 25464 12782
rect 25412 12718 25464 12724
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 25056 12442 25084 12582
rect 25044 12436 25096 12442
rect 25044 12378 25096 12384
rect 25516 12345 25544 17070
rect 25964 16788 26016 16794
rect 25964 16730 26016 16736
rect 25596 16720 25648 16726
rect 25596 16662 25648 16668
rect 25608 15638 25636 16662
rect 25688 16448 25740 16454
rect 25688 16390 25740 16396
rect 25700 16182 25728 16390
rect 25688 16176 25740 16182
rect 25688 16118 25740 16124
rect 25596 15632 25648 15638
rect 25596 15574 25648 15580
rect 25596 12708 25648 12714
rect 25596 12650 25648 12656
rect 25608 12442 25636 12650
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25502 12336 25558 12345
rect 25044 12300 25096 12306
rect 25502 12271 25558 12280
rect 25044 12242 25096 12248
rect 24860 11756 24912 11762
rect 24860 11698 24912 11704
rect 24872 11218 24900 11698
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24872 10674 24900 11154
rect 25056 10742 25084 12242
rect 25412 12096 25464 12102
rect 25412 12038 25464 12044
rect 25424 11694 25452 12038
rect 25412 11688 25464 11694
rect 25412 11630 25464 11636
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 25044 10736 25096 10742
rect 25044 10678 25096 10684
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24872 9654 24900 9998
rect 24964 9994 24992 10542
rect 25056 10130 25084 10678
rect 25148 10130 25176 11494
rect 25320 10464 25372 10470
rect 25320 10406 25372 10412
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 25136 10124 25188 10130
rect 25136 10066 25188 10072
rect 25228 10124 25280 10130
rect 25228 10066 25280 10072
rect 24952 9988 25004 9994
rect 24952 9930 25004 9936
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 24964 9586 24992 9930
rect 25056 9926 25084 10066
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 25240 9518 25268 10066
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 24952 9376 25004 9382
rect 24952 9318 25004 9324
rect 24964 8498 24992 9318
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 24964 8090 24992 8434
rect 24952 8084 25004 8090
rect 24952 8026 25004 8032
rect 25332 7834 25360 10406
rect 25700 8974 25728 16118
rect 25976 14958 26004 16730
rect 26252 16658 26280 17734
rect 26514 17600 26570 17734
rect 27158 17600 27214 18000
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 26240 16040 26292 16046
rect 26240 15982 26292 15988
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 25964 14952 26016 14958
rect 25964 14894 26016 14900
rect 25884 14074 25912 14894
rect 26252 14618 26280 15982
rect 26344 15366 26372 17070
rect 26976 17060 27028 17066
rect 26976 17002 27028 17008
rect 26700 16992 26752 16998
rect 26700 16934 26752 16940
rect 26712 16658 26740 16934
rect 26988 16658 27016 17002
rect 26700 16652 26752 16658
rect 26700 16594 26752 16600
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 26976 16652 27028 16658
rect 26976 16594 27028 16600
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26620 15570 26648 15846
rect 26896 15706 26924 16594
rect 26884 15700 26936 15706
rect 26884 15642 26936 15648
rect 26424 15564 26476 15570
rect 26424 15506 26476 15512
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26700 15564 26752 15570
rect 26700 15506 26752 15512
rect 26792 15564 26844 15570
rect 26792 15506 26844 15512
rect 26884 15564 26936 15570
rect 26884 15506 26936 15512
rect 26332 15360 26384 15366
rect 26332 15302 26384 15308
rect 26240 14612 26292 14618
rect 26240 14554 26292 14560
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 26344 14006 26372 15302
rect 26436 14906 26464 15506
rect 26620 14958 26648 15506
rect 26608 14952 26660 14958
rect 26436 14878 26556 14906
rect 26608 14894 26660 14900
rect 26424 14816 26476 14822
rect 26424 14758 26476 14764
rect 26436 14550 26464 14758
rect 26424 14544 26476 14550
rect 26424 14486 26476 14492
rect 26424 14408 26476 14414
rect 26424 14350 26476 14356
rect 26332 14000 26384 14006
rect 26332 13942 26384 13948
rect 25964 13864 26016 13870
rect 26056 13864 26108 13870
rect 25964 13806 26016 13812
rect 26054 13832 26056 13841
rect 26108 13832 26110 13841
rect 26238 13832 26294 13841
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25792 12306 25820 13126
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 25884 12306 25912 12582
rect 25976 12442 26004 13806
rect 26054 13767 26110 13776
rect 26160 13790 26238 13818
rect 25964 12436 26016 12442
rect 25964 12378 26016 12384
rect 26160 12345 26188 13790
rect 26238 13767 26294 13776
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26252 12374 26280 13670
rect 26240 12368 26292 12374
rect 26146 12336 26202 12345
rect 25780 12300 25832 12306
rect 25780 12242 25832 12248
rect 25872 12300 25924 12306
rect 26240 12310 26292 12316
rect 26146 12271 26202 12280
rect 25872 12242 25924 12248
rect 26240 12232 26292 12238
rect 26240 12174 26292 12180
rect 26252 11898 26280 12174
rect 26240 11892 26292 11898
rect 26240 11834 26292 11840
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 26252 11354 26280 11630
rect 26240 11348 26292 11354
rect 26240 11290 26292 11296
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 25884 10266 25912 11086
rect 26436 10810 26464 14350
rect 26528 14006 26556 14878
rect 26712 14498 26740 15506
rect 26804 14618 26832 15506
rect 26792 14612 26844 14618
rect 26792 14554 26844 14560
rect 26620 14470 26740 14498
rect 26620 14278 26648 14470
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26516 14000 26568 14006
rect 26516 13942 26568 13948
rect 26620 13870 26648 14214
rect 26790 13968 26846 13977
rect 26896 13954 26924 15506
rect 26846 13926 26924 13954
rect 26790 13903 26846 13912
rect 26804 13870 26832 13903
rect 26516 13864 26568 13870
rect 26516 13806 26568 13812
rect 26608 13864 26660 13870
rect 26608 13806 26660 13812
rect 26700 13864 26752 13870
rect 26700 13806 26752 13812
rect 26792 13864 26844 13870
rect 27172 13841 27200 17600
rect 27262 16892 27570 16901
rect 27262 16890 27268 16892
rect 27324 16890 27348 16892
rect 27404 16890 27428 16892
rect 27484 16890 27508 16892
rect 27564 16890 27570 16892
rect 27324 16838 27326 16890
rect 27506 16838 27508 16890
rect 27262 16836 27268 16838
rect 27324 16836 27348 16838
rect 27404 16836 27428 16838
rect 27484 16836 27508 16838
rect 27564 16836 27570 16838
rect 27262 16827 27570 16836
rect 27262 15804 27570 15813
rect 27262 15802 27268 15804
rect 27324 15802 27348 15804
rect 27404 15802 27428 15804
rect 27484 15802 27508 15804
rect 27564 15802 27570 15804
rect 27324 15750 27326 15802
rect 27506 15750 27508 15802
rect 27262 15748 27268 15750
rect 27324 15748 27348 15750
rect 27404 15748 27428 15750
rect 27484 15748 27508 15750
rect 27564 15748 27570 15750
rect 27262 15739 27570 15748
rect 27262 14716 27570 14725
rect 27262 14714 27268 14716
rect 27324 14714 27348 14716
rect 27404 14714 27428 14716
rect 27484 14714 27508 14716
rect 27564 14714 27570 14716
rect 27324 14662 27326 14714
rect 27506 14662 27508 14714
rect 27262 14660 27268 14662
rect 27324 14660 27348 14662
rect 27404 14660 27428 14662
rect 27484 14660 27508 14662
rect 27564 14660 27570 14662
rect 27262 14651 27570 14660
rect 26792 13806 26844 13812
rect 27158 13832 27214 13841
rect 26528 13394 26556 13806
rect 26516 13388 26568 13394
rect 26516 13330 26568 13336
rect 26528 12986 26556 13330
rect 26516 12980 26568 12986
rect 26516 12922 26568 12928
rect 26712 11694 26740 13806
rect 27158 13767 27214 13776
rect 27262 13628 27570 13637
rect 27262 13626 27268 13628
rect 27324 13626 27348 13628
rect 27404 13626 27428 13628
rect 27484 13626 27508 13628
rect 27564 13626 27570 13628
rect 27324 13574 27326 13626
rect 27506 13574 27508 13626
rect 27262 13572 27268 13574
rect 27324 13572 27348 13574
rect 27404 13572 27428 13574
rect 27484 13572 27508 13574
rect 27564 13572 27570 13574
rect 27262 13563 27570 13572
rect 27262 12540 27570 12549
rect 27262 12538 27268 12540
rect 27324 12538 27348 12540
rect 27404 12538 27428 12540
rect 27484 12538 27508 12540
rect 27564 12538 27570 12540
rect 27324 12486 27326 12538
rect 27506 12486 27508 12538
rect 27262 12484 27268 12486
rect 27324 12484 27348 12486
rect 27404 12484 27428 12486
rect 27484 12484 27508 12486
rect 27564 12484 27570 12486
rect 27262 12475 27570 12484
rect 26700 11688 26752 11694
rect 26700 11630 26752 11636
rect 27262 11452 27570 11461
rect 27262 11450 27268 11452
rect 27324 11450 27348 11452
rect 27404 11450 27428 11452
rect 27484 11450 27508 11452
rect 27564 11450 27570 11452
rect 27324 11398 27326 11450
rect 27506 11398 27508 11450
rect 27262 11396 27268 11398
rect 27324 11396 27348 11398
rect 27404 11396 27428 11398
rect 27484 11396 27508 11398
rect 27564 11396 27570 11398
rect 27262 11387 27570 11396
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 26436 10130 26464 10746
rect 27262 10364 27570 10373
rect 27262 10362 27268 10364
rect 27324 10362 27348 10364
rect 27404 10362 27428 10364
rect 27484 10362 27508 10364
rect 27564 10362 27570 10364
rect 27324 10310 27326 10362
rect 27506 10310 27508 10362
rect 27262 10308 27268 10310
rect 27324 10308 27348 10310
rect 27404 10308 27428 10310
rect 27484 10308 27508 10310
rect 27564 10308 27570 10310
rect 27262 10299 27570 10308
rect 25872 10124 25924 10130
rect 25872 10066 25924 10072
rect 26424 10124 26476 10130
rect 26424 10066 26476 10072
rect 25780 9036 25832 9042
rect 25780 8978 25832 8984
rect 25412 8968 25464 8974
rect 25412 8910 25464 8916
rect 25688 8968 25740 8974
rect 25688 8910 25740 8916
rect 25424 8634 25452 8910
rect 25596 8900 25648 8906
rect 25596 8842 25648 8848
rect 25504 8832 25556 8838
rect 25504 8774 25556 8780
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25424 8022 25452 8570
rect 25516 8362 25544 8774
rect 25504 8356 25556 8362
rect 25504 8298 25556 8304
rect 25412 8016 25464 8022
rect 25412 7958 25464 7964
rect 24596 7806 24716 7834
rect 24584 7744 24636 7750
rect 24584 7686 24636 7692
rect 24596 7342 24624 7686
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 24688 6882 24716 7806
rect 25240 7806 25360 7834
rect 25240 6934 25268 7806
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25332 7342 25360 7686
rect 25320 7336 25372 7342
rect 25320 7278 25372 7284
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24596 6854 24716 6882
rect 25228 6928 25280 6934
rect 25228 6870 25280 6876
rect 24768 6860 24820 6866
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 24400 6316 24452 6322
rect 24400 6258 24452 6264
rect 24412 5914 24440 6258
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 23388 5840 23440 5846
rect 23388 5782 23440 5788
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23296 5092 23348 5098
rect 23296 5034 23348 5040
rect 23400 5030 23428 5170
rect 23676 5166 23704 5850
rect 24504 5778 24532 6802
rect 24492 5772 24544 5778
rect 24492 5714 24544 5720
rect 24596 5658 24624 6854
rect 24768 6802 24820 6808
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24688 6458 24716 6734
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24780 6186 24808 6802
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 24952 6656 25004 6662
rect 24952 6598 25004 6604
rect 24964 6458 24992 6598
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 24504 5630 24624 5658
rect 24308 5568 24360 5574
rect 24308 5510 24360 5516
rect 23904 5468 24212 5477
rect 23904 5466 23910 5468
rect 23966 5466 23990 5468
rect 24046 5466 24070 5468
rect 24126 5466 24150 5468
rect 24206 5466 24212 5468
rect 23966 5414 23968 5466
rect 24148 5414 24150 5466
rect 23904 5412 23910 5414
rect 23966 5412 23990 5414
rect 24046 5412 24070 5414
rect 24126 5412 24150 5414
rect 24206 5412 24212 5414
rect 23904 5403 24212 5412
rect 24320 5166 24348 5510
rect 24504 5166 24532 5630
rect 24964 5370 24992 6394
rect 25148 5914 25176 6734
rect 25136 5908 25188 5914
rect 25136 5850 25188 5856
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 25240 5234 25268 6870
rect 25424 6458 25452 7958
rect 25504 7948 25556 7954
rect 25504 7890 25556 7896
rect 25516 7546 25544 7890
rect 25504 7540 25556 7546
rect 25504 7482 25556 7488
rect 25608 6866 25636 8842
rect 25700 8294 25728 8910
rect 25688 8288 25740 8294
rect 25688 8230 25740 8236
rect 25792 7478 25820 8978
rect 25780 7472 25832 7478
rect 25780 7414 25832 7420
rect 25780 7336 25832 7342
rect 25780 7278 25832 7284
rect 25688 7200 25740 7206
rect 25688 7142 25740 7148
rect 25596 6860 25648 6866
rect 25596 6802 25648 6808
rect 25412 6452 25464 6458
rect 25412 6394 25464 6400
rect 25424 5846 25452 6394
rect 25700 6254 25728 7142
rect 25792 7002 25820 7278
rect 25780 6996 25832 7002
rect 25780 6938 25832 6944
rect 25884 6798 25912 10066
rect 26422 10024 26478 10033
rect 26422 9959 26424 9968
rect 26476 9959 26478 9968
rect 26424 9930 26476 9936
rect 27262 9276 27570 9285
rect 27262 9274 27268 9276
rect 27324 9274 27348 9276
rect 27404 9274 27428 9276
rect 27484 9274 27508 9276
rect 27564 9274 27570 9276
rect 27324 9222 27326 9274
rect 27506 9222 27508 9274
rect 27262 9220 27268 9222
rect 27324 9220 27348 9222
rect 27404 9220 27428 9222
rect 27484 9220 27508 9222
rect 27564 9220 27570 9222
rect 27262 9211 27570 9220
rect 26424 9104 26476 9110
rect 26424 9046 26476 9052
rect 26436 8090 26464 9046
rect 26516 8288 26568 8294
rect 26516 8230 26568 8236
rect 26424 8084 26476 8090
rect 26424 8026 26476 8032
rect 26528 7954 26556 8230
rect 27262 8188 27570 8197
rect 27262 8186 27268 8188
rect 27324 8186 27348 8188
rect 27404 8186 27428 8188
rect 27484 8186 27508 8188
rect 27564 8186 27570 8188
rect 27324 8134 27326 8186
rect 27506 8134 27508 8186
rect 27262 8132 27268 8134
rect 27324 8132 27348 8134
rect 27404 8132 27428 8134
rect 27484 8132 27508 8134
rect 27564 8132 27570 8134
rect 27262 8123 27570 8132
rect 26516 7948 26568 7954
rect 26516 7890 26568 7896
rect 27262 7100 27570 7109
rect 27262 7098 27268 7100
rect 27324 7098 27348 7100
rect 27404 7098 27428 7100
rect 27484 7098 27508 7100
rect 27564 7098 27570 7100
rect 27324 7046 27326 7098
rect 27506 7046 27508 7098
rect 27262 7044 27268 7046
rect 27324 7044 27348 7046
rect 27404 7044 27428 7046
rect 27484 7044 27508 7046
rect 27564 7044 27570 7046
rect 27262 7035 27570 7044
rect 25872 6792 25924 6798
rect 25872 6734 25924 6740
rect 25884 6458 25912 6734
rect 25872 6452 25924 6458
rect 25872 6394 25924 6400
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 27262 6012 27570 6021
rect 27262 6010 27268 6012
rect 27324 6010 27348 6012
rect 27404 6010 27428 6012
rect 27484 6010 27508 6012
rect 27564 6010 27570 6012
rect 27324 5958 27326 6010
rect 27506 5958 27508 6010
rect 27262 5956 27268 5958
rect 27324 5956 27348 5958
rect 27404 5956 27428 5958
rect 27484 5956 27508 5958
rect 27564 5956 27570 5958
rect 27262 5947 27570 5956
rect 25412 5840 25464 5846
rect 25412 5782 25464 5788
rect 25688 5772 25740 5778
rect 25688 5714 25740 5720
rect 25700 5370 25728 5714
rect 25688 5364 25740 5370
rect 25688 5306 25740 5312
rect 25228 5228 25280 5234
rect 25228 5170 25280 5176
rect 23664 5160 23716 5166
rect 23664 5102 23716 5108
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 24308 5160 24360 5166
rect 24308 5102 24360 5108
rect 24492 5160 24544 5166
rect 24492 5102 24544 5108
rect 23388 5024 23440 5030
rect 23388 4966 23440 4972
rect 23664 5024 23716 5030
rect 23664 4966 23716 4972
rect 23676 4078 23704 4966
rect 24044 4826 24072 5102
rect 24032 4820 24084 4826
rect 24032 4762 24084 4768
rect 24504 4758 24532 5102
rect 27262 4924 27570 4933
rect 27262 4922 27268 4924
rect 27324 4922 27348 4924
rect 27404 4922 27428 4924
rect 27484 4922 27508 4924
rect 27564 4922 27570 4924
rect 27324 4870 27326 4922
rect 27506 4870 27508 4922
rect 27262 4868 27268 4870
rect 27324 4868 27348 4870
rect 27404 4868 27428 4870
rect 27484 4868 27508 4870
rect 27564 4868 27570 4870
rect 27262 4859 27570 4868
rect 24492 4752 24544 4758
rect 24492 4694 24544 4700
rect 23904 4380 24212 4389
rect 23904 4378 23910 4380
rect 23966 4378 23990 4380
rect 24046 4378 24070 4380
rect 24126 4378 24150 4380
rect 24206 4378 24212 4380
rect 23966 4326 23968 4378
rect 24148 4326 24150 4378
rect 23904 4324 23910 4326
rect 23966 4324 23990 4326
rect 24046 4324 24070 4326
rect 24126 4324 24150 4326
rect 24206 4324 24212 4326
rect 23904 4315 24212 4324
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 27262 3836 27570 3845
rect 27262 3834 27268 3836
rect 27324 3834 27348 3836
rect 27404 3834 27428 3836
rect 27484 3834 27508 3836
rect 27564 3834 27570 3836
rect 27324 3782 27326 3834
rect 27506 3782 27508 3834
rect 27262 3780 27268 3782
rect 27324 3780 27348 3782
rect 27404 3780 27428 3782
rect 27484 3780 27508 3782
rect 27564 3780 27570 3782
rect 27262 3771 27570 3780
rect 23904 3292 24212 3301
rect 23904 3290 23910 3292
rect 23966 3290 23990 3292
rect 24046 3290 24070 3292
rect 24126 3290 24150 3292
rect 24206 3290 24212 3292
rect 23966 3238 23968 3290
rect 24148 3238 24150 3290
rect 23904 3236 23910 3238
rect 23966 3236 23990 3238
rect 24046 3236 24070 3238
rect 24126 3236 24150 3238
rect 24206 3236 24212 3238
rect 23904 3227 24212 3236
rect 27262 2748 27570 2757
rect 27262 2746 27268 2748
rect 27324 2746 27348 2748
rect 27404 2746 27428 2748
rect 27484 2746 27508 2748
rect 27564 2746 27570 2748
rect 27324 2694 27326 2746
rect 27506 2694 27508 2746
rect 27262 2692 27268 2694
rect 27324 2692 27348 2694
rect 27404 2692 27428 2694
rect 27484 2692 27508 2694
rect 27564 2692 27570 2694
rect 27262 2683 27570 2692
rect 23904 2204 24212 2213
rect 23904 2202 23910 2204
rect 23966 2202 23990 2204
rect 24046 2202 24070 2204
rect 24126 2202 24150 2204
rect 24206 2202 24212 2204
rect 23966 2150 23968 2202
rect 24148 2150 24150 2202
rect 23904 2148 23910 2150
rect 23966 2148 23990 2150
rect 24046 2148 24070 2150
rect 24126 2148 24150 2150
rect 24206 2148 24212 2150
rect 23904 2139 24212 2148
rect 23572 1828 23624 1834
rect 23572 1770 23624 1776
rect 22006 1391 22008 1400
rect 22060 1391 22062 1400
rect 22928 1420 22980 1426
rect 22008 1362 22060 1368
rect 22928 1362 22980 1368
rect 23584 400 23612 1770
rect 27262 1660 27570 1669
rect 27262 1658 27268 1660
rect 27324 1658 27348 1660
rect 27404 1658 27428 1660
rect 27484 1658 27508 1660
rect 27564 1658 27570 1660
rect 27324 1606 27326 1658
rect 27506 1606 27508 1658
rect 27262 1604 27268 1606
rect 27324 1604 27348 1606
rect 27404 1604 27428 1606
rect 27484 1604 27508 1606
rect 27564 1604 27570 1606
rect 27262 1595 27570 1604
rect 25320 1488 25372 1494
rect 25320 1430 25372 1436
rect 23904 1116 24212 1125
rect 23904 1114 23910 1116
rect 23966 1114 23990 1116
rect 24046 1114 24070 1116
rect 24126 1114 24150 1116
rect 24206 1114 24212 1116
rect 23966 1062 23968 1114
rect 24148 1062 24150 1114
rect 23904 1060 23910 1062
rect 23966 1060 23990 1062
rect 24046 1060 24070 1062
rect 24126 1060 24150 1062
rect 24206 1060 24212 1062
rect 23904 1051 24212 1060
rect 25332 400 25360 1430
rect 27068 740 27120 746
rect 27068 682 27120 688
rect 27080 400 27108 682
rect 27262 572 27570 581
rect 27262 570 27268 572
rect 27324 570 27348 572
rect 27404 570 27428 572
rect 27484 570 27508 572
rect 27564 570 27570 572
rect 27324 518 27326 570
rect 27506 518 27508 570
rect 27262 516 27268 518
rect 27324 516 27348 518
rect 27404 516 27428 518
rect 27484 516 27508 518
rect 27564 516 27570 518
rect 27262 507 27570 516
rect 846 0 902 400
rect 2594 0 2650 400
rect 4342 0 4398 400
rect 6090 0 6146 400
rect 7838 0 7894 400
rect 9586 0 9642 400
rect 11334 0 11390 400
rect 13082 0 13138 400
rect 14830 0 14886 400
rect 16578 0 16634 400
rect 18326 0 18382 400
rect 20074 0 20130 400
rect 21822 0 21878 400
rect 23570 0 23626 400
rect 25318 0 25374 400
rect 27066 0 27122 400
<< via2 >>
rect 3762 17434 3818 17436
rect 3842 17434 3898 17436
rect 3922 17434 3978 17436
rect 4002 17434 4058 17436
rect 3762 17382 3808 17434
rect 3808 17382 3818 17434
rect 3842 17382 3872 17434
rect 3872 17382 3884 17434
rect 3884 17382 3898 17434
rect 3922 17382 3936 17434
rect 3936 17382 3948 17434
rect 3948 17382 3978 17434
rect 4002 17382 4012 17434
rect 4012 17382 4058 17434
rect 3762 17380 3818 17382
rect 3842 17380 3898 17382
rect 3922 17380 3978 17382
rect 4002 17380 4058 17382
rect 7120 16890 7176 16892
rect 7200 16890 7256 16892
rect 7280 16890 7336 16892
rect 7360 16890 7416 16892
rect 7120 16838 7166 16890
rect 7166 16838 7176 16890
rect 7200 16838 7230 16890
rect 7230 16838 7242 16890
rect 7242 16838 7256 16890
rect 7280 16838 7294 16890
rect 7294 16838 7306 16890
rect 7306 16838 7336 16890
rect 7360 16838 7370 16890
rect 7370 16838 7416 16890
rect 7120 16836 7176 16838
rect 7200 16836 7256 16838
rect 7280 16836 7336 16838
rect 7360 16836 7416 16838
rect 3762 16346 3818 16348
rect 3842 16346 3898 16348
rect 3922 16346 3978 16348
rect 4002 16346 4058 16348
rect 3762 16294 3808 16346
rect 3808 16294 3818 16346
rect 3842 16294 3872 16346
rect 3872 16294 3884 16346
rect 3884 16294 3898 16346
rect 3922 16294 3936 16346
rect 3936 16294 3948 16346
rect 3948 16294 3978 16346
rect 4002 16294 4012 16346
rect 4012 16294 4058 16346
rect 3762 16292 3818 16294
rect 3842 16292 3898 16294
rect 3922 16292 3978 16294
rect 4002 16292 4058 16294
rect 3762 15258 3818 15260
rect 3842 15258 3898 15260
rect 3922 15258 3978 15260
rect 4002 15258 4058 15260
rect 3762 15206 3808 15258
rect 3808 15206 3818 15258
rect 3842 15206 3872 15258
rect 3872 15206 3884 15258
rect 3884 15206 3898 15258
rect 3922 15206 3936 15258
rect 3936 15206 3948 15258
rect 3948 15206 3978 15258
rect 4002 15206 4012 15258
rect 4012 15206 4058 15258
rect 3762 15204 3818 15206
rect 3842 15204 3898 15206
rect 3922 15204 3978 15206
rect 4002 15204 4058 15206
rect 3762 14170 3818 14172
rect 3842 14170 3898 14172
rect 3922 14170 3978 14172
rect 4002 14170 4058 14172
rect 3762 14118 3808 14170
rect 3808 14118 3818 14170
rect 3842 14118 3872 14170
rect 3872 14118 3884 14170
rect 3884 14118 3898 14170
rect 3922 14118 3936 14170
rect 3936 14118 3948 14170
rect 3948 14118 3978 14170
rect 4002 14118 4012 14170
rect 4012 14118 4058 14170
rect 3762 14116 3818 14118
rect 3842 14116 3898 14118
rect 3922 14116 3978 14118
rect 4002 14116 4058 14118
rect 3762 13082 3818 13084
rect 3842 13082 3898 13084
rect 3922 13082 3978 13084
rect 4002 13082 4058 13084
rect 3762 13030 3808 13082
rect 3808 13030 3818 13082
rect 3842 13030 3872 13082
rect 3872 13030 3884 13082
rect 3884 13030 3898 13082
rect 3922 13030 3936 13082
rect 3936 13030 3948 13082
rect 3948 13030 3978 13082
rect 4002 13030 4012 13082
rect 4012 13030 4058 13082
rect 3762 13028 3818 13030
rect 3842 13028 3898 13030
rect 3922 13028 3978 13030
rect 4002 13028 4058 13030
rect 3422 12824 3478 12880
rect 6182 13912 6238 13968
rect 4710 12860 4712 12880
rect 4712 12860 4764 12880
rect 4764 12860 4766 12880
rect 4710 12824 4766 12860
rect 7120 15802 7176 15804
rect 7200 15802 7256 15804
rect 7280 15802 7336 15804
rect 7360 15802 7416 15804
rect 7120 15750 7166 15802
rect 7166 15750 7176 15802
rect 7200 15750 7230 15802
rect 7230 15750 7242 15802
rect 7242 15750 7256 15802
rect 7280 15750 7294 15802
rect 7294 15750 7306 15802
rect 7306 15750 7336 15802
rect 7360 15750 7370 15802
rect 7370 15750 7416 15802
rect 7120 15748 7176 15750
rect 7200 15748 7256 15750
rect 7280 15748 7336 15750
rect 7360 15748 7416 15750
rect 7120 14714 7176 14716
rect 7200 14714 7256 14716
rect 7280 14714 7336 14716
rect 7360 14714 7416 14716
rect 7120 14662 7166 14714
rect 7166 14662 7176 14714
rect 7200 14662 7230 14714
rect 7230 14662 7242 14714
rect 7242 14662 7256 14714
rect 7280 14662 7294 14714
rect 7294 14662 7306 14714
rect 7306 14662 7336 14714
rect 7360 14662 7370 14714
rect 7370 14662 7416 14714
rect 7120 14660 7176 14662
rect 7200 14660 7256 14662
rect 7280 14660 7336 14662
rect 7360 14660 7416 14662
rect 7120 13626 7176 13628
rect 7200 13626 7256 13628
rect 7280 13626 7336 13628
rect 7360 13626 7416 13628
rect 7120 13574 7166 13626
rect 7166 13574 7176 13626
rect 7200 13574 7230 13626
rect 7230 13574 7242 13626
rect 7242 13574 7256 13626
rect 7280 13574 7294 13626
rect 7294 13574 7306 13626
rect 7306 13574 7336 13626
rect 7360 13574 7370 13626
rect 7370 13574 7416 13626
rect 7120 13572 7176 13574
rect 7200 13572 7256 13574
rect 7280 13572 7336 13574
rect 7360 13572 7416 13574
rect 3762 11994 3818 11996
rect 3842 11994 3898 11996
rect 3922 11994 3978 11996
rect 4002 11994 4058 11996
rect 3762 11942 3808 11994
rect 3808 11942 3818 11994
rect 3842 11942 3872 11994
rect 3872 11942 3884 11994
rect 3884 11942 3898 11994
rect 3922 11942 3936 11994
rect 3936 11942 3948 11994
rect 3948 11942 3978 11994
rect 4002 11942 4012 11994
rect 4012 11942 4058 11994
rect 3762 11940 3818 11942
rect 3842 11940 3898 11942
rect 3922 11940 3978 11942
rect 4002 11940 4058 11942
rect 7120 12538 7176 12540
rect 7200 12538 7256 12540
rect 7280 12538 7336 12540
rect 7360 12538 7416 12540
rect 7120 12486 7166 12538
rect 7166 12486 7176 12538
rect 7200 12486 7230 12538
rect 7230 12486 7242 12538
rect 7242 12486 7256 12538
rect 7280 12486 7294 12538
rect 7294 12486 7306 12538
rect 7306 12486 7336 12538
rect 7360 12486 7370 12538
rect 7370 12486 7416 12538
rect 7120 12484 7176 12486
rect 7200 12484 7256 12486
rect 7280 12484 7336 12486
rect 7360 12484 7416 12486
rect 10478 17434 10534 17436
rect 10558 17434 10614 17436
rect 10638 17434 10694 17436
rect 10718 17434 10774 17436
rect 10478 17382 10524 17434
rect 10524 17382 10534 17434
rect 10558 17382 10588 17434
rect 10588 17382 10600 17434
rect 10600 17382 10614 17434
rect 10638 17382 10652 17434
rect 10652 17382 10664 17434
rect 10664 17382 10694 17434
rect 10718 17382 10728 17434
rect 10728 17382 10774 17434
rect 10478 17380 10534 17382
rect 10558 17380 10614 17382
rect 10638 17380 10694 17382
rect 10718 17380 10774 17382
rect 10478 16346 10534 16348
rect 10558 16346 10614 16348
rect 10638 16346 10694 16348
rect 10718 16346 10774 16348
rect 10478 16294 10524 16346
rect 10524 16294 10534 16346
rect 10558 16294 10588 16346
rect 10588 16294 10600 16346
rect 10600 16294 10614 16346
rect 10638 16294 10652 16346
rect 10652 16294 10664 16346
rect 10664 16294 10694 16346
rect 10718 16294 10728 16346
rect 10728 16294 10774 16346
rect 10478 16292 10534 16294
rect 10558 16292 10614 16294
rect 10638 16292 10694 16294
rect 10718 16292 10774 16294
rect 7930 15000 7986 15056
rect 8206 13948 8208 13968
rect 8208 13948 8260 13968
rect 8260 13948 8262 13968
rect 8206 13912 8262 13948
rect 7470 12300 7526 12336
rect 7470 12280 7472 12300
rect 7472 12280 7524 12300
rect 7524 12280 7526 12300
rect 3762 10906 3818 10908
rect 3842 10906 3898 10908
rect 3922 10906 3978 10908
rect 4002 10906 4058 10908
rect 3762 10854 3808 10906
rect 3808 10854 3818 10906
rect 3842 10854 3872 10906
rect 3872 10854 3884 10906
rect 3884 10854 3898 10906
rect 3922 10854 3936 10906
rect 3936 10854 3948 10906
rect 3948 10854 3978 10906
rect 4002 10854 4012 10906
rect 4012 10854 4058 10906
rect 3762 10852 3818 10854
rect 3842 10852 3898 10854
rect 3922 10852 3978 10854
rect 4002 10852 4058 10854
rect 3762 9818 3818 9820
rect 3842 9818 3898 9820
rect 3922 9818 3978 9820
rect 4002 9818 4058 9820
rect 3762 9766 3808 9818
rect 3808 9766 3818 9818
rect 3842 9766 3872 9818
rect 3872 9766 3884 9818
rect 3884 9766 3898 9818
rect 3922 9766 3936 9818
rect 3936 9766 3948 9818
rect 3948 9766 3978 9818
rect 4002 9766 4012 9818
rect 4012 9766 4058 9818
rect 3762 9764 3818 9766
rect 3842 9764 3898 9766
rect 3922 9764 3978 9766
rect 4002 9764 4058 9766
rect 5170 9052 5172 9072
rect 5172 9052 5224 9072
rect 5224 9052 5226 9072
rect 5170 9016 5226 9052
rect 3762 8730 3818 8732
rect 3842 8730 3898 8732
rect 3922 8730 3978 8732
rect 4002 8730 4058 8732
rect 3762 8678 3808 8730
rect 3808 8678 3818 8730
rect 3842 8678 3872 8730
rect 3872 8678 3884 8730
rect 3884 8678 3898 8730
rect 3922 8678 3936 8730
rect 3936 8678 3948 8730
rect 3948 8678 3978 8730
rect 4002 8678 4012 8730
rect 4012 8678 4058 8730
rect 3762 8676 3818 8678
rect 3842 8676 3898 8678
rect 3922 8676 3978 8678
rect 4002 8676 4058 8678
rect 3514 8336 3570 8392
rect 3762 7642 3818 7644
rect 3842 7642 3898 7644
rect 3922 7642 3978 7644
rect 4002 7642 4058 7644
rect 3762 7590 3808 7642
rect 3808 7590 3818 7642
rect 3842 7590 3872 7642
rect 3872 7590 3884 7642
rect 3884 7590 3898 7642
rect 3922 7590 3936 7642
rect 3936 7590 3948 7642
rect 3948 7590 3978 7642
rect 4002 7590 4012 7642
rect 4012 7590 4058 7642
rect 3762 7588 3818 7590
rect 3842 7588 3898 7590
rect 3922 7588 3978 7590
rect 4002 7588 4058 7590
rect 3762 6554 3818 6556
rect 3842 6554 3898 6556
rect 3922 6554 3978 6556
rect 4002 6554 4058 6556
rect 3762 6502 3808 6554
rect 3808 6502 3818 6554
rect 3842 6502 3872 6554
rect 3872 6502 3884 6554
rect 3884 6502 3898 6554
rect 3922 6502 3936 6554
rect 3936 6502 3948 6554
rect 3948 6502 3978 6554
rect 4002 6502 4012 6554
rect 4012 6502 4058 6554
rect 3762 6500 3818 6502
rect 3842 6500 3898 6502
rect 3922 6500 3978 6502
rect 4002 6500 4058 6502
rect 7120 11450 7176 11452
rect 7200 11450 7256 11452
rect 7280 11450 7336 11452
rect 7360 11450 7416 11452
rect 7120 11398 7166 11450
rect 7166 11398 7176 11450
rect 7200 11398 7230 11450
rect 7230 11398 7242 11450
rect 7242 11398 7256 11450
rect 7280 11398 7294 11450
rect 7294 11398 7306 11450
rect 7306 11398 7336 11450
rect 7360 11398 7370 11450
rect 7370 11398 7416 11450
rect 7120 11396 7176 11398
rect 7200 11396 7256 11398
rect 7280 11396 7336 11398
rect 7360 11396 7416 11398
rect 3762 5466 3818 5468
rect 3842 5466 3898 5468
rect 3922 5466 3978 5468
rect 4002 5466 4058 5468
rect 3762 5414 3808 5466
rect 3808 5414 3818 5466
rect 3842 5414 3872 5466
rect 3872 5414 3884 5466
rect 3884 5414 3898 5466
rect 3922 5414 3936 5466
rect 3936 5414 3948 5466
rect 3948 5414 3978 5466
rect 4002 5414 4012 5466
rect 4012 5414 4058 5466
rect 3762 5412 3818 5414
rect 3842 5412 3898 5414
rect 3922 5412 3978 5414
rect 4002 5412 4058 5414
rect 3762 4378 3818 4380
rect 3842 4378 3898 4380
rect 3922 4378 3978 4380
rect 4002 4378 4058 4380
rect 3762 4326 3808 4378
rect 3808 4326 3818 4378
rect 3842 4326 3872 4378
rect 3872 4326 3884 4378
rect 3884 4326 3898 4378
rect 3922 4326 3936 4378
rect 3936 4326 3948 4378
rect 3948 4326 3978 4378
rect 4002 4326 4012 4378
rect 4012 4326 4058 4378
rect 3762 4324 3818 4326
rect 3842 4324 3898 4326
rect 3922 4324 3978 4326
rect 4002 4324 4058 4326
rect 3762 3290 3818 3292
rect 3842 3290 3898 3292
rect 3922 3290 3978 3292
rect 4002 3290 4058 3292
rect 3762 3238 3808 3290
rect 3808 3238 3818 3290
rect 3842 3238 3872 3290
rect 3872 3238 3884 3290
rect 3884 3238 3898 3290
rect 3922 3238 3936 3290
rect 3936 3238 3948 3290
rect 3948 3238 3978 3290
rect 4002 3238 4012 3290
rect 4012 3238 4058 3290
rect 3762 3236 3818 3238
rect 3842 3236 3898 3238
rect 3922 3236 3978 3238
rect 4002 3236 4058 3238
rect 3762 2202 3818 2204
rect 3842 2202 3898 2204
rect 3922 2202 3978 2204
rect 4002 2202 4058 2204
rect 3762 2150 3808 2202
rect 3808 2150 3818 2202
rect 3842 2150 3872 2202
rect 3872 2150 3884 2202
rect 3884 2150 3898 2202
rect 3922 2150 3936 2202
rect 3936 2150 3948 2202
rect 3948 2150 3978 2202
rect 4002 2150 4012 2202
rect 4012 2150 4058 2202
rect 3762 2148 3818 2150
rect 3842 2148 3898 2150
rect 3922 2148 3978 2150
rect 4002 2148 4058 2150
rect 846 1808 902 1864
rect 6366 6180 6422 6216
rect 6366 6160 6368 6180
rect 6368 6160 6420 6180
rect 6420 6160 6422 6180
rect 5998 1944 6054 2000
rect 3762 1114 3818 1116
rect 3842 1114 3898 1116
rect 3922 1114 3978 1116
rect 4002 1114 4058 1116
rect 3762 1062 3808 1114
rect 3808 1062 3818 1114
rect 3842 1062 3872 1114
rect 3872 1062 3884 1114
rect 3884 1062 3898 1114
rect 3922 1062 3936 1114
rect 3936 1062 3948 1114
rect 3948 1062 3978 1114
rect 4002 1062 4012 1114
rect 4012 1062 4058 1114
rect 3762 1060 3818 1062
rect 3842 1060 3898 1062
rect 3922 1060 3978 1062
rect 4002 1060 4058 1062
rect 7120 10362 7176 10364
rect 7200 10362 7256 10364
rect 7280 10362 7336 10364
rect 7360 10362 7416 10364
rect 7120 10310 7166 10362
rect 7166 10310 7176 10362
rect 7200 10310 7230 10362
rect 7230 10310 7242 10362
rect 7242 10310 7256 10362
rect 7280 10310 7294 10362
rect 7294 10310 7306 10362
rect 7306 10310 7336 10362
rect 7360 10310 7370 10362
rect 7370 10310 7416 10362
rect 7120 10308 7176 10310
rect 7200 10308 7256 10310
rect 7280 10308 7336 10310
rect 7360 10308 7416 10310
rect 7746 11600 7802 11656
rect 7838 11192 7894 11248
rect 7120 9274 7176 9276
rect 7200 9274 7256 9276
rect 7280 9274 7336 9276
rect 7360 9274 7416 9276
rect 7120 9222 7166 9274
rect 7166 9222 7176 9274
rect 7200 9222 7230 9274
rect 7230 9222 7242 9274
rect 7242 9222 7256 9274
rect 7280 9222 7294 9274
rect 7294 9222 7306 9274
rect 7306 9222 7336 9274
rect 7360 9222 7370 9274
rect 7370 9222 7416 9274
rect 7120 9220 7176 9222
rect 7200 9220 7256 9222
rect 7280 9220 7336 9222
rect 7360 9220 7416 9222
rect 7120 8186 7176 8188
rect 7200 8186 7256 8188
rect 7280 8186 7336 8188
rect 7360 8186 7416 8188
rect 7120 8134 7166 8186
rect 7166 8134 7176 8186
rect 7200 8134 7230 8186
rect 7230 8134 7242 8186
rect 7242 8134 7256 8186
rect 7280 8134 7294 8186
rect 7294 8134 7306 8186
rect 7306 8134 7336 8186
rect 7360 8134 7370 8186
rect 7370 8134 7416 8186
rect 7120 8132 7176 8134
rect 7200 8132 7256 8134
rect 7280 8132 7336 8134
rect 7360 8132 7416 8134
rect 7120 7098 7176 7100
rect 7200 7098 7256 7100
rect 7280 7098 7336 7100
rect 7360 7098 7416 7100
rect 7120 7046 7166 7098
rect 7166 7046 7176 7098
rect 7200 7046 7230 7098
rect 7230 7046 7242 7098
rect 7242 7046 7256 7098
rect 7280 7046 7294 7098
rect 7294 7046 7306 7098
rect 7306 7046 7336 7098
rect 7360 7046 7370 7098
rect 7370 7046 7416 7098
rect 7120 7044 7176 7046
rect 7200 7044 7256 7046
rect 7280 7044 7336 7046
rect 7360 7044 7416 7046
rect 7120 6010 7176 6012
rect 7200 6010 7256 6012
rect 7280 6010 7336 6012
rect 7360 6010 7416 6012
rect 7120 5958 7166 6010
rect 7166 5958 7176 6010
rect 7200 5958 7230 6010
rect 7230 5958 7242 6010
rect 7242 5958 7256 6010
rect 7280 5958 7294 6010
rect 7294 5958 7306 6010
rect 7306 5958 7336 6010
rect 7360 5958 7370 6010
rect 7370 5958 7416 6010
rect 7120 5956 7176 5958
rect 7200 5956 7256 5958
rect 7280 5956 7336 5958
rect 7360 5956 7416 5958
rect 7120 4922 7176 4924
rect 7200 4922 7256 4924
rect 7280 4922 7336 4924
rect 7360 4922 7416 4924
rect 7120 4870 7166 4922
rect 7166 4870 7176 4922
rect 7200 4870 7230 4922
rect 7230 4870 7242 4922
rect 7242 4870 7256 4922
rect 7280 4870 7294 4922
rect 7294 4870 7306 4922
rect 7306 4870 7336 4922
rect 7360 4870 7370 4922
rect 7370 4870 7416 4922
rect 7120 4868 7176 4870
rect 7200 4868 7256 4870
rect 7280 4868 7336 4870
rect 7360 4868 7416 4870
rect 6458 2488 6514 2544
rect 9862 14492 9864 14512
rect 9864 14492 9916 14512
rect 9916 14492 9918 14512
rect 9862 14456 9918 14492
rect 10322 15272 10378 15328
rect 10478 15258 10534 15260
rect 10558 15258 10614 15260
rect 10638 15258 10694 15260
rect 10718 15258 10774 15260
rect 10478 15206 10524 15258
rect 10524 15206 10534 15258
rect 10558 15206 10588 15258
rect 10588 15206 10600 15258
rect 10600 15206 10614 15258
rect 10638 15206 10652 15258
rect 10652 15206 10664 15258
rect 10664 15206 10694 15258
rect 10718 15206 10728 15258
rect 10728 15206 10774 15258
rect 10478 15204 10534 15206
rect 10558 15204 10614 15206
rect 10638 15204 10694 15206
rect 10718 15204 10774 15206
rect 10478 14170 10534 14172
rect 10558 14170 10614 14172
rect 10638 14170 10694 14172
rect 10718 14170 10774 14172
rect 10478 14118 10524 14170
rect 10524 14118 10534 14170
rect 10558 14118 10588 14170
rect 10588 14118 10600 14170
rect 10600 14118 10614 14170
rect 10638 14118 10652 14170
rect 10652 14118 10664 14170
rect 10664 14118 10694 14170
rect 10718 14118 10728 14170
rect 10728 14118 10774 14170
rect 10478 14116 10534 14118
rect 10558 14116 10614 14118
rect 10638 14116 10694 14118
rect 10718 14116 10774 14118
rect 9586 11328 9642 11384
rect 10478 13082 10534 13084
rect 10558 13082 10614 13084
rect 10638 13082 10694 13084
rect 10718 13082 10774 13084
rect 10478 13030 10524 13082
rect 10524 13030 10534 13082
rect 10558 13030 10588 13082
rect 10588 13030 10600 13082
rect 10600 13030 10614 13082
rect 10638 13030 10652 13082
rect 10652 13030 10664 13082
rect 10664 13030 10694 13082
rect 10718 13030 10728 13082
rect 10728 13030 10774 13082
rect 10478 13028 10534 13030
rect 10558 13028 10614 13030
rect 10638 13028 10694 13030
rect 10718 13028 10774 13030
rect 10046 12280 10102 12336
rect 7120 3834 7176 3836
rect 7200 3834 7256 3836
rect 7280 3834 7336 3836
rect 7360 3834 7416 3836
rect 7120 3782 7166 3834
rect 7166 3782 7176 3834
rect 7200 3782 7230 3834
rect 7230 3782 7242 3834
rect 7242 3782 7256 3834
rect 7280 3782 7294 3834
rect 7294 3782 7306 3834
rect 7306 3782 7336 3834
rect 7360 3782 7370 3834
rect 7370 3782 7416 3834
rect 7120 3780 7176 3782
rect 7200 3780 7256 3782
rect 7280 3780 7336 3782
rect 7360 3780 7416 3782
rect 7120 2746 7176 2748
rect 7200 2746 7256 2748
rect 7280 2746 7336 2748
rect 7360 2746 7416 2748
rect 7120 2694 7166 2746
rect 7166 2694 7176 2746
rect 7200 2694 7230 2746
rect 7230 2694 7242 2746
rect 7242 2694 7256 2746
rect 7280 2694 7294 2746
rect 7294 2694 7306 2746
rect 7306 2694 7336 2746
rect 7360 2694 7370 2746
rect 7370 2694 7416 2746
rect 7120 2692 7176 2694
rect 7200 2692 7256 2694
rect 7280 2692 7336 2694
rect 7360 2692 7416 2694
rect 7120 1658 7176 1660
rect 7200 1658 7256 1660
rect 7280 1658 7336 1660
rect 7360 1658 7416 1660
rect 7120 1606 7166 1658
rect 7166 1606 7176 1658
rect 7200 1606 7230 1658
rect 7230 1606 7242 1658
rect 7242 1606 7256 1658
rect 7280 1606 7294 1658
rect 7294 1606 7306 1658
rect 7306 1606 7336 1658
rect 7360 1606 7370 1658
rect 7370 1606 7416 1658
rect 7120 1604 7176 1606
rect 7200 1604 7256 1606
rect 7280 1604 7336 1606
rect 7360 1604 7416 1606
rect 7470 1400 7526 1456
rect 7930 1400 7986 1456
rect 7120 570 7176 572
rect 7200 570 7256 572
rect 7280 570 7336 572
rect 7360 570 7416 572
rect 7120 518 7166 570
rect 7166 518 7176 570
rect 7200 518 7230 570
rect 7230 518 7242 570
rect 7242 518 7256 570
rect 7280 518 7294 570
rect 7294 518 7306 570
rect 7306 518 7336 570
rect 7360 518 7370 570
rect 7370 518 7416 570
rect 7120 516 7176 518
rect 7200 516 7256 518
rect 7280 516 7336 518
rect 7360 516 7416 518
rect 8850 4664 8906 4720
rect 9218 6840 9274 6896
rect 9862 7812 9918 7848
rect 9862 7792 9864 7812
rect 9864 7792 9916 7812
rect 9916 7792 9918 7812
rect 9402 6840 9458 6896
rect 9310 4684 9366 4720
rect 9310 4664 9312 4684
rect 9312 4664 9364 4684
rect 9364 4664 9366 4684
rect 10478 11994 10534 11996
rect 10558 11994 10614 11996
rect 10638 11994 10694 11996
rect 10718 11994 10774 11996
rect 10478 11942 10524 11994
rect 10524 11942 10534 11994
rect 10558 11942 10588 11994
rect 10588 11942 10600 11994
rect 10600 11942 10614 11994
rect 10638 11942 10652 11994
rect 10652 11942 10664 11994
rect 10664 11942 10694 11994
rect 10718 11942 10728 11994
rect 10728 11942 10774 11994
rect 10478 11940 10534 11942
rect 10558 11940 10614 11942
rect 10638 11940 10694 11942
rect 10718 11940 10774 11942
rect 10478 10906 10534 10908
rect 10558 10906 10614 10908
rect 10638 10906 10694 10908
rect 10718 10906 10774 10908
rect 10478 10854 10524 10906
rect 10524 10854 10534 10906
rect 10558 10854 10588 10906
rect 10588 10854 10600 10906
rect 10600 10854 10614 10906
rect 10638 10854 10652 10906
rect 10652 10854 10664 10906
rect 10664 10854 10694 10906
rect 10718 10854 10728 10906
rect 10728 10854 10774 10906
rect 10478 10852 10534 10854
rect 10558 10852 10614 10854
rect 10638 10852 10694 10854
rect 10718 10852 10774 10854
rect 10478 9818 10534 9820
rect 10558 9818 10614 9820
rect 10638 9818 10694 9820
rect 10718 9818 10774 9820
rect 10478 9766 10524 9818
rect 10524 9766 10534 9818
rect 10558 9766 10588 9818
rect 10588 9766 10600 9818
rect 10600 9766 10614 9818
rect 10638 9766 10652 9818
rect 10652 9766 10664 9818
rect 10664 9766 10694 9818
rect 10718 9766 10728 9818
rect 10728 9766 10774 9818
rect 10478 9764 10534 9766
rect 10558 9764 10614 9766
rect 10638 9764 10694 9766
rect 10718 9764 10774 9766
rect 10478 8730 10534 8732
rect 10558 8730 10614 8732
rect 10638 8730 10694 8732
rect 10718 8730 10774 8732
rect 10478 8678 10524 8730
rect 10524 8678 10534 8730
rect 10558 8678 10588 8730
rect 10588 8678 10600 8730
rect 10600 8678 10614 8730
rect 10638 8678 10652 8730
rect 10652 8678 10664 8730
rect 10664 8678 10694 8730
rect 10718 8678 10728 8730
rect 10728 8678 10774 8730
rect 10478 8676 10534 8678
rect 10558 8676 10614 8678
rect 10638 8676 10694 8678
rect 10718 8676 10774 8678
rect 10478 7642 10534 7644
rect 10558 7642 10614 7644
rect 10638 7642 10694 7644
rect 10718 7642 10774 7644
rect 10478 7590 10524 7642
rect 10524 7590 10534 7642
rect 10558 7590 10588 7642
rect 10588 7590 10600 7642
rect 10600 7590 10614 7642
rect 10638 7590 10652 7642
rect 10652 7590 10664 7642
rect 10664 7590 10694 7642
rect 10718 7590 10728 7642
rect 10728 7590 10774 7642
rect 10478 7588 10534 7590
rect 10558 7588 10614 7590
rect 10638 7588 10694 7590
rect 10718 7588 10774 7590
rect 10478 6554 10534 6556
rect 10558 6554 10614 6556
rect 10638 6554 10694 6556
rect 10718 6554 10774 6556
rect 10478 6502 10524 6554
rect 10524 6502 10534 6554
rect 10558 6502 10588 6554
rect 10588 6502 10600 6554
rect 10600 6502 10614 6554
rect 10638 6502 10652 6554
rect 10652 6502 10664 6554
rect 10664 6502 10694 6554
rect 10718 6502 10728 6554
rect 10728 6502 10774 6554
rect 10478 6500 10534 6502
rect 10558 6500 10614 6502
rect 10638 6500 10694 6502
rect 10718 6500 10774 6502
rect 10598 6296 10654 6352
rect 10782 5636 10838 5672
rect 10782 5616 10784 5636
rect 10784 5616 10836 5636
rect 10836 5616 10838 5636
rect 10478 5466 10534 5468
rect 10558 5466 10614 5468
rect 10638 5466 10694 5468
rect 10718 5466 10774 5468
rect 10478 5414 10524 5466
rect 10524 5414 10534 5466
rect 10558 5414 10588 5466
rect 10588 5414 10600 5466
rect 10600 5414 10614 5466
rect 10638 5414 10652 5466
rect 10652 5414 10664 5466
rect 10664 5414 10694 5466
rect 10718 5414 10728 5466
rect 10728 5414 10774 5466
rect 10478 5412 10534 5414
rect 10558 5412 10614 5414
rect 10638 5412 10694 5414
rect 10718 5412 10774 5414
rect 10478 4378 10534 4380
rect 10558 4378 10614 4380
rect 10638 4378 10694 4380
rect 10718 4378 10774 4380
rect 10478 4326 10524 4378
rect 10524 4326 10534 4378
rect 10558 4326 10588 4378
rect 10588 4326 10600 4378
rect 10600 4326 10614 4378
rect 10638 4326 10652 4378
rect 10652 4326 10664 4378
rect 10664 4326 10694 4378
rect 10718 4326 10728 4378
rect 10728 4326 10774 4378
rect 10478 4324 10534 4326
rect 10558 4324 10614 4326
rect 10638 4324 10694 4326
rect 10718 4324 10774 4326
rect 10478 3290 10534 3292
rect 10558 3290 10614 3292
rect 10638 3290 10694 3292
rect 10718 3290 10774 3292
rect 10478 3238 10524 3290
rect 10524 3238 10534 3290
rect 10558 3238 10588 3290
rect 10588 3238 10600 3290
rect 10600 3238 10614 3290
rect 10638 3238 10652 3290
rect 10652 3238 10664 3290
rect 10664 3238 10694 3290
rect 10718 3238 10728 3290
rect 10728 3238 10774 3290
rect 10478 3236 10534 3238
rect 10558 3236 10614 3238
rect 10638 3236 10694 3238
rect 10718 3236 10774 3238
rect 13836 16890 13892 16892
rect 13916 16890 13972 16892
rect 13996 16890 14052 16892
rect 14076 16890 14132 16892
rect 13836 16838 13882 16890
rect 13882 16838 13892 16890
rect 13916 16838 13946 16890
rect 13946 16838 13958 16890
rect 13958 16838 13972 16890
rect 13996 16838 14010 16890
rect 14010 16838 14022 16890
rect 14022 16838 14052 16890
rect 14076 16838 14086 16890
rect 14086 16838 14132 16890
rect 13836 16836 13892 16838
rect 13916 16836 13972 16838
rect 13996 16836 14052 16838
rect 14076 16836 14132 16838
rect 14002 16652 14058 16688
rect 14002 16632 14004 16652
rect 14004 16632 14056 16652
rect 14056 16632 14058 16652
rect 12714 15000 12770 15056
rect 11426 5208 11482 5264
rect 12438 11328 12494 11384
rect 12438 9560 12494 9616
rect 12070 8472 12126 8528
rect 12438 9324 12440 9344
rect 12440 9324 12492 9344
rect 12492 9324 12494 9344
rect 12438 9288 12494 9324
rect 11886 6296 11942 6352
rect 8942 2352 8998 2408
rect 10478 2202 10534 2204
rect 10558 2202 10614 2204
rect 10638 2202 10694 2204
rect 10718 2202 10774 2204
rect 10478 2150 10524 2202
rect 10524 2150 10534 2202
rect 10558 2150 10588 2202
rect 10588 2150 10600 2202
rect 10600 2150 10614 2202
rect 10638 2150 10652 2202
rect 10652 2150 10664 2202
rect 10664 2150 10694 2202
rect 10718 2150 10728 2202
rect 10728 2150 10774 2202
rect 10478 2148 10534 2150
rect 10558 2148 10614 2150
rect 10638 2148 10694 2150
rect 10718 2148 10774 2150
rect 10478 1114 10534 1116
rect 10558 1114 10614 1116
rect 10638 1114 10694 1116
rect 10718 1114 10774 1116
rect 10478 1062 10524 1114
rect 10524 1062 10534 1114
rect 10558 1062 10588 1114
rect 10588 1062 10600 1114
rect 10600 1062 10614 1114
rect 10638 1062 10652 1114
rect 10652 1062 10664 1114
rect 10664 1062 10694 1114
rect 10718 1062 10728 1114
rect 10728 1062 10774 1114
rect 10478 1060 10534 1062
rect 10558 1060 10614 1062
rect 10638 1060 10694 1062
rect 10718 1060 10774 1062
rect 13836 15802 13892 15804
rect 13916 15802 13972 15804
rect 13996 15802 14052 15804
rect 14076 15802 14132 15804
rect 13836 15750 13882 15802
rect 13882 15750 13892 15802
rect 13916 15750 13946 15802
rect 13946 15750 13958 15802
rect 13958 15750 13972 15802
rect 13996 15750 14010 15802
rect 14010 15750 14022 15802
rect 14022 15750 14052 15802
rect 14076 15750 14086 15802
rect 14086 15750 14132 15802
rect 13836 15748 13892 15750
rect 13916 15748 13972 15750
rect 13996 15748 14052 15750
rect 14076 15748 14132 15750
rect 13836 14714 13892 14716
rect 13916 14714 13972 14716
rect 13996 14714 14052 14716
rect 14076 14714 14132 14716
rect 13836 14662 13882 14714
rect 13882 14662 13892 14714
rect 13916 14662 13946 14714
rect 13946 14662 13958 14714
rect 13958 14662 13972 14714
rect 13996 14662 14010 14714
rect 14010 14662 14022 14714
rect 14022 14662 14052 14714
rect 14076 14662 14086 14714
rect 14086 14662 14132 14714
rect 13836 14660 13892 14662
rect 13916 14660 13972 14662
rect 13996 14660 14052 14662
rect 14076 14660 14132 14662
rect 14002 14456 14058 14512
rect 13836 13626 13892 13628
rect 13916 13626 13972 13628
rect 13996 13626 14052 13628
rect 14076 13626 14132 13628
rect 13836 13574 13882 13626
rect 13882 13574 13892 13626
rect 13916 13574 13946 13626
rect 13946 13574 13958 13626
rect 13958 13574 13972 13626
rect 13996 13574 14010 13626
rect 14010 13574 14022 13626
rect 14022 13574 14052 13626
rect 14076 13574 14086 13626
rect 14086 13574 14132 13626
rect 13836 13572 13892 13574
rect 13916 13572 13972 13574
rect 13996 13572 14052 13574
rect 14076 13572 14132 13574
rect 13358 13096 13414 13152
rect 13836 12538 13892 12540
rect 13916 12538 13972 12540
rect 13996 12538 14052 12540
rect 14076 12538 14132 12540
rect 13836 12486 13882 12538
rect 13882 12486 13892 12538
rect 13916 12486 13946 12538
rect 13946 12486 13958 12538
rect 13958 12486 13972 12538
rect 13996 12486 14010 12538
rect 14010 12486 14022 12538
rect 14022 12486 14052 12538
rect 14076 12486 14086 12538
rect 14086 12486 14132 12538
rect 13836 12484 13892 12486
rect 13916 12484 13972 12486
rect 13996 12484 14052 12486
rect 14076 12484 14132 12486
rect 14094 11756 14150 11792
rect 14094 11736 14096 11756
rect 14096 11736 14148 11756
rect 14148 11736 14150 11756
rect 13836 11450 13892 11452
rect 13916 11450 13972 11452
rect 13996 11450 14052 11452
rect 14076 11450 14132 11452
rect 13836 11398 13882 11450
rect 13882 11398 13892 11450
rect 13916 11398 13946 11450
rect 13946 11398 13958 11450
rect 13958 11398 13972 11450
rect 13996 11398 14010 11450
rect 14010 11398 14022 11450
rect 14022 11398 14052 11450
rect 14076 11398 14086 11450
rect 14086 11398 14132 11450
rect 13836 11396 13892 11398
rect 13916 11396 13972 11398
rect 13996 11396 14052 11398
rect 14076 11396 14132 11398
rect 12806 6840 12862 6896
rect 13836 10362 13892 10364
rect 13916 10362 13972 10364
rect 13996 10362 14052 10364
rect 14076 10362 14132 10364
rect 13836 10310 13882 10362
rect 13882 10310 13892 10362
rect 13916 10310 13946 10362
rect 13946 10310 13958 10362
rect 13958 10310 13972 10362
rect 13996 10310 14010 10362
rect 14010 10310 14022 10362
rect 14022 10310 14052 10362
rect 14076 10310 14086 10362
rect 14086 10310 14132 10362
rect 13836 10308 13892 10310
rect 13916 10308 13972 10310
rect 13996 10308 14052 10310
rect 14076 10308 14132 10310
rect 13358 9288 13414 9344
rect 13836 9274 13892 9276
rect 13916 9274 13972 9276
rect 13996 9274 14052 9276
rect 14076 9274 14132 9276
rect 13836 9222 13882 9274
rect 13882 9222 13892 9274
rect 13916 9222 13946 9274
rect 13946 9222 13958 9274
rect 13958 9222 13972 9274
rect 13996 9222 14010 9274
rect 14010 9222 14022 9274
rect 14022 9222 14052 9274
rect 14076 9222 14086 9274
rect 14086 9222 14132 9274
rect 13836 9220 13892 9222
rect 13916 9220 13972 9222
rect 13996 9220 14052 9222
rect 14076 9220 14132 9222
rect 13836 8186 13892 8188
rect 13916 8186 13972 8188
rect 13996 8186 14052 8188
rect 14076 8186 14132 8188
rect 13836 8134 13882 8186
rect 13882 8134 13892 8186
rect 13916 8134 13946 8186
rect 13946 8134 13958 8186
rect 13958 8134 13972 8186
rect 13996 8134 14010 8186
rect 14010 8134 14022 8186
rect 14022 8134 14052 8186
rect 14076 8134 14086 8186
rect 14086 8134 14132 8186
rect 13836 8132 13892 8134
rect 13916 8132 13972 8134
rect 13996 8132 14052 8134
rect 14076 8132 14132 8134
rect 13818 7828 13820 7848
rect 13820 7828 13872 7848
rect 13872 7828 13874 7848
rect 13818 7792 13874 7828
rect 13836 7098 13892 7100
rect 13916 7098 13972 7100
rect 13996 7098 14052 7100
rect 14076 7098 14132 7100
rect 13836 7046 13882 7098
rect 13882 7046 13892 7098
rect 13916 7046 13946 7098
rect 13946 7046 13958 7098
rect 13958 7046 13972 7098
rect 13996 7046 14010 7098
rect 14010 7046 14022 7098
rect 14022 7046 14052 7098
rect 14076 7046 14086 7098
rect 14086 7046 14132 7098
rect 13836 7044 13892 7046
rect 13916 7044 13972 7046
rect 13996 7044 14052 7046
rect 14076 7044 14132 7046
rect 13836 6010 13892 6012
rect 13916 6010 13972 6012
rect 13996 6010 14052 6012
rect 14076 6010 14132 6012
rect 13836 5958 13882 6010
rect 13882 5958 13892 6010
rect 13916 5958 13946 6010
rect 13946 5958 13958 6010
rect 13958 5958 13972 6010
rect 13996 5958 14010 6010
rect 14010 5958 14022 6010
rect 14022 5958 14052 6010
rect 14076 5958 14086 6010
rect 14086 5958 14132 6010
rect 13836 5956 13892 5958
rect 13916 5956 13972 5958
rect 13996 5956 14052 5958
rect 14076 5956 14132 5958
rect 13836 4922 13892 4924
rect 13916 4922 13972 4924
rect 13996 4922 14052 4924
rect 14076 4922 14132 4924
rect 13836 4870 13882 4922
rect 13882 4870 13892 4922
rect 13916 4870 13946 4922
rect 13946 4870 13958 4922
rect 13958 4870 13972 4922
rect 13996 4870 14010 4922
rect 14010 4870 14022 4922
rect 14022 4870 14052 4922
rect 14076 4870 14086 4922
rect 14086 4870 14132 4922
rect 13836 4868 13892 4870
rect 13916 4868 13972 4870
rect 13996 4868 14052 4870
rect 14076 4868 14132 4870
rect 13836 3834 13892 3836
rect 13916 3834 13972 3836
rect 13996 3834 14052 3836
rect 14076 3834 14132 3836
rect 13836 3782 13882 3834
rect 13882 3782 13892 3834
rect 13916 3782 13946 3834
rect 13946 3782 13958 3834
rect 13958 3782 13972 3834
rect 13996 3782 14010 3834
rect 14010 3782 14022 3834
rect 14022 3782 14052 3834
rect 14076 3782 14086 3834
rect 14086 3782 14132 3834
rect 13836 3780 13892 3782
rect 13916 3780 13972 3782
rect 13996 3780 14052 3782
rect 14076 3780 14132 3782
rect 13836 2746 13892 2748
rect 13916 2746 13972 2748
rect 13996 2746 14052 2748
rect 14076 2746 14132 2748
rect 13836 2694 13882 2746
rect 13882 2694 13892 2746
rect 13916 2694 13946 2746
rect 13946 2694 13958 2746
rect 13958 2694 13972 2746
rect 13996 2694 14010 2746
rect 14010 2694 14022 2746
rect 14022 2694 14052 2746
rect 14076 2694 14086 2746
rect 14086 2694 14132 2746
rect 13836 2692 13892 2694
rect 13916 2692 13972 2694
rect 13996 2692 14052 2694
rect 14076 2692 14132 2694
rect 17194 17434 17250 17436
rect 17274 17434 17330 17436
rect 17354 17434 17410 17436
rect 17434 17434 17490 17436
rect 17194 17382 17240 17434
rect 17240 17382 17250 17434
rect 17274 17382 17304 17434
rect 17304 17382 17316 17434
rect 17316 17382 17330 17434
rect 17354 17382 17368 17434
rect 17368 17382 17380 17434
rect 17380 17382 17410 17434
rect 17434 17382 17444 17434
rect 17444 17382 17490 17434
rect 17194 17380 17250 17382
rect 17274 17380 17330 17382
rect 17354 17380 17410 17382
rect 17434 17380 17490 17382
rect 19522 17176 19578 17232
rect 23910 17434 23966 17436
rect 23990 17434 24046 17436
rect 24070 17434 24126 17436
rect 24150 17434 24206 17436
rect 23910 17382 23956 17434
rect 23956 17382 23966 17434
rect 23990 17382 24020 17434
rect 24020 17382 24032 17434
rect 24032 17382 24046 17434
rect 24070 17382 24084 17434
rect 24084 17382 24096 17434
rect 24096 17382 24126 17434
rect 24150 17382 24160 17434
rect 24160 17382 24206 17434
rect 23910 17380 23966 17382
rect 23990 17380 24046 17382
rect 24070 17380 24126 17382
rect 24150 17380 24206 17382
rect 24030 17212 24032 17232
rect 24032 17212 24084 17232
rect 24084 17212 24086 17232
rect 24030 17176 24086 17212
rect 14646 11056 14702 11112
rect 14462 9596 14464 9616
rect 14464 9596 14516 9616
rect 14516 9596 14518 9616
rect 14462 9560 14518 9596
rect 14462 6840 14518 6896
rect 14830 14476 14886 14512
rect 14830 14456 14832 14476
rect 14832 14456 14884 14476
rect 14884 14456 14886 14476
rect 15014 13388 15070 13424
rect 15014 13368 15016 13388
rect 15016 13368 15068 13388
rect 15068 13368 15070 13388
rect 14922 11600 14978 11656
rect 15106 11056 15162 11112
rect 15474 13096 15530 13152
rect 16210 13368 16266 13424
rect 15934 12300 15990 12336
rect 15934 12280 15936 12300
rect 15936 12280 15988 12300
rect 15988 12280 15990 12300
rect 15750 9444 15806 9480
rect 15750 9424 15752 9444
rect 15752 9424 15804 9444
rect 15804 9424 15806 9444
rect 16394 12280 16450 12336
rect 17194 16346 17250 16348
rect 17274 16346 17330 16348
rect 17354 16346 17410 16348
rect 17434 16346 17490 16348
rect 17194 16294 17240 16346
rect 17240 16294 17250 16346
rect 17274 16294 17304 16346
rect 17304 16294 17316 16346
rect 17316 16294 17330 16346
rect 17354 16294 17368 16346
rect 17368 16294 17380 16346
rect 17380 16294 17410 16346
rect 17434 16294 17444 16346
rect 17444 16294 17490 16346
rect 17194 16292 17250 16294
rect 17274 16292 17330 16294
rect 17354 16292 17410 16294
rect 17434 16292 17490 16294
rect 17194 15258 17250 15260
rect 17274 15258 17330 15260
rect 17354 15258 17410 15260
rect 17434 15258 17490 15260
rect 17194 15206 17240 15258
rect 17240 15206 17250 15258
rect 17274 15206 17304 15258
rect 17304 15206 17316 15258
rect 17316 15206 17330 15258
rect 17354 15206 17368 15258
rect 17368 15206 17380 15258
rect 17380 15206 17410 15258
rect 17434 15206 17444 15258
rect 17444 15206 17490 15258
rect 17194 15204 17250 15206
rect 17274 15204 17330 15206
rect 17354 15204 17410 15206
rect 17434 15204 17490 15206
rect 17194 14170 17250 14172
rect 17274 14170 17330 14172
rect 17354 14170 17410 14172
rect 17434 14170 17490 14172
rect 17194 14118 17240 14170
rect 17240 14118 17250 14170
rect 17274 14118 17304 14170
rect 17304 14118 17316 14170
rect 17316 14118 17330 14170
rect 17354 14118 17368 14170
rect 17368 14118 17380 14170
rect 17380 14118 17410 14170
rect 17434 14118 17444 14170
rect 17444 14118 17490 14170
rect 17194 14116 17250 14118
rect 17274 14116 17330 14118
rect 17354 14116 17410 14118
rect 17434 14116 17490 14118
rect 17194 13082 17250 13084
rect 17274 13082 17330 13084
rect 17354 13082 17410 13084
rect 17434 13082 17490 13084
rect 17194 13030 17240 13082
rect 17240 13030 17250 13082
rect 17274 13030 17304 13082
rect 17304 13030 17316 13082
rect 17316 13030 17330 13082
rect 17354 13030 17368 13082
rect 17368 13030 17380 13082
rect 17380 13030 17410 13082
rect 17434 13030 17444 13082
rect 17444 13030 17490 13082
rect 17194 13028 17250 13030
rect 17274 13028 17330 13030
rect 17354 13028 17410 13030
rect 17434 13028 17490 13030
rect 17194 11994 17250 11996
rect 17274 11994 17330 11996
rect 17354 11994 17410 11996
rect 17434 11994 17490 11996
rect 17194 11942 17240 11994
rect 17240 11942 17250 11994
rect 17274 11942 17304 11994
rect 17304 11942 17316 11994
rect 17316 11942 17330 11994
rect 17354 11942 17368 11994
rect 17368 11942 17380 11994
rect 17380 11942 17410 11994
rect 17434 11942 17444 11994
rect 17444 11942 17490 11994
rect 17194 11940 17250 11942
rect 17274 11940 17330 11942
rect 17354 11940 17410 11942
rect 17434 11940 17490 11942
rect 16578 11192 16634 11248
rect 17194 10906 17250 10908
rect 17274 10906 17330 10908
rect 17354 10906 17410 10908
rect 17434 10906 17490 10908
rect 17194 10854 17240 10906
rect 17240 10854 17250 10906
rect 17274 10854 17304 10906
rect 17304 10854 17316 10906
rect 17316 10854 17330 10906
rect 17354 10854 17368 10906
rect 17368 10854 17380 10906
rect 17380 10854 17410 10906
rect 17434 10854 17444 10906
rect 17444 10854 17490 10906
rect 17194 10852 17250 10854
rect 17274 10852 17330 10854
rect 17354 10852 17410 10854
rect 17434 10852 17490 10854
rect 17194 9818 17250 9820
rect 17274 9818 17330 9820
rect 17354 9818 17410 9820
rect 17434 9818 17490 9820
rect 17194 9766 17240 9818
rect 17240 9766 17250 9818
rect 17274 9766 17304 9818
rect 17304 9766 17316 9818
rect 17316 9766 17330 9818
rect 17354 9766 17368 9818
rect 17368 9766 17380 9818
rect 17380 9766 17410 9818
rect 17434 9766 17444 9818
rect 17444 9766 17490 9818
rect 17194 9764 17250 9766
rect 17274 9764 17330 9766
rect 17354 9764 17410 9766
rect 17434 9764 17490 9766
rect 16578 9016 16634 9072
rect 14646 2644 14702 2680
rect 14646 2624 14648 2644
rect 14648 2624 14700 2644
rect 14700 2624 14702 2644
rect 13836 1658 13892 1660
rect 13916 1658 13972 1660
rect 13996 1658 14052 1660
rect 14076 1658 14132 1660
rect 13836 1606 13882 1658
rect 13882 1606 13892 1658
rect 13916 1606 13946 1658
rect 13946 1606 13958 1658
rect 13958 1606 13972 1658
rect 13996 1606 14010 1658
rect 14010 1606 14022 1658
rect 14022 1606 14052 1658
rect 14076 1606 14086 1658
rect 14086 1606 14132 1658
rect 13836 1604 13892 1606
rect 13916 1604 13972 1606
rect 13996 1604 14052 1606
rect 14076 1604 14132 1606
rect 15290 1808 15346 1864
rect 13836 570 13892 572
rect 13916 570 13972 572
rect 13996 570 14052 572
rect 14076 570 14132 572
rect 13836 518 13882 570
rect 13882 518 13892 570
rect 13916 518 13946 570
rect 13946 518 13958 570
rect 13958 518 13972 570
rect 13996 518 14010 570
rect 14010 518 14022 570
rect 14022 518 14052 570
rect 14076 518 14086 570
rect 14086 518 14132 570
rect 13836 516 13892 518
rect 13916 516 13972 518
rect 13996 516 14052 518
rect 14076 516 14132 518
rect 17130 9016 17186 9072
rect 17194 8730 17250 8732
rect 17274 8730 17330 8732
rect 17354 8730 17410 8732
rect 17434 8730 17490 8732
rect 17194 8678 17240 8730
rect 17240 8678 17250 8730
rect 17274 8678 17304 8730
rect 17304 8678 17316 8730
rect 17316 8678 17330 8730
rect 17354 8678 17368 8730
rect 17368 8678 17380 8730
rect 17380 8678 17410 8730
rect 17434 8678 17444 8730
rect 17444 8678 17490 8730
rect 17194 8676 17250 8678
rect 17274 8676 17330 8678
rect 17354 8676 17410 8678
rect 17434 8676 17490 8678
rect 17590 8472 17646 8528
rect 17194 7642 17250 7644
rect 17274 7642 17330 7644
rect 17354 7642 17410 7644
rect 17434 7642 17490 7644
rect 17194 7590 17240 7642
rect 17240 7590 17250 7642
rect 17274 7590 17304 7642
rect 17304 7590 17316 7642
rect 17316 7590 17330 7642
rect 17354 7590 17368 7642
rect 17368 7590 17380 7642
rect 17380 7590 17410 7642
rect 17434 7590 17444 7642
rect 17444 7590 17490 7642
rect 17194 7588 17250 7590
rect 17274 7588 17330 7590
rect 17354 7588 17410 7590
rect 17434 7588 17490 7590
rect 17194 6554 17250 6556
rect 17274 6554 17330 6556
rect 17354 6554 17410 6556
rect 17434 6554 17490 6556
rect 17194 6502 17240 6554
rect 17240 6502 17250 6554
rect 17274 6502 17304 6554
rect 17304 6502 17316 6554
rect 17316 6502 17330 6554
rect 17354 6502 17368 6554
rect 17368 6502 17380 6554
rect 17380 6502 17410 6554
rect 17434 6502 17444 6554
rect 17444 6502 17490 6554
rect 17194 6500 17250 6502
rect 17274 6500 17330 6502
rect 17354 6500 17410 6502
rect 17434 6500 17490 6502
rect 16946 5616 17002 5672
rect 17314 5652 17316 5672
rect 17316 5652 17368 5672
rect 17368 5652 17370 5672
rect 17314 5616 17370 5652
rect 17194 5466 17250 5468
rect 17274 5466 17330 5468
rect 17354 5466 17410 5468
rect 17434 5466 17490 5468
rect 17194 5414 17240 5466
rect 17240 5414 17250 5466
rect 17274 5414 17304 5466
rect 17304 5414 17316 5466
rect 17316 5414 17330 5466
rect 17354 5414 17368 5466
rect 17368 5414 17380 5466
rect 17380 5414 17410 5466
rect 17434 5414 17444 5466
rect 17444 5414 17490 5466
rect 17194 5412 17250 5414
rect 17274 5412 17330 5414
rect 17354 5412 17410 5414
rect 17434 5412 17490 5414
rect 17774 8336 17830 8392
rect 17194 4378 17250 4380
rect 17274 4378 17330 4380
rect 17354 4378 17410 4380
rect 17434 4378 17490 4380
rect 17194 4326 17240 4378
rect 17240 4326 17250 4378
rect 17274 4326 17304 4378
rect 17304 4326 17316 4378
rect 17316 4326 17330 4378
rect 17354 4326 17368 4378
rect 17368 4326 17380 4378
rect 17380 4326 17410 4378
rect 17434 4326 17444 4378
rect 17444 4326 17490 4378
rect 17194 4324 17250 4326
rect 17274 4324 17330 4326
rect 17354 4324 17410 4326
rect 17434 4324 17490 4326
rect 17194 3290 17250 3292
rect 17274 3290 17330 3292
rect 17354 3290 17410 3292
rect 17434 3290 17490 3292
rect 17194 3238 17240 3290
rect 17240 3238 17250 3290
rect 17274 3238 17304 3290
rect 17304 3238 17316 3290
rect 17316 3238 17330 3290
rect 17354 3238 17368 3290
rect 17368 3238 17380 3290
rect 17380 3238 17410 3290
rect 17434 3238 17444 3290
rect 17444 3238 17490 3290
rect 17194 3236 17250 3238
rect 17274 3236 17330 3238
rect 17354 3236 17410 3238
rect 17434 3236 17490 3238
rect 16118 856 16174 912
rect 17194 2202 17250 2204
rect 17274 2202 17330 2204
rect 17354 2202 17410 2204
rect 17434 2202 17490 2204
rect 17194 2150 17240 2202
rect 17240 2150 17250 2202
rect 17274 2150 17304 2202
rect 17304 2150 17316 2202
rect 17316 2150 17330 2202
rect 17354 2150 17368 2202
rect 17368 2150 17380 2202
rect 17380 2150 17410 2202
rect 17434 2150 17444 2202
rect 17444 2150 17490 2202
rect 17194 2148 17250 2150
rect 17274 2148 17330 2150
rect 17354 2148 17410 2150
rect 17434 2148 17490 2150
rect 19338 16632 19394 16688
rect 19890 16632 19946 16688
rect 20552 16890 20608 16892
rect 20632 16890 20688 16892
rect 20712 16890 20768 16892
rect 20792 16890 20848 16892
rect 20552 16838 20598 16890
rect 20598 16838 20608 16890
rect 20632 16838 20662 16890
rect 20662 16838 20674 16890
rect 20674 16838 20688 16890
rect 20712 16838 20726 16890
rect 20726 16838 20738 16890
rect 20738 16838 20768 16890
rect 20792 16838 20802 16890
rect 20802 16838 20848 16890
rect 20552 16836 20608 16838
rect 20632 16836 20688 16838
rect 20712 16836 20768 16838
rect 20792 16836 20848 16838
rect 20552 15802 20608 15804
rect 20632 15802 20688 15804
rect 20712 15802 20768 15804
rect 20792 15802 20848 15804
rect 20552 15750 20598 15802
rect 20598 15750 20608 15802
rect 20632 15750 20662 15802
rect 20662 15750 20674 15802
rect 20674 15750 20688 15802
rect 20712 15750 20726 15802
rect 20726 15750 20738 15802
rect 20738 15750 20768 15802
rect 20792 15750 20802 15802
rect 20802 15750 20848 15802
rect 20552 15748 20608 15750
rect 20632 15748 20688 15750
rect 20712 15748 20768 15750
rect 20792 15748 20848 15750
rect 19338 13776 19394 13832
rect 18786 11736 18842 11792
rect 19338 11636 19340 11656
rect 19340 11636 19392 11656
rect 19392 11636 19394 11656
rect 19338 11600 19394 11636
rect 18878 11056 18934 11112
rect 19246 11056 19302 11112
rect 18418 1944 18474 2000
rect 18970 1420 19026 1456
rect 18970 1400 18972 1420
rect 18972 1400 19024 1420
rect 19024 1400 19026 1420
rect 17194 1114 17250 1116
rect 17274 1114 17330 1116
rect 17354 1114 17410 1116
rect 17434 1114 17490 1116
rect 17194 1062 17240 1114
rect 17240 1062 17250 1114
rect 17274 1062 17304 1114
rect 17304 1062 17316 1114
rect 17316 1062 17330 1114
rect 17354 1062 17368 1114
rect 17368 1062 17380 1114
rect 17380 1062 17410 1114
rect 17434 1062 17444 1114
rect 17444 1062 17490 1114
rect 17194 1060 17250 1062
rect 17274 1060 17330 1062
rect 17354 1060 17410 1062
rect 17434 1060 17490 1062
rect 19890 11636 19892 11656
rect 19892 11636 19944 11656
rect 19944 11636 19946 11656
rect 19890 11600 19946 11636
rect 20552 14714 20608 14716
rect 20632 14714 20688 14716
rect 20712 14714 20768 14716
rect 20792 14714 20848 14716
rect 20552 14662 20598 14714
rect 20598 14662 20608 14714
rect 20632 14662 20662 14714
rect 20662 14662 20674 14714
rect 20674 14662 20688 14714
rect 20712 14662 20726 14714
rect 20726 14662 20738 14714
rect 20738 14662 20768 14714
rect 20792 14662 20802 14714
rect 20802 14662 20848 14714
rect 20552 14660 20608 14662
rect 20632 14660 20688 14662
rect 20712 14660 20768 14662
rect 20792 14660 20848 14662
rect 20718 13812 20720 13832
rect 20720 13812 20772 13832
rect 20772 13812 20774 13832
rect 20718 13776 20774 13812
rect 20552 13626 20608 13628
rect 20632 13626 20688 13628
rect 20712 13626 20768 13628
rect 20792 13626 20848 13628
rect 20552 13574 20598 13626
rect 20598 13574 20608 13626
rect 20632 13574 20662 13626
rect 20662 13574 20674 13626
rect 20674 13574 20688 13626
rect 20712 13574 20726 13626
rect 20726 13574 20738 13626
rect 20738 13574 20768 13626
rect 20792 13574 20802 13626
rect 20802 13574 20848 13626
rect 20552 13572 20608 13574
rect 20632 13572 20688 13574
rect 20712 13572 20768 13574
rect 20792 13572 20848 13574
rect 20552 12538 20608 12540
rect 20632 12538 20688 12540
rect 20712 12538 20768 12540
rect 20792 12538 20848 12540
rect 20552 12486 20598 12538
rect 20598 12486 20608 12538
rect 20632 12486 20662 12538
rect 20662 12486 20674 12538
rect 20674 12486 20688 12538
rect 20712 12486 20726 12538
rect 20726 12486 20738 12538
rect 20738 12486 20768 12538
rect 20792 12486 20802 12538
rect 20802 12486 20848 12538
rect 20552 12484 20608 12486
rect 20632 12484 20688 12486
rect 20712 12484 20768 12486
rect 20792 12484 20848 12486
rect 20552 11450 20608 11452
rect 20632 11450 20688 11452
rect 20712 11450 20768 11452
rect 20792 11450 20848 11452
rect 20552 11398 20598 11450
rect 20598 11398 20608 11450
rect 20632 11398 20662 11450
rect 20662 11398 20674 11450
rect 20674 11398 20688 11450
rect 20712 11398 20726 11450
rect 20726 11398 20738 11450
rect 20738 11398 20768 11450
rect 20792 11398 20802 11450
rect 20802 11398 20848 11450
rect 20552 11396 20608 11398
rect 20632 11396 20688 11398
rect 20712 11396 20768 11398
rect 20792 11396 20848 11398
rect 20552 10362 20608 10364
rect 20632 10362 20688 10364
rect 20712 10362 20768 10364
rect 20792 10362 20848 10364
rect 20552 10310 20598 10362
rect 20598 10310 20608 10362
rect 20632 10310 20662 10362
rect 20662 10310 20674 10362
rect 20674 10310 20688 10362
rect 20712 10310 20726 10362
rect 20726 10310 20738 10362
rect 20738 10310 20768 10362
rect 20792 10310 20802 10362
rect 20802 10310 20848 10362
rect 20552 10308 20608 10310
rect 20632 10308 20688 10310
rect 20712 10308 20768 10310
rect 20792 10308 20848 10310
rect 20552 9274 20608 9276
rect 20632 9274 20688 9276
rect 20712 9274 20768 9276
rect 20792 9274 20848 9276
rect 20552 9222 20598 9274
rect 20598 9222 20608 9274
rect 20632 9222 20662 9274
rect 20662 9222 20674 9274
rect 20674 9222 20688 9274
rect 20712 9222 20726 9274
rect 20726 9222 20738 9274
rect 20738 9222 20768 9274
rect 20792 9222 20802 9274
rect 20802 9222 20848 9274
rect 20552 9220 20608 9222
rect 20632 9220 20688 9222
rect 20712 9220 20768 9222
rect 20792 9220 20848 9222
rect 20552 8186 20608 8188
rect 20632 8186 20688 8188
rect 20712 8186 20768 8188
rect 20792 8186 20848 8188
rect 20552 8134 20598 8186
rect 20598 8134 20608 8186
rect 20632 8134 20662 8186
rect 20662 8134 20674 8186
rect 20674 8134 20688 8186
rect 20712 8134 20726 8186
rect 20726 8134 20738 8186
rect 20738 8134 20768 8186
rect 20792 8134 20802 8186
rect 20802 8134 20848 8186
rect 20552 8132 20608 8134
rect 20632 8132 20688 8134
rect 20712 8132 20768 8134
rect 20792 8132 20848 8134
rect 20552 7098 20608 7100
rect 20632 7098 20688 7100
rect 20712 7098 20768 7100
rect 20792 7098 20848 7100
rect 20552 7046 20598 7098
rect 20598 7046 20608 7098
rect 20632 7046 20662 7098
rect 20662 7046 20674 7098
rect 20674 7046 20688 7098
rect 20712 7046 20726 7098
rect 20726 7046 20738 7098
rect 20738 7046 20768 7098
rect 20792 7046 20802 7098
rect 20802 7046 20848 7098
rect 20552 7044 20608 7046
rect 20632 7044 20688 7046
rect 20712 7044 20768 7046
rect 20792 7044 20848 7046
rect 20552 6010 20608 6012
rect 20632 6010 20688 6012
rect 20712 6010 20768 6012
rect 20792 6010 20848 6012
rect 20552 5958 20598 6010
rect 20598 5958 20608 6010
rect 20632 5958 20662 6010
rect 20662 5958 20674 6010
rect 20674 5958 20688 6010
rect 20712 5958 20726 6010
rect 20726 5958 20738 6010
rect 20738 5958 20768 6010
rect 20792 5958 20802 6010
rect 20802 5958 20848 6010
rect 20552 5956 20608 5958
rect 20632 5956 20688 5958
rect 20712 5956 20768 5958
rect 20792 5956 20848 5958
rect 20552 4922 20608 4924
rect 20632 4922 20688 4924
rect 20712 4922 20768 4924
rect 20792 4922 20848 4924
rect 20552 4870 20598 4922
rect 20598 4870 20608 4922
rect 20632 4870 20662 4922
rect 20662 4870 20674 4922
rect 20674 4870 20688 4922
rect 20712 4870 20726 4922
rect 20726 4870 20738 4922
rect 20738 4870 20768 4922
rect 20792 4870 20802 4922
rect 20802 4870 20848 4922
rect 20552 4868 20608 4870
rect 20632 4868 20688 4870
rect 20712 4868 20768 4870
rect 20792 4868 20848 4870
rect 20552 3834 20608 3836
rect 20632 3834 20688 3836
rect 20712 3834 20768 3836
rect 20792 3834 20848 3836
rect 20552 3782 20598 3834
rect 20598 3782 20608 3834
rect 20632 3782 20662 3834
rect 20662 3782 20674 3834
rect 20674 3782 20688 3834
rect 20712 3782 20726 3834
rect 20726 3782 20738 3834
rect 20738 3782 20768 3834
rect 20792 3782 20802 3834
rect 20802 3782 20848 3834
rect 20552 3780 20608 3782
rect 20632 3780 20688 3782
rect 20712 3780 20768 3782
rect 20792 3780 20848 3782
rect 20552 2746 20608 2748
rect 20632 2746 20688 2748
rect 20712 2746 20768 2748
rect 20792 2746 20848 2748
rect 20552 2694 20598 2746
rect 20598 2694 20608 2746
rect 20632 2694 20662 2746
rect 20662 2694 20674 2746
rect 20674 2694 20688 2746
rect 20712 2694 20726 2746
rect 20726 2694 20738 2746
rect 20738 2694 20768 2746
rect 20792 2694 20802 2746
rect 20802 2694 20848 2746
rect 20552 2692 20608 2694
rect 20632 2692 20688 2694
rect 20712 2692 20768 2694
rect 20792 2692 20848 2694
rect 20258 1964 20314 2000
rect 20258 1944 20260 1964
rect 20260 1944 20312 1964
rect 20312 1944 20314 1964
rect 20552 1658 20608 1660
rect 20632 1658 20688 1660
rect 20712 1658 20768 1660
rect 20792 1658 20848 1660
rect 20552 1606 20598 1658
rect 20598 1606 20608 1658
rect 20632 1606 20662 1658
rect 20662 1606 20674 1658
rect 20674 1606 20688 1658
rect 20712 1606 20726 1658
rect 20726 1606 20738 1658
rect 20738 1606 20768 1658
rect 20792 1606 20802 1658
rect 20802 1606 20848 1658
rect 20552 1604 20608 1606
rect 20632 1604 20688 1606
rect 20712 1604 20768 1606
rect 20792 1604 20848 1606
rect 21730 13812 21732 13832
rect 21732 13812 21784 13832
rect 21784 13812 21786 13832
rect 21730 13776 21786 13812
rect 21638 12552 21694 12608
rect 22006 10124 22062 10160
rect 22006 10104 22008 10124
rect 22008 10104 22060 10124
rect 22060 10104 22062 10124
rect 23910 16346 23966 16348
rect 23990 16346 24046 16348
rect 24070 16346 24126 16348
rect 24150 16346 24206 16348
rect 23910 16294 23956 16346
rect 23956 16294 23966 16346
rect 23990 16294 24020 16346
rect 24020 16294 24032 16346
rect 24032 16294 24046 16346
rect 24070 16294 24084 16346
rect 24084 16294 24096 16346
rect 24096 16294 24126 16346
rect 24150 16294 24160 16346
rect 24160 16294 24206 16346
rect 23910 16292 23966 16294
rect 23990 16292 24046 16294
rect 24070 16292 24126 16294
rect 24150 16292 24206 16294
rect 23910 15258 23966 15260
rect 23990 15258 24046 15260
rect 24070 15258 24126 15260
rect 24150 15258 24206 15260
rect 23910 15206 23956 15258
rect 23956 15206 23966 15258
rect 23990 15206 24020 15258
rect 24020 15206 24032 15258
rect 24032 15206 24046 15258
rect 24070 15206 24084 15258
rect 24084 15206 24096 15258
rect 24096 15206 24126 15258
rect 24150 15206 24160 15258
rect 24160 15206 24206 15258
rect 23910 15204 23966 15206
rect 23990 15204 24046 15206
rect 24070 15204 24126 15206
rect 24150 15204 24206 15206
rect 23910 14170 23966 14172
rect 23990 14170 24046 14172
rect 24070 14170 24126 14172
rect 24150 14170 24206 14172
rect 23910 14118 23956 14170
rect 23956 14118 23966 14170
rect 23990 14118 24020 14170
rect 24020 14118 24032 14170
rect 24032 14118 24046 14170
rect 24070 14118 24084 14170
rect 24084 14118 24096 14170
rect 24096 14118 24126 14170
rect 24150 14118 24160 14170
rect 24160 14118 24206 14170
rect 23910 14116 23966 14118
rect 23990 14116 24046 14118
rect 24070 14116 24126 14118
rect 24150 14116 24206 14118
rect 23570 13776 23626 13832
rect 24306 13776 24362 13832
rect 23910 13082 23966 13084
rect 23990 13082 24046 13084
rect 24070 13082 24126 13084
rect 24150 13082 24206 13084
rect 23910 13030 23956 13082
rect 23956 13030 23966 13082
rect 23990 13030 24020 13082
rect 24020 13030 24032 13082
rect 24032 13030 24046 13082
rect 24070 13030 24084 13082
rect 24084 13030 24096 13082
rect 24096 13030 24126 13082
rect 24150 13030 24160 13082
rect 24160 13030 24206 13082
rect 23910 13028 23966 13030
rect 23990 13028 24046 13030
rect 24070 13028 24126 13030
rect 24150 13028 24206 13030
rect 23910 11994 23966 11996
rect 23990 11994 24046 11996
rect 24070 11994 24126 11996
rect 24150 11994 24206 11996
rect 23910 11942 23956 11994
rect 23956 11942 23966 11994
rect 23990 11942 24020 11994
rect 24020 11942 24032 11994
rect 24032 11942 24046 11994
rect 24070 11942 24084 11994
rect 24084 11942 24096 11994
rect 24096 11942 24126 11994
rect 24150 11942 24160 11994
rect 24160 11942 24206 11994
rect 23910 11940 23966 11942
rect 23990 11940 24046 11942
rect 24070 11940 24126 11942
rect 24150 11940 24206 11942
rect 23386 10124 23442 10160
rect 23386 10104 23388 10124
rect 23388 10104 23440 10124
rect 23440 10104 23442 10124
rect 23910 10906 23966 10908
rect 23990 10906 24046 10908
rect 24070 10906 24126 10908
rect 24150 10906 24206 10908
rect 23910 10854 23956 10906
rect 23956 10854 23966 10906
rect 23990 10854 24020 10906
rect 24020 10854 24032 10906
rect 24032 10854 24046 10906
rect 24070 10854 24084 10906
rect 24084 10854 24096 10906
rect 24096 10854 24126 10906
rect 24150 10854 24160 10906
rect 24160 10854 24206 10906
rect 23910 10852 23966 10854
rect 23990 10852 24046 10854
rect 24070 10852 24126 10854
rect 24150 10852 24206 10854
rect 24398 9968 24454 10024
rect 23910 9818 23966 9820
rect 23990 9818 24046 9820
rect 24070 9818 24126 9820
rect 24150 9818 24206 9820
rect 23910 9766 23956 9818
rect 23956 9766 23966 9818
rect 23990 9766 24020 9818
rect 24020 9766 24032 9818
rect 24032 9766 24046 9818
rect 24070 9766 24084 9818
rect 24084 9766 24096 9818
rect 24096 9766 24126 9818
rect 24150 9766 24160 9818
rect 24160 9766 24206 9818
rect 23910 9764 23966 9766
rect 23990 9764 24046 9766
rect 24070 9764 24126 9766
rect 24150 9764 24206 9766
rect 21730 7384 21786 7440
rect 20552 570 20608 572
rect 20632 570 20688 572
rect 20712 570 20768 572
rect 20792 570 20848 572
rect 20552 518 20598 570
rect 20598 518 20608 570
rect 20632 518 20662 570
rect 20662 518 20674 570
rect 20674 518 20688 570
rect 20712 518 20726 570
rect 20726 518 20738 570
rect 20738 518 20768 570
rect 20792 518 20802 570
rect 20802 518 20848 570
rect 20552 516 20608 518
rect 20632 516 20688 518
rect 20712 516 20768 518
rect 20792 516 20848 518
rect 22006 1420 22062 1456
rect 23910 8730 23966 8732
rect 23990 8730 24046 8732
rect 24070 8730 24126 8732
rect 24150 8730 24206 8732
rect 23910 8678 23956 8730
rect 23956 8678 23966 8730
rect 23990 8678 24020 8730
rect 24020 8678 24032 8730
rect 24032 8678 24046 8730
rect 24070 8678 24084 8730
rect 24084 8678 24096 8730
rect 24096 8678 24126 8730
rect 24150 8678 24160 8730
rect 24160 8678 24206 8730
rect 23910 8676 23966 8678
rect 23990 8676 24046 8678
rect 24070 8676 24126 8678
rect 24150 8676 24206 8678
rect 23910 7642 23966 7644
rect 23990 7642 24046 7644
rect 24070 7642 24126 7644
rect 24150 7642 24206 7644
rect 23910 7590 23956 7642
rect 23956 7590 23966 7642
rect 23990 7590 24020 7642
rect 24020 7590 24032 7642
rect 24032 7590 24046 7642
rect 24070 7590 24084 7642
rect 24084 7590 24096 7642
rect 24096 7590 24126 7642
rect 24150 7590 24160 7642
rect 24160 7590 24206 7642
rect 23910 7588 23966 7590
rect 23990 7588 24046 7590
rect 24070 7588 24126 7590
rect 24150 7588 24206 7590
rect 23910 6554 23966 6556
rect 23990 6554 24046 6556
rect 24070 6554 24126 6556
rect 24150 6554 24206 6556
rect 23910 6502 23956 6554
rect 23956 6502 23966 6554
rect 23990 6502 24020 6554
rect 24020 6502 24032 6554
rect 24032 6502 24046 6554
rect 24070 6502 24084 6554
rect 24084 6502 24096 6554
rect 24096 6502 24126 6554
rect 24150 6502 24160 6554
rect 24160 6502 24206 6554
rect 23910 6500 23966 6502
rect 23990 6500 24046 6502
rect 24070 6500 24126 6502
rect 24150 6500 24206 6502
rect 25502 12280 25558 12336
rect 26054 13812 26056 13832
rect 26056 13812 26108 13832
rect 26108 13812 26110 13832
rect 26054 13776 26110 13812
rect 26238 13776 26294 13832
rect 26146 12280 26202 12336
rect 26790 13912 26846 13968
rect 27268 16890 27324 16892
rect 27348 16890 27404 16892
rect 27428 16890 27484 16892
rect 27508 16890 27564 16892
rect 27268 16838 27314 16890
rect 27314 16838 27324 16890
rect 27348 16838 27378 16890
rect 27378 16838 27390 16890
rect 27390 16838 27404 16890
rect 27428 16838 27442 16890
rect 27442 16838 27454 16890
rect 27454 16838 27484 16890
rect 27508 16838 27518 16890
rect 27518 16838 27564 16890
rect 27268 16836 27324 16838
rect 27348 16836 27404 16838
rect 27428 16836 27484 16838
rect 27508 16836 27564 16838
rect 27268 15802 27324 15804
rect 27348 15802 27404 15804
rect 27428 15802 27484 15804
rect 27508 15802 27564 15804
rect 27268 15750 27314 15802
rect 27314 15750 27324 15802
rect 27348 15750 27378 15802
rect 27378 15750 27390 15802
rect 27390 15750 27404 15802
rect 27428 15750 27442 15802
rect 27442 15750 27454 15802
rect 27454 15750 27484 15802
rect 27508 15750 27518 15802
rect 27518 15750 27564 15802
rect 27268 15748 27324 15750
rect 27348 15748 27404 15750
rect 27428 15748 27484 15750
rect 27508 15748 27564 15750
rect 27268 14714 27324 14716
rect 27348 14714 27404 14716
rect 27428 14714 27484 14716
rect 27508 14714 27564 14716
rect 27268 14662 27314 14714
rect 27314 14662 27324 14714
rect 27348 14662 27378 14714
rect 27378 14662 27390 14714
rect 27390 14662 27404 14714
rect 27428 14662 27442 14714
rect 27442 14662 27454 14714
rect 27454 14662 27484 14714
rect 27508 14662 27518 14714
rect 27518 14662 27564 14714
rect 27268 14660 27324 14662
rect 27348 14660 27404 14662
rect 27428 14660 27484 14662
rect 27508 14660 27564 14662
rect 27158 13776 27214 13832
rect 27268 13626 27324 13628
rect 27348 13626 27404 13628
rect 27428 13626 27484 13628
rect 27508 13626 27564 13628
rect 27268 13574 27314 13626
rect 27314 13574 27324 13626
rect 27348 13574 27378 13626
rect 27378 13574 27390 13626
rect 27390 13574 27404 13626
rect 27428 13574 27442 13626
rect 27442 13574 27454 13626
rect 27454 13574 27484 13626
rect 27508 13574 27518 13626
rect 27518 13574 27564 13626
rect 27268 13572 27324 13574
rect 27348 13572 27404 13574
rect 27428 13572 27484 13574
rect 27508 13572 27564 13574
rect 27268 12538 27324 12540
rect 27348 12538 27404 12540
rect 27428 12538 27484 12540
rect 27508 12538 27564 12540
rect 27268 12486 27314 12538
rect 27314 12486 27324 12538
rect 27348 12486 27378 12538
rect 27378 12486 27390 12538
rect 27390 12486 27404 12538
rect 27428 12486 27442 12538
rect 27442 12486 27454 12538
rect 27454 12486 27484 12538
rect 27508 12486 27518 12538
rect 27518 12486 27564 12538
rect 27268 12484 27324 12486
rect 27348 12484 27404 12486
rect 27428 12484 27484 12486
rect 27508 12484 27564 12486
rect 27268 11450 27324 11452
rect 27348 11450 27404 11452
rect 27428 11450 27484 11452
rect 27508 11450 27564 11452
rect 27268 11398 27314 11450
rect 27314 11398 27324 11450
rect 27348 11398 27378 11450
rect 27378 11398 27390 11450
rect 27390 11398 27404 11450
rect 27428 11398 27442 11450
rect 27442 11398 27454 11450
rect 27454 11398 27484 11450
rect 27508 11398 27518 11450
rect 27518 11398 27564 11450
rect 27268 11396 27324 11398
rect 27348 11396 27404 11398
rect 27428 11396 27484 11398
rect 27508 11396 27564 11398
rect 27268 10362 27324 10364
rect 27348 10362 27404 10364
rect 27428 10362 27484 10364
rect 27508 10362 27564 10364
rect 27268 10310 27314 10362
rect 27314 10310 27324 10362
rect 27348 10310 27378 10362
rect 27378 10310 27390 10362
rect 27390 10310 27404 10362
rect 27428 10310 27442 10362
rect 27442 10310 27454 10362
rect 27454 10310 27484 10362
rect 27508 10310 27518 10362
rect 27518 10310 27564 10362
rect 27268 10308 27324 10310
rect 27348 10308 27404 10310
rect 27428 10308 27484 10310
rect 27508 10308 27564 10310
rect 23910 5466 23966 5468
rect 23990 5466 24046 5468
rect 24070 5466 24126 5468
rect 24150 5466 24206 5468
rect 23910 5414 23956 5466
rect 23956 5414 23966 5466
rect 23990 5414 24020 5466
rect 24020 5414 24032 5466
rect 24032 5414 24046 5466
rect 24070 5414 24084 5466
rect 24084 5414 24096 5466
rect 24096 5414 24126 5466
rect 24150 5414 24160 5466
rect 24160 5414 24206 5466
rect 23910 5412 23966 5414
rect 23990 5412 24046 5414
rect 24070 5412 24126 5414
rect 24150 5412 24206 5414
rect 26422 9988 26478 10024
rect 26422 9968 26424 9988
rect 26424 9968 26476 9988
rect 26476 9968 26478 9988
rect 27268 9274 27324 9276
rect 27348 9274 27404 9276
rect 27428 9274 27484 9276
rect 27508 9274 27564 9276
rect 27268 9222 27314 9274
rect 27314 9222 27324 9274
rect 27348 9222 27378 9274
rect 27378 9222 27390 9274
rect 27390 9222 27404 9274
rect 27428 9222 27442 9274
rect 27442 9222 27454 9274
rect 27454 9222 27484 9274
rect 27508 9222 27518 9274
rect 27518 9222 27564 9274
rect 27268 9220 27324 9222
rect 27348 9220 27404 9222
rect 27428 9220 27484 9222
rect 27508 9220 27564 9222
rect 27268 8186 27324 8188
rect 27348 8186 27404 8188
rect 27428 8186 27484 8188
rect 27508 8186 27564 8188
rect 27268 8134 27314 8186
rect 27314 8134 27324 8186
rect 27348 8134 27378 8186
rect 27378 8134 27390 8186
rect 27390 8134 27404 8186
rect 27428 8134 27442 8186
rect 27442 8134 27454 8186
rect 27454 8134 27484 8186
rect 27508 8134 27518 8186
rect 27518 8134 27564 8186
rect 27268 8132 27324 8134
rect 27348 8132 27404 8134
rect 27428 8132 27484 8134
rect 27508 8132 27564 8134
rect 27268 7098 27324 7100
rect 27348 7098 27404 7100
rect 27428 7098 27484 7100
rect 27508 7098 27564 7100
rect 27268 7046 27314 7098
rect 27314 7046 27324 7098
rect 27348 7046 27378 7098
rect 27378 7046 27390 7098
rect 27390 7046 27404 7098
rect 27428 7046 27442 7098
rect 27442 7046 27454 7098
rect 27454 7046 27484 7098
rect 27508 7046 27518 7098
rect 27518 7046 27564 7098
rect 27268 7044 27324 7046
rect 27348 7044 27404 7046
rect 27428 7044 27484 7046
rect 27508 7044 27564 7046
rect 27268 6010 27324 6012
rect 27348 6010 27404 6012
rect 27428 6010 27484 6012
rect 27508 6010 27564 6012
rect 27268 5958 27314 6010
rect 27314 5958 27324 6010
rect 27348 5958 27378 6010
rect 27378 5958 27390 6010
rect 27390 5958 27404 6010
rect 27428 5958 27442 6010
rect 27442 5958 27454 6010
rect 27454 5958 27484 6010
rect 27508 5958 27518 6010
rect 27518 5958 27564 6010
rect 27268 5956 27324 5958
rect 27348 5956 27404 5958
rect 27428 5956 27484 5958
rect 27508 5956 27564 5958
rect 27268 4922 27324 4924
rect 27348 4922 27404 4924
rect 27428 4922 27484 4924
rect 27508 4922 27564 4924
rect 27268 4870 27314 4922
rect 27314 4870 27324 4922
rect 27348 4870 27378 4922
rect 27378 4870 27390 4922
rect 27390 4870 27404 4922
rect 27428 4870 27442 4922
rect 27442 4870 27454 4922
rect 27454 4870 27484 4922
rect 27508 4870 27518 4922
rect 27518 4870 27564 4922
rect 27268 4868 27324 4870
rect 27348 4868 27404 4870
rect 27428 4868 27484 4870
rect 27508 4868 27564 4870
rect 23910 4378 23966 4380
rect 23990 4378 24046 4380
rect 24070 4378 24126 4380
rect 24150 4378 24206 4380
rect 23910 4326 23956 4378
rect 23956 4326 23966 4378
rect 23990 4326 24020 4378
rect 24020 4326 24032 4378
rect 24032 4326 24046 4378
rect 24070 4326 24084 4378
rect 24084 4326 24096 4378
rect 24096 4326 24126 4378
rect 24150 4326 24160 4378
rect 24160 4326 24206 4378
rect 23910 4324 23966 4326
rect 23990 4324 24046 4326
rect 24070 4324 24126 4326
rect 24150 4324 24206 4326
rect 27268 3834 27324 3836
rect 27348 3834 27404 3836
rect 27428 3834 27484 3836
rect 27508 3834 27564 3836
rect 27268 3782 27314 3834
rect 27314 3782 27324 3834
rect 27348 3782 27378 3834
rect 27378 3782 27390 3834
rect 27390 3782 27404 3834
rect 27428 3782 27442 3834
rect 27442 3782 27454 3834
rect 27454 3782 27484 3834
rect 27508 3782 27518 3834
rect 27518 3782 27564 3834
rect 27268 3780 27324 3782
rect 27348 3780 27404 3782
rect 27428 3780 27484 3782
rect 27508 3780 27564 3782
rect 23910 3290 23966 3292
rect 23990 3290 24046 3292
rect 24070 3290 24126 3292
rect 24150 3290 24206 3292
rect 23910 3238 23956 3290
rect 23956 3238 23966 3290
rect 23990 3238 24020 3290
rect 24020 3238 24032 3290
rect 24032 3238 24046 3290
rect 24070 3238 24084 3290
rect 24084 3238 24096 3290
rect 24096 3238 24126 3290
rect 24150 3238 24160 3290
rect 24160 3238 24206 3290
rect 23910 3236 23966 3238
rect 23990 3236 24046 3238
rect 24070 3236 24126 3238
rect 24150 3236 24206 3238
rect 27268 2746 27324 2748
rect 27348 2746 27404 2748
rect 27428 2746 27484 2748
rect 27508 2746 27564 2748
rect 27268 2694 27314 2746
rect 27314 2694 27324 2746
rect 27348 2694 27378 2746
rect 27378 2694 27390 2746
rect 27390 2694 27404 2746
rect 27428 2694 27442 2746
rect 27442 2694 27454 2746
rect 27454 2694 27484 2746
rect 27508 2694 27518 2746
rect 27518 2694 27564 2746
rect 27268 2692 27324 2694
rect 27348 2692 27404 2694
rect 27428 2692 27484 2694
rect 27508 2692 27564 2694
rect 23910 2202 23966 2204
rect 23990 2202 24046 2204
rect 24070 2202 24126 2204
rect 24150 2202 24206 2204
rect 23910 2150 23956 2202
rect 23956 2150 23966 2202
rect 23990 2150 24020 2202
rect 24020 2150 24032 2202
rect 24032 2150 24046 2202
rect 24070 2150 24084 2202
rect 24084 2150 24096 2202
rect 24096 2150 24126 2202
rect 24150 2150 24160 2202
rect 24160 2150 24206 2202
rect 23910 2148 23966 2150
rect 23990 2148 24046 2150
rect 24070 2148 24126 2150
rect 24150 2148 24206 2150
rect 22006 1400 22008 1420
rect 22008 1400 22060 1420
rect 22060 1400 22062 1420
rect 27268 1658 27324 1660
rect 27348 1658 27404 1660
rect 27428 1658 27484 1660
rect 27508 1658 27564 1660
rect 27268 1606 27314 1658
rect 27314 1606 27324 1658
rect 27348 1606 27378 1658
rect 27378 1606 27390 1658
rect 27390 1606 27404 1658
rect 27428 1606 27442 1658
rect 27442 1606 27454 1658
rect 27454 1606 27484 1658
rect 27508 1606 27518 1658
rect 27518 1606 27564 1658
rect 27268 1604 27324 1606
rect 27348 1604 27404 1606
rect 27428 1604 27484 1606
rect 27508 1604 27564 1606
rect 23910 1114 23966 1116
rect 23990 1114 24046 1116
rect 24070 1114 24126 1116
rect 24150 1114 24206 1116
rect 23910 1062 23956 1114
rect 23956 1062 23966 1114
rect 23990 1062 24020 1114
rect 24020 1062 24032 1114
rect 24032 1062 24046 1114
rect 24070 1062 24084 1114
rect 24084 1062 24096 1114
rect 24096 1062 24126 1114
rect 24150 1062 24160 1114
rect 24160 1062 24206 1114
rect 23910 1060 23966 1062
rect 23990 1060 24046 1062
rect 24070 1060 24126 1062
rect 24150 1060 24206 1062
rect 27268 570 27324 572
rect 27348 570 27404 572
rect 27428 570 27484 572
rect 27508 570 27564 572
rect 27268 518 27314 570
rect 27314 518 27324 570
rect 27348 518 27378 570
rect 27378 518 27390 570
rect 27390 518 27404 570
rect 27428 518 27442 570
rect 27442 518 27454 570
rect 27454 518 27484 570
rect 27508 518 27518 570
rect 27518 518 27564 570
rect 27268 516 27324 518
rect 27348 516 27404 518
rect 27428 516 27484 518
rect 27508 516 27564 518
<< metal3 >>
rect 3752 17440 4068 17441
rect 3752 17376 3758 17440
rect 3822 17376 3838 17440
rect 3902 17376 3918 17440
rect 3982 17376 3998 17440
rect 4062 17376 4068 17440
rect 3752 17375 4068 17376
rect 10468 17440 10784 17441
rect 10468 17376 10474 17440
rect 10538 17376 10554 17440
rect 10618 17376 10634 17440
rect 10698 17376 10714 17440
rect 10778 17376 10784 17440
rect 10468 17375 10784 17376
rect 17184 17440 17500 17441
rect 17184 17376 17190 17440
rect 17254 17376 17270 17440
rect 17334 17376 17350 17440
rect 17414 17376 17430 17440
rect 17494 17376 17500 17440
rect 17184 17375 17500 17376
rect 23900 17440 24216 17441
rect 23900 17376 23906 17440
rect 23970 17376 23986 17440
rect 24050 17376 24066 17440
rect 24130 17376 24146 17440
rect 24210 17376 24216 17440
rect 23900 17375 24216 17376
rect 19517 17234 19583 17237
rect 24025 17234 24091 17237
rect 19517 17232 24091 17234
rect 19517 17176 19522 17232
rect 19578 17176 24030 17232
rect 24086 17176 24091 17232
rect 19517 17174 24091 17176
rect 19517 17171 19583 17174
rect 24025 17171 24091 17174
rect 7110 16896 7426 16897
rect 7110 16832 7116 16896
rect 7180 16832 7196 16896
rect 7260 16832 7276 16896
rect 7340 16832 7356 16896
rect 7420 16832 7426 16896
rect 7110 16831 7426 16832
rect 13826 16896 14142 16897
rect 13826 16832 13832 16896
rect 13896 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14142 16896
rect 13826 16831 14142 16832
rect 20542 16896 20858 16897
rect 20542 16832 20548 16896
rect 20612 16832 20628 16896
rect 20692 16832 20708 16896
rect 20772 16832 20788 16896
rect 20852 16832 20858 16896
rect 20542 16831 20858 16832
rect 27258 16896 27574 16897
rect 27258 16832 27264 16896
rect 27328 16832 27344 16896
rect 27408 16832 27424 16896
rect 27488 16832 27504 16896
rect 27568 16832 27574 16896
rect 27258 16831 27574 16832
rect 13997 16690 14063 16693
rect 19333 16692 19399 16693
rect 14406 16690 14412 16692
rect 13997 16688 14412 16690
rect 13997 16632 14002 16688
rect 14058 16632 14412 16688
rect 13997 16630 14412 16632
rect 13997 16627 14063 16630
rect 14406 16628 14412 16630
rect 14476 16628 14482 16692
rect 19333 16688 19380 16692
rect 19444 16690 19450 16692
rect 19885 16690 19951 16693
rect 20294 16690 20300 16692
rect 19333 16632 19338 16688
rect 19333 16628 19380 16632
rect 19444 16630 19490 16690
rect 19885 16688 20300 16690
rect 19885 16632 19890 16688
rect 19946 16632 20300 16688
rect 19885 16630 20300 16632
rect 19444 16628 19450 16630
rect 19333 16627 19399 16628
rect 19885 16627 19951 16630
rect 20294 16628 20300 16630
rect 20364 16628 20370 16692
rect 3752 16352 4068 16353
rect 3752 16288 3758 16352
rect 3822 16288 3838 16352
rect 3902 16288 3918 16352
rect 3982 16288 3998 16352
rect 4062 16288 4068 16352
rect 3752 16287 4068 16288
rect 10468 16352 10784 16353
rect 10468 16288 10474 16352
rect 10538 16288 10554 16352
rect 10618 16288 10634 16352
rect 10698 16288 10714 16352
rect 10778 16288 10784 16352
rect 10468 16287 10784 16288
rect 17184 16352 17500 16353
rect 17184 16288 17190 16352
rect 17254 16288 17270 16352
rect 17334 16288 17350 16352
rect 17414 16288 17430 16352
rect 17494 16288 17500 16352
rect 17184 16287 17500 16288
rect 23900 16352 24216 16353
rect 23900 16288 23906 16352
rect 23970 16288 23986 16352
rect 24050 16288 24066 16352
rect 24130 16288 24146 16352
rect 24210 16288 24216 16352
rect 23900 16287 24216 16288
rect 7110 15808 7426 15809
rect 7110 15744 7116 15808
rect 7180 15744 7196 15808
rect 7260 15744 7276 15808
rect 7340 15744 7356 15808
rect 7420 15744 7426 15808
rect 7110 15743 7426 15744
rect 13826 15808 14142 15809
rect 13826 15744 13832 15808
rect 13896 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14142 15808
rect 13826 15743 14142 15744
rect 20542 15808 20858 15809
rect 20542 15744 20548 15808
rect 20612 15744 20628 15808
rect 20692 15744 20708 15808
rect 20772 15744 20788 15808
rect 20852 15744 20858 15808
rect 20542 15743 20858 15744
rect 27258 15808 27574 15809
rect 27258 15744 27264 15808
rect 27328 15744 27344 15808
rect 27408 15744 27424 15808
rect 27488 15744 27504 15808
rect 27568 15744 27574 15808
rect 27258 15743 27574 15744
rect 10174 15268 10180 15332
rect 10244 15330 10250 15332
rect 10317 15330 10383 15333
rect 10244 15328 10383 15330
rect 10244 15272 10322 15328
rect 10378 15272 10383 15328
rect 10244 15270 10383 15272
rect 10244 15268 10250 15270
rect 10317 15267 10383 15270
rect 3752 15264 4068 15265
rect 3752 15200 3758 15264
rect 3822 15200 3838 15264
rect 3902 15200 3918 15264
rect 3982 15200 3998 15264
rect 4062 15200 4068 15264
rect 3752 15199 4068 15200
rect 10468 15264 10784 15265
rect 10468 15200 10474 15264
rect 10538 15200 10554 15264
rect 10618 15200 10634 15264
rect 10698 15200 10714 15264
rect 10778 15200 10784 15264
rect 10468 15199 10784 15200
rect 17184 15264 17500 15265
rect 17184 15200 17190 15264
rect 17254 15200 17270 15264
rect 17334 15200 17350 15264
rect 17414 15200 17430 15264
rect 17494 15200 17500 15264
rect 17184 15199 17500 15200
rect 23900 15264 24216 15265
rect 23900 15200 23906 15264
rect 23970 15200 23986 15264
rect 24050 15200 24066 15264
rect 24130 15200 24146 15264
rect 24210 15200 24216 15264
rect 23900 15199 24216 15200
rect 7925 15058 7991 15061
rect 12709 15058 12775 15061
rect 7925 15056 12775 15058
rect 7925 15000 7930 15056
rect 7986 15000 12714 15056
rect 12770 15000 12775 15056
rect 7925 14998 12775 15000
rect 7925 14995 7991 14998
rect 12709 14995 12775 14998
rect 7110 14720 7426 14721
rect 7110 14656 7116 14720
rect 7180 14656 7196 14720
rect 7260 14656 7276 14720
rect 7340 14656 7356 14720
rect 7420 14656 7426 14720
rect 7110 14655 7426 14656
rect 13826 14720 14142 14721
rect 13826 14656 13832 14720
rect 13896 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14142 14720
rect 13826 14655 14142 14656
rect 20542 14720 20858 14721
rect 20542 14656 20548 14720
rect 20612 14656 20628 14720
rect 20692 14656 20708 14720
rect 20772 14656 20788 14720
rect 20852 14656 20858 14720
rect 20542 14655 20858 14656
rect 27258 14720 27574 14721
rect 27258 14656 27264 14720
rect 27328 14656 27344 14720
rect 27408 14656 27424 14720
rect 27488 14656 27504 14720
rect 27568 14656 27574 14720
rect 27258 14655 27574 14656
rect 9857 14514 9923 14517
rect 13997 14514 14063 14517
rect 14825 14514 14891 14517
rect 9857 14512 14891 14514
rect 9857 14456 9862 14512
rect 9918 14456 14002 14512
rect 14058 14456 14830 14512
rect 14886 14456 14891 14512
rect 9857 14454 14891 14456
rect 9857 14451 9923 14454
rect 13997 14451 14063 14454
rect 14825 14451 14891 14454
rect 3752 14176 4068 14177
rect 3752 14112 3758 14176
rect 3822 14112 3838 14176
rect 3902 14112 3918 14176
rect 3982 14112 3998 14176
rect 4062 14112 4068 14176
rect 3752 14111 4068 14112
rect 10468 14176 10784 14177
rect 10468 14112 10474 14176
rect 10538 14112 10554 14176
rect 10618 14112 10634 14176
rect 10698 14112 10714 14176
rect 10778 14112 10784 14176
rect 10468 14111 10784 14112
rect 17184 14176 17500 14177
rect 17184 14112 17190 14176
rect 17254 14112 17270 14176
rect 17334 14112 17350 14176
rect 17414 14112 17430 14176
rect 17494 14112 17500 14176
rect 17184 14111 17500 14112
rect 23900 14176 24216 14177
rect 23900 14112 23906 14176
rect 23970 14112 23986 14176
rect 24050 14112 24066 14176
rect 24130 14112 24146 14176
rect 24210 14112 24216 14176
rect 23900 14111 24216 14112
rect 6177 13970 6243 13973
rect 8201 13970 8267 13973
rect 26785 13970 26851 13973
rect 6177 13968 8267 13970
rect 6177 13912 6182 13968
rect 6238 13912 8206 13968
rect 8262 13912 8267 13968
rect 6177 13910 8267 13912
rect 6177 13907 6243 13910
rect 8201 13907 8267 13910
rect 26006 13968 26851 13970
rect 26006 13912 26790 13968
rect 26846 13912 26851 13968
rect 26006 13910 26851 13912
rect 26006 13837 26066 13910
rect 26785 13907 26851 13910
rect 19333 13834 19399 13837
rect 20713 13834 20779 13837
rect 21725 13834 21791 13837
rect 23565 13834 23631 13837
rect 19333 13832 23631 13834
rect 19333 13776 19338 13832
rect 19394 13776 20718 13832
rect 20774 13776 21730 13832
rect 21786 13776 23570 13832
rect 23626 13776 23631 13832
rect 19333 13774 23631 13776
rect 19333 13771 19399 13774
rect 20713 13771 20779 13774
rect 21725 13771 21791 13774
rect 23565 13771 23631 13774
rect 24301 13834 24367 13837
rect 26006 13834 26115 13837
rect 24301 13832 26115 13834
rect 24301 13776 24306 13832
rect 24362 13776 26054 13832
rect 26110 13776 26115 13832
rect 24301 13774 26115 13776
rect 24301 13771 24367 13774
rect 26049 13771 26115 13774
rect 26233 13834 26299 13837
rect 27153 13834 27219 13837
rect 26233 13832 27219 13834
rect 26233 13776 26238 13832
rect 26294 13776 27158 13832
rect 27214 13776 27219 13832
rect 26233 13774 27219 13776
rect 26233 13771 26299 13774
rect 27153 13771 27219 13774
rect 7110 13632 7426 13633
rect 7110 13568 7116 13632
rect 7180 13568 7196 13632
rect 7260 13568 7276 13632
rect 7340 13568 7356 13632
rect 7420 13568 7426 13632
rect 7110 13567 7426 13568
rect 13826 13632 14142 13633
rect 13826 13568 13832 13632
rect 13896 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14142 13632
rect 13826 13567 14142 13568
rect 20542 13632 20858 13633
rect 20542 13568 20548 13632
rect 20612 13568 20628 13632
rect 20692 13568 20708 13632
rect 20772 13568 20788 13632
rect 20852 13568 20858 13632
rect 20542 13567 20858 13568
rect 27258 13632 27574 13633
rect 27258 13568 27264 13632
rect 27328 13568 27344 13632
rect 27408 13568 27424 13632
rect 27488 13568 27504 13632
rect 27568 13568 27574 13632
rect 27258 13567 27574 13568
rect 15009 13426 15075 13429
rect 16205 13426 16271 13429
rect 15009 13424 16271 13426
rect 15009 13368 15014 13424
rect 15070 13368 16210 13424
rect 16266 13368 16271 13424
rect 15009 13366 16271 13368
rect 15009 13363 15075 13366
rect 16205 13363 16271 13366
rect 13353 13154 13419 13157
rect 15469 13154 15535 13157
rect 13353 13152 15535 13154
rect 13353 13096 13358 13152
rect 13414 13096 15474 13152
rect 15530 13096 15535 13152
rect 13353 13094 15535 13096
rect 13353 13091 13419 13094
rect 15469 13091 15535 13094
rect 3752 13088 4068 13089
rect 3752 13024 3758 13088
rect 3822 13024 3838 13088
rect 3902 13024 3918 13088
rect 3982 13024 3998 13088
rect 4062 13024 4068 13088
rect 3752 13023 4068 13024
rect 10468 13088 10784 13089
rect 10468 13024 10474 13088
rect 10538 13024 10554 13088
rect 10618 13024 10634 13088
rect 10698 13024 10714 13088
rect 10778 13024 10784 13088
rect 10468 13023 10784 13024
rect 17184 13088 17500 13089
rect 17184 13024 17190 13088
rect 17254 13024 17270 13088
rect 17334 13024 17350 13088
rect 17414 13024 17430 13088
rect 17494 13024 17500 13088
rect 17184 13023 17500 13024
rect 23900 13088 24216 13089
rect 23900 13024 23906 13088
rect 23970 13024 23986 13088
rect 24050 13024 24066 13088
rect 24130 13024 24146 13088
rect 24210 13024 24216 13088
rect 23900 13023 24216 13024
rect 3417 12882 3483 12885
rect 4705 12882 4771 12885
rect 3417 12880 4771 12882
rect 3417 12824 3422 12880
rect 3478 12824 4710 12880
rect 4766 12824 4771 12880
rect 3417 12822 4771 12824
rect 3417 12819 3483 12822
rect 4705 12819 4771 12822
rect 21633 12612 21699 12613
rect 21582 12548 21588 12612
rect 21652 12610 21699 12612
rect 21652 12608 21744 12610
rect 21694 12552 21744 12608
rect 21652 12550 21744 12552
rect 21652 12548 21699 12550
rect 21633 12547 21699 12548
rect 7110 12544 7426 12545
rect 7110 12480 7116 12544
rect 7180 12480 7196 12544
rect 7260 12480 7276 12544
rect 7340 12480 7356 12544
rect 7420 12480 7426 12544
rect 7110 12479 7426 12480
rect 13826 12544 14142 12545
rect 13826 12480 13832 12544
rect 13896 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14142 12544
rect 13826 12479 14142 12480
rect 20542 12544 20858 12545
rect 20542 12480 20548 12544
rect 20612 12480 20628 12544
rect 20692 12480 20708 12544
rect 20772 12480 20788 12544
rect 20852 12480 20858 12544
rect 20542 12479 20858 12480
rect 27258 12544 27574 12545
rect 27258 12480 27264 12544
rect 27328 12480 27344 12544
rect 27408 12480 27424 12544
rect 27488 12480 27504 12544
rect 27568 12480 27574 12544
rect 27258 12479 27574 12480
rect 7465 12338 7531 12341
rect 10041 12338 10107 12341
rect 7465 12336 10107 12338
rect 7465 12280 7470 12336
rect 7526 12280 10046 12336
rect 10102 12280 10107 12336
rect 7465 12278 10107 12280
rect 7465 12275 7531 12278
rect 10041 12275 10107 12278
rect 15929 12338 15995 12341
rect 16389 12338 16455 12341
rect 25497 12338 25563 12341
rect 15929 12336 25563 12338
rect 15929 12280 15934 12336
rect 15990 12280 16394 12336
rect 16450 12280 25502 12336
rect 25558 12280 25563 12336
rect 15929 12278 25563 12280
rect 15929 12275 15995 12278
rect 16389 12275 16455 12278
rect 25497 12275 25563 12278
rect 26141 12340 26207 12341
rect 26141 12336 26188 12340
rect 26252 12338 26258 12340
rect 26141 12280 26146 12336
rect 26141 12276 26188 12280
rect 26252 12278 26298 12338
rect 26252 12276 26258 12278
rect 26141 12275 26207 12276
rect 3752 12000 4068 12001
rect 3752 11936 3758 12000
rect 3822 11936 3838 12000
rect 3902 11936 3918 12000
rect 3982 11936 3998 12000
rect 4062 11936 4068 12000
rect 3752 11935 4068 11936
rect 10468 12000 10784 12001
rect 10468 11936 10474 12000
rect 10538 11936 10554 12000
rect 10618 11936 10634 12000
rect 10698 11936 10714 12000
rect 10778 11936 10784 12000
rect 10468 11935 10784 11936
rect 17184 12000 17500 12001
rect 17184 11936 17190 12000
rect 17254 11936 17270 12000
rect 17334 11936 17350 12000
rect 17414 11936 17430 12000
rect 17494 11936 17500 12000
rect 17184 11935 17500 11936
rect 23900 12000 24216 12001
rect 23900 11936 23906 12000
rect 23970 11936 23986 12000
rect 24050 11936 24066 12000
rect 24130 11936 24146 12000
rect 24210 11936 24216 12000
rect 23900 11935 24216 11936
rect 14089 11794 14155 11797
rect 18781 11794 18847 11797
rect 14089 11792 18847 11794
rect 14089 11736 14094 11792
rect 14150 11736 18786 11792
rect 18842 11736 18847 11792
rect 14089 11734 18847 11736
rect 14089 11731 14155 11734
rect 18781 11731 18847 11734
rect 7741 11658 7807 11661
rect 14917 11658 14983 11661
rect 7741 11656 14983 11658
rect 7741 11600 7746 11656
rect 7802 11600 14922 11656
rect 14978 11600 14983 11656
rect 7741 11598 14983 11600
rect 7741 11595 7807 11598
rect 14917 11595 14983 11598
rect 19333 11658 19399 11661
rect 19885 11658 19951 11661
rect 19333 11656 19951 11658
rect 19333 11600 19338 11656
rect 19394 11600 19890 11656
rect 19946 11600 19951 11656
rect 19333 11598 19951 11600
rect 19333 11595 19399 11598
rect 19885 11595 19951 11598
rect 7110 11456 7426 11457
rect 7110 11392 7116 11456
rect 7180 11392 7196 11456
rect 7260 11392 7276 11456
rect 7340 11392 7356 11456
rect 7420 11392 7426 11456
rect 7110 11391 7426 11392
rect 13826 11456 14142 11457
rect 13826 11392 13832 11456
rect 13896 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14142 11456
rect 13826 11391 14142 11392
rect 20542 11456 20858 11457
rect 20542 11392 20548 11456
rect 20612 11392 20628 11456
rect 20692 11392 20708 11456
rect 20772 11392 20788 11456
rect 20852 11392 20858 11456
rect 20542 11391 20858 11392
rect 27258 11456 27574 11457
rect 27258 11392 27264 11456
rect 27328 11392 27344 11456
rect 27408 11392 27424 11456
rect 27488 11392 27504 11456
rect 27568 11392 27574 11456
rect 27258 11391 27574 11392
rect 9581 11386 9647 11389
rect 12433 11386 12499 11389
rect 9581 11384 12499 11386
rect 9581 11328 9586 11384
rect 9642 11328 12438 11384
rect 12494 11328 12499 11384
rect 9581 11326 12499 11328
rect 9581 11323 9647 11326
rect 12433 11323 12499 11326
rect 7833 11250 7899 11253
rect 16246 11250 16252 11252
rect 7833 11248 16252 11250
rect 7833 11192 7838 11248
rect 7894 11192 16252 11248
rect 7833 11190 16252 11192
rect 7833 11187 7899 11190
rect 16246 11188 16252 11190
rect 16316 11250 16322 11252
rect 16573 11250 16639 11253
rect 16316 11248 16639 11250
rect 16316 11192 16578 11248
rect 16634 11192 16639 11248
rect 16316 11190 16639 11192
rect 16316 11188 16322 11190
rect 16573 11187 16639 11190
rect 14641 11114 14707 11117
rect 14774 11114 14780 11116
rect 14641 11112 14780 11114
rect 14641 11056 14646 11112
rect 14702 11056 14780 11112
rect 14641 11054 14780 11056
rect 14641 11051 14707 11054
rect 14774 11052 14780 11054
rect 14844 11052 14850 11116
rect 15101 11114 15167 11117
rect 18873 11114 18939 11117
rect 19241 11114 19307 11117
rect 15101 11112 19307 11114
rect 15101 11056 15106 11112
rect 15162 11056 18878 11112
rect 18934 11056 19246 11112
rect 19302 11056 19307 11112
rect 15101 11054 19307 11056
rect 15101 11051 15167 11054
rect 18873 11051 18939 11054
rect 19241 11051 19307 11054
rect 3752 10912 4068 10913
rect 3752 10848 3758 10912
rect 3822 10848 3838 10912
rect 3902 10848 3918 10912
rect 3982 10848 3998 10912
rect 4062 10848 4068 10912
rect 3752 10847 4068 10848
rect 10468 10912 10784 10913
rect 10468 10848 10474 10912
rect 10538 10848 10554 10912
rect 10618 10848 10634 10912
rect 10698 10848 10714 10912
rect 10778 10848 10784 10912
rect 10468 10847 10784 10848
rect 17184 10912 17500 10913
rect 17184 10848 17190 10912
rect 17254 10848 17270 10912
rect 17334 10848 17350 10912
rect 17414 10848 17430 10912
rect 17494 10848 17500 10912
rect 17184 10847 17500 10848
rect 23900 10912 24216 10913
rect 23900 10848 23906 10912
rect 23970 10848 23986 10912
rect 24050 10848 24066 10912
rect 24130 10848 24146 10912
rect 24210 10848 24216 10912
rect 23900 10847 24216 10848
rect 7110 10368 7426 10369
rect 7110 10304 7116 10368
rect 7180 10304 7196 10368
rect 7260 10304 7276 10368
rect 7340 10304 7356 10368
rect 7420 10304 7426 10368
rect 7110 10303 7426 10304
rect 13826 10368 14142 10369
rect 13826 10304 13832 10368
rect 13896 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14142 10368
rect 13826 10303 14142 10304
rect 20542 10368 20858 10369
rect 20542 10304 20548 10368
rect 20612 10304 20628 10368
rect 20692 10304 20708 10368
rect 20772 10304 20788 10368
rect 20852 10304 20858 10368
rect 20542 10303 20858 10304
rect 27258 10368 27574 10369
rect 27258 10304 27264 10368
rect 27328 10304 27344 10368
rect 27408 10304 27424 10368
rect 27488 10304 27504 10368
rect 27568 10304 27574 10368
rect 27258 10303 27574 10304
rect 22001 10162 22067 10165
rect 23381 10162 23447 10165
rect 22001 10160 23447 10162
rect 22001 10104 22006 10160
rect 22062 10104 23386 10160
rect 23442 10104 23447 10160
rect 22001 10102 23447 10104
rect 22001 10099 22067 10102
rect 23381 10099 23447 10102
rect 24393 10026 24459 10029
rect 26417 10026 26483 10029
rect 24393 10024 26483 10026
rect 24393 9968 24398 10024
rect 24454 9968 26422 10024
rect 26478 9968 26483 10024
rect 24393 9966 26483 9968
rect 24393 9963 24459 9966
rect 26417 9963 26483 9966
rect 3752 9824 4068 9825
rect 3752 9760 3758 9824
rect 3822 9760 3838 9824
rect 3902 9760 3918 9824
rect 3982 9760 3998 9824
rect 4062 9760 4068 9824
rect 3752 9759 4068 9760
rect 10468 9824 10784 9825
rect 10468 9760 10474 9824
rect 10538 9760 10554 9824
rect 10618 9760 10634 9824
rect 10698 9760 10714 9824
rect 10778 9760 10784 9824
rect 10468 9759 10784 9760
rect 17184 9824 17500 9825
rect 17184 9760 17190 9824
rect 17254 9760 17270 9824
rect 17334 9760 17350 9824
rect 17414 9760 17430 9824
rect 17494 9760 17500 9824
rect 17184 9759 17500 9760
rect 23900 9824 24216 9825
rect 23900 9760 23906 9824
rect 23970 9760 23986 9824
rect 24050 9760 24066 9824
rect 24130 9760 24146 9824
rect 24210 9760 24216 9824
rect 23900 9759 24216 9760
rect 11462 9556 11468 9620
rect 11532 9618 11538 9620
rect 12433 9618 12499 9621
rect 14457 9618 14523 9621
rect 21582 9618 21588 9620
rect 11532 9616 21588 9618
rect 11532 9560 12438 9616
rect 12494 9560 14462 9616
rect 14518 9560 21588 9616
rect 11532 9558 21588 9560
rect 11532 9556 11538 9558
rect 12433 9555 12499 9558
rect 14457 9555 14523 9558
rect 21582 9556 21588 9558
rect 21652 9556 21658 9620
rect 15745 9482 15811 9485
rect 26182 9482 26188 9484
rect 15745 9480 26188 9482
rect 15745 9424 15750 9480
rect 15806 9424 26188 9480
rect 15745 9422 26188 9424
rect 15745 9419 15811 9422
rect 26182 9420 26188 9422
rect 26252 9420 26258 9484
rect 12433 9346 12499 9349
rect 13353 9346 13419 9349
rect 12433 9344 13419 9346
rect 12433 9288 12438 9344
rect 12494 9288 13358 9344
rect 13414 9288 13419 9344
rect 12433 9286 13419 9288
rect 12433 9283 12499 9286
rect 13353 9283 13419 9286
rect 7110 9280 7426 9281
rect 7110 9216 7116 9280
rect 7180 9216 7196 9280
rect 7260 9216 7276 9280
rect 7340 9216 7356 9280
rect 7420 9216 7426 9280
rect 7110 9215 7426 9216
rect 13826 9280 14142 9281
rect 13826 9216 13832 9280
rect 13896 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14142 9280
rect 13826 9215 14142 9216
rect 20542 9280 20858 9281
rect 20542 9216 20548 9280
rect 20612 9216 20628 9280
rect 20692 9216 20708 9280
rect 20772 9216 20788 9280
rect 20852 9216 20858 9280
rect 20542 9215 20858 9216
rect 27258 9280 27574 9281
rect 27258 9216 27264 9280
rect 27328 9216 27344 9280
rect 27408 9216 27424 9280
rect 27488 9216 27504 9280
rect 27568 9216 27574 9280
rect 27258 9215 27574 9216
rect 5165 9074 5231 9077
rect 10174 9074 10180 9076
rect 5165 9072 10180 9074
rect 5165 9016 5170 9072
rect 5226 9016 10180 9072
rect 5165 9014 10180 9016
rect 5165 9011 5231 9014
rect 10174 9012 10180 9014
rect 10244 9074 10250 9076
rect 16573 9074 16639 9077
rect 17125 9074 17191 9077
rect 10244 9072 17191 9074
rect 10244 9016 16578 9072
rect 16634 9016 17130 9072
rect 17186 9016 17191 9072
rect 10244 9014 17191 9016
rect 10244 9012 10250 9014
rect 16573 9011 16639 9014
rect 17125 9011 17191 9014
rect 3752 8736 4068 8737
rect 3752 8672 3758 8736
rect 3822 8672 3838 8736
rect 3902 8672 3918 8736
rect 3982 8672 3998 8736
rect 4062 8672 4068 8736
rect 3752 8671 4068 8672
rect 10468 8736 10784 8737
rect 10468 8672 10474 8736
rect 10538 8672 10554 8736
rect 10618 8672 10634 8736
rect 10698 8672 10714 8736
rect 10778 8672 10784 8736
rect 10468 8671 10784 8672
rect 17184 8736 17500 8737
rect 17184 8672 17190 8736
rect 17254 8672 17270 8736
rect 17334 8672 17350 8736
rect 17414 8672 17430 8736
rect 17494 8672 17500 8736
rect 17184 8671 17500 8672
rect 23900 8736 24216 8737
rect 23900 8672 23906 8736
rect 23970 8672 23986 8736
rect 24050 8672 24066 8736
rect 24130 8672 24146 8736
rect 24210 8672 24216 8736
rect 23900 8671 24216 8672
rect 12065 8530 12131 8533
rect 17585 8530 17651 8533
rect 12065 8528 17651 8530
rect 12065 8472 12070 8528
rect 12126 8472 17590 8528
rect 17646 8472 17651 8528
rect 12065 8470 17651 8472
rect 12065 8467 12131 8470
rect 17585 8467 17651 8470
rect 3509 8394 3575 8397
rect 17769 8394 17835 8397
rect 3509 8392 17835 8394
rect 3509 8336 3514 8392
rect 3570 8336 17774 8392
rect 17830 8336 17835 8392
rect 3509 8334 17835 8336
rect 3509 8331 3575 8334
rect 17769 8331 17835 8334
rect 7110 8192 7426 8193
rect 7110 8128 7116 8192
rect 7180 8128 7196 8192
rect 7260 8128 7276 8192
rect 7340 8128 7356 8192
rect 7420 8128 7426 8192
rect 7110 8127 7426 8128
rect 13826 8192 14142 8193
rect 13826 8128 13832 8192
rect 13896 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14142 8192
rect 13826 8127 14142 8128
rect 20542 8192 20858 8193
rect 20542 8128 20548 8192
rect 20612 8128 20628 8192
rect 20692 8128 20708 8192
rect 20772 8128 20788 8192
rect 20852 8128 20858 8192
rect 20542 8127 20858 8128
rect 27258 8192 27574 8193
rect 27258 8128 27264 8192
rect 27328 8128 27344 8192
rect 27408 8128 27424 8192
rect 27488 8128 27504 8192
rect 27568 8128 27574 8192
rect 27258 8127 27574 8128
rect 9857 7850 9923 7853
rect 13813 7850 13879 7853
rect 9857 7848 13879 7850
rect 9857 7792 9862 7848
rect 9918 7792 13818 7848
rect 13874 7792 13879 7848
rect 9857 7790 13879 7792
rect 9857 7787 9923 7790
rect 13813 7787 13879 7790
rect 3752 7648 4068 7649
rect 3752 7584 3758 7648
rect 3822 7584 3838 7648
rect 3902 7584 3918 7648
rect 3982 7584 3998 7648
rect 4062 7584 4068 7648
rect 3752 7583 4068 7584
rect 10468 7648 10784 7649
rect 10468 7584 10474 7648
rect 10538 7584 10554 7648
rect 10618 7584 10634 7648
rect 10698 7584 10714 7648
rect 10778 7584 10784 7648
rect 10468 7583 10784 7584
rect 17184 7648 17500 7649
rect 17184 7584 17190 7648
rect 17254 7584 17270 7648
rect 17334 7584 17350 7648
rect 17414 7584 17430 7648
rect 17494 7584 17500 7648
rect 17184 7583 17500 7584
rect 23900 7648 24216 7649
rect 23900 7584 23906 7648
rect 23970 7584 23986 7648
rect 24050 7584 24066 7648
rect 24130 7584 24146 7648
rect 24210 7584 24216 7648
rect 23900 7583 24216 7584
rect 21582 7380 21588 7444
rect 21652 7442 21658 7444
rect 21725 7442 21791 7445
rect 21652 7440 21791 7442
rect 21652 7384 21730 7440
rect 21786 7384 21791 7440
rect 21652 7382 21791 7384
rect 21652 7380 21658 7382
rect 21725 7379 21791 7382
rect 7110 7104 7426 7105
rect 7110 7040 7116 7104
rect 7180 7040 7196 7104
rect 7260 7040 7276 7104
rect 7340 7040 7356 7104
rect 7420 7040 7426 7104
rect 7110 7039 7426 7040
rect 13826 7104 14142 7105
rect 13826 7040 13832 7104
rect 13896 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14142 7104
rect 13826 7039 14142 7040
rect 20542 7104 20858 7105
rect 20542 7040 20548 7104
rect 20612 7040 20628 7104
rect 20692 7040 20708 7104
rect 20772 7040 20788 7104
rect 20852 7040 20858 7104
rect 20542 7039 20858 7040
rect 27258 7104 27574 7105
rect 27258 7040 27264 7104
rect 27328 7040 27344 7104
rect 27408 7040 27424 7104
rect 27488 7040 27504 7104
rect 27568 7040 27574 7104
rect 27258 7039 27574 7040
rect 9213 6898 9279 6901
rect 9397 6898 9463 6901
rect 12801 6898 12867 6901
rect 14457 6900 14523 6901
rect 9213 6896 12867 6898
rect 9213 6840 9218 6896
rect 9274 6840 9402 6896
rect 9458 6840 12806 6896
rect 12862 6840 12867 6896
rect 9213 6838 12867 6840
rect 9213 6835 9279 6838
rect 9397 6835 9463 6838
rect 12801 6835 12867 6838
rect 14406 6836 14412 6900
rect 14476 6898 14523 6900
rect 14476 6896 14568 6898
rect 14518 6840 14568 6896
rect 14476 6838 14568 6840
rect 14476 6836 14523 6838
rect 14457 6835 14523 6836
rect 3752 6560 4068 6561
rect 3752 6496 3758 6560
rect 3822 6496 3838 6560
rect 3902 6496 3918 6560
rect 3982 6496 3998 6560
rect 4062 6496 4068 6560
rect 3752 6495 4068 6496
rect 10468 6560 10784 6561
rect 10468 6496 10474 6560
rect 10538 6496 10554 6560
rect 10618 6496 10634 6560
rect 10698 6496 10714 6560
rect 10778 6496 10784 6560
rect 10468 6495 10784 6496
rect 17184 6560 17500 6561
rect 17184 6496 17190 6560
rect 17254 6496 17270 6560
rect 17334 6496 17350 6560
rect 17414 6496 17430 6560
rect 17494 6496 17500 6560
rect 17184 6495 17500 6496
rect 23900 6560 24216 6561
rect 23900 6496 23906 6560
rect 23970 6496 23986 6560
rect 24050 6496 24066 6560
rect 24130 6496 24146 6560
rect 24210 6496 24216 6560
rect 23900 6495 24216 6496
rect 10593 6354 10659 6357
rect 11881 6354 11947 6357
rect 10593 6352 11947 6354
rect 10593 6296 10598 6352
rect 10654 6296 11886 6352
rect 11942 6296 11947 6352
rect 10593 6294 11947 6296
rect 10593 6291 10659 6294
rect 11881 6291 11947 6294
rect 6361 6218 6427 6221
rect 11462 6218 11468 6220
rect 6361 6216 11468 6218
rect 6361 6160 6366 6216
rect 6422 6160 11468 6216
rect 6361 6158 11468 6160
rect 6361 6155 6427 6158
rect 11462 6156 11468 6158
rect 11532 6156 11538 6220
rect 7110 6016 7426 6017
rect 7110 5952 7116 6016
rect 7180 5952 7196 6016
rect 7260 5952 7276 6016
rect 7340 5952 7356 6016
rect 7420 5952 7426 6016
rect 7110 5951 7426 5952
rect 13826 6016 14142 6017
rect 13826 5952 13832 6016
rect 13896 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14142 6016
rect 13826 5951 14142 5952
rect 20542 6016 20858 6017
rect 20542 5952 20548 6016
rect 20612 5952 20628 6016
rect 20692 5952 20708 6016
rect 20772 5952 20788 6016
rect 20852 5952 20858 6016
rect 20542 5951 20858 5952
rect 27258 6016 27574 6017
rect 27258 5952 27264 6016
rect 27328 5952 27344 6016
rect 27408 5952 27424 6016
rect 27488 5952 27504 6016
rect 27568 5952 27574 6016
rect 27258 5951 27574 5952
rect 10777 5674 10843 5677
rect 16941 5674 17007 5677
rect 17309 5674 17375 5677
rect 10777 5672 17375 5674
rect 10777 5616 10782 5672
rect 10838 5616 16946 5672
rect 17002 5616 17314 5672
rect 17370 5616 17375 5672
rect 10777 5614 17375 5616
rect 10777 5611 10843 5614
rect 16941 5611 17007 5614
rect 17309 5611 17375 5614
rect 3752 5472 4068 5473
rect 3752 5408 3758 5472
rect 3822 5408 3838 5472
rect 3902 5408 3918 5472
rect 3982 5408 3998 5472
rect 4062 5408 4068 5472
rect 3752 5407 4068 5408
rect 10468 5472 10784 5473
rect 10468 5408 10474 5472
rect 10538 5408 10554 5472
rect 10618 5408 10634 5472
rect 10698 5408 10714 5472
rect 10778 5408 10784 5472
rect 10468 5407 10784 5408
rect 17184 5472 17500 5473
rect 17184 5408 17190 5472
rect 17254 5408 17270 5472
rect 17334 5408 17350 5472
rect 17414 5408 17430 5472
rect 17494 5408 17500 5472
rect 17184 5407 17500 5408
rect 23900 5472 24216 5473
rect 23900 5408 23906 5472
rect 23970 5408 23986 5472
rect 24050 5408 24066 5472
rect 24130 5408 24146 5472
rect 24210 5408 24216 5472
rect 23900 5407 24216 5408
rect 11421 5268 11487 5269
rect 11421 5266 11468 5268
rect 11376 5264 11468 5266
rect 11376 5208 11426 5264
rect 11376 5206 11468 5208
rect 11421 5204 11468 5206
rect 11532 5204 11538 5268
rect 11421 5203 11487 5204
rect 7110 4928 7426 4929
rect 7110 4864 7116 4928
rect 7180 4864 7196 4928
rect 7260 4864 7276 4928
rect 7340 4864 7356 4928
rect 7420 4864 7426 4928
rect 7110 4863 7426 4864
rect 13826 4928 14142 4929
rect 13826 4864 13832 4928
rect 13896 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14142 4928
rect 13826 4863 14142 4864
rect 20542 4928 20858 4929
rect 20542 4864 20548 4928
rect 20612 4864 20628 4928
rect 20692 4864 20708 4928
rect 20772 4864 20788 4928
rect 20852 4864 20858 4928
rect 20542 4863 20858 4864
rect 27258 4928 27574 4929
rect 27258 4864 27264 4928
rect 27328 4864 27344 4928
rect 27408 4864 27424 4928
rect 27488 4864 27504 4928
rect 27568 4864 27574 4928
rect 27258 4863 27574 4864
rect 8845 4722 8911 4725
rect 9305 4722 9371 4725
rect 8845 4720 9371 4722
rect 8845 4664 8850 4720
rect 8906 4664 9310 4720
rect 9366 4664 9371 4720
rect 8845 4662 9371 4664
rect 8845 4659 8911 4662
rect 9305 4659 9371 4662
rect 3752 4384 4068 4385
rect 3752 4320 3758 4384
rect 3822 4320 3838 4384
rect 3902 4320 3918 4384
rect 3982 4320 3998 4384
rect 4062 4320 4068 4384
rect 3752 4319 4068 4320
rect 10468 4384 10784 4385
rect 10468 4320 10474 4384
rect 10538 4320 10554 4384
rect 10618 4320 10634 4384
rect 10698 4320 10714 4384
rect 10778 4320 10784 4384
rect 10468 4319 10784 4320
rect 17184 4384 17500 4385
rect 17184 4320 17190 4384
rect 17254 4320 17270 4384
rect 17334 4320 17350 4384
rect 17414 4320 17430 4384
rect 17494 4320 17500 4384
rect 17184 4319 17500 4320
rect 23900 4384 24216 4385
rect 23900 4320 23906 4384
rect 23970 4320 23986 4384
rect 24050 4320 24066 4384
rect 24130 4320 24146 4384
rect 24210 4320 24216 4384
rect 23900 4319 24216 4320
rect 7110 3840 7426 3841
rect 7110 3776 7116 3840
rect 7180 3776 7196 3840
rect 7260 3776 7276 3840
rect 7340 3776 7356 3840
rect 7420 3776 7426 3840
rect 7110 3775 7426 3776
rect 13826 3840 14142 3841
rect 13826 3776 13832 3840
rect 13896 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14142 3840
rect 13826 3775 14142 3776
rect 20542 3840 20858 3841
rect 20542 3776 20548 3840
rect 20612 3776 20628 3840
rect 20692 3776 20708 3840
rect 20772 3776 20788 3840
rect 20852 3776 20858 3840
rect 20542 3775 20858 3776
rect 27258 3840 27574 3841
rect 27258 3776 27264 3840
rect 27328 3776 27344 3840
rect 27408 3776 27424 3840
rect 27488 3776 27504 3840
rect 27568 3776 27574 3840
rect 27258 3775 27574 3776
rect 3752 3296 4068 3297
rect 3752 3232 3758 3296
rect 3822 3232 3838 3296
rect 3902 3232 3918 3296
rect 3982 3232 3998 3296
rect 4062 3232 4068 3296
rect 3752 3231 4068 3232
rect 10468 3296 10784 3297
rect 10468 3232 10474 3296
rect 10538 3232 10554 3296
rect 10618 3232 10634 3296
rect 10698 3232 10714 3296
rect 10778 3232 10784 3296
rect 10468 3231 10784 3232
rect 17184 3296 17500 3297
rect 17184 3232 17190 3296
rect 17254 3232 17270 3296
rect 17334 3232 17350 3296
rect 17414 3232 17430 3296
rect 17494 3232 17500 3296
rect 17184 3231 17500 3232
rect 23900 3296 24216 3297
rect 23900 3232 23906 3296
rect 23970 3232 23986 3296
rect 24050 3232 24066 3296
rect 24130 3232 24146 3296
rect 24210 3232 24216 3296
rect 23900 3231 24216 3232
rect 7110 2752 7426 2753
rect 7110 2688 7116 2752
rect 7180 2688 7196 2752
rect 7260 2688 7276 2752
rect 7340 2688 7356 2752
rect 7420 2688 7426 2752
rect 7110 2687 7426 2688
rect 13826 2752 14142 2753
rect 13826 2688 13832 2752
rect 13896 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14142 2752
rect 13826 2687 14142 2688
rect 20542 2752 20858 2753
rect 20542 2688 20548 2752
rect 20612 2688 20628 2752
rect 20692 2688 20708 2752
rect 20772 2688 20788 2752
rect 20852 2688 20858 2752
rect 20542 2687 20858 2688
rect 27258 2752 27574 2753
rect 27258 2688 27264 2752
rect 27328 2688 27344 2752
rect 27408 2688 27424 2752
rect 27488 2688 27504 2752
rect 27568 2688 27574 2752
rect 27258 2687 27574 2688
rect 14641 2682 14707 2685
rect 14774 2682 14780 2684
rect 14641 2680 14780 2682
rect 14641 2624 14646 2680
rect 14702 2624 14780 2680
rect 14641 2622 14780 2624
rect 14641 2619 14707 2622
rect 14774 2620 14780 2622
rect 14844 2620 14850 2684
rect 6453 2546 6519 2549
rect 19374 2546 19380 2548
rect 6453 2544 19380 2546
rect 6453 2488 6458 2544
rect 6514 2488 19380 2544
rect 6453 2486 19380 2488
rect 6453 2483 6519 2486
rect 19374 2484 19380 2486
rect 19444 2484 19450 2548
rect 8937 2410 9003 2413
rect 20294 2410 20300 2412
rect 8937 2408 20300 2410
rect 8937 2352 8942 2408
rect 8998 2352 20300 2408
rect 8937 2350 20300 2352
rect 8937 2347 9003 2350
rect 20294 2348 20300 2350
rect 20364 2348 20370 2412
rect 3752 2208 4068 2209
rect 3752 2144 3758 2208
rect 3822 2144 3838 2208
rect 3902 2144 3918 2208
rect 3982 2144 3998 2208
rect 4062 2144 4068 2208
rect 3752 2143 4068 2144
rect 10468 2208 10784 2209
rect 10468 2144 10474 2208
rect 10538 2144 10554 2208
rect 10618 2144 10634 2208
rect 10698 2144 10714 2208
rect 10778 2144 10784 2208
rect 10468 2143 10784 2144
rect 17184 2208 17500 2209
rect 17184 2144 17190 2208
rect 17254 2144 17270 2208
rect 17334 2144 17350 2208
rect 17414 2144 17430 2208
rect 17494 2144 17500 2208
rect 17184 2143 17500 2144
rect 23900 2208 24216 2209
rect 23900 2144 23906 2208
rect 23970 2144 23986 2208
rect 24050 2144 24066 2208
rect 24130 2144 24146 2208
rect 24210 2144 24216 2208
rect 23900 2143 24216 2144
rect 5993 2002 6059 2005
rect 18413 2002 18479 2005
rect 20253 2004 20319 2005
rect 20253 2002 20300 2004
rect 5993 2000 18479 2002
rect 5993 1944 5998 2000
rect 6054 1944 18418 2000
rect 18474 1944 18479 2000
rect 5993 1942 18479 1944
rect 20208 2000 20300 2002
rect 20208 1944 20258 2000
rect 20208 1942 20300 1944
rect 5993 1939 6059 1942
rect 18413 1939 18479 1942
rect 20253 1940 20300 1942
rect 20364 1940 20370 2004
rect 20253 1939 20319 1940
rect 841 1866 907 1869
rect 15285 1866 15351 1869
rect 841 1864 15351 1866
rect 841 1808 846 1864
rect 902 1808 15290 1864
rect 15346 1808 15351 1864
rect 841 1806 15351 1808
rect 841 1803 907 1806
rect 15285 1803 15351 1806
rect 7110 1664 7426 1665
rect 7110 1600 7116 1664
rect 7180 1600 7196 1664
rect 7260 1600 7276 1664
rect 7340 1600 7356 1664
rect 7420 1600 7426 1664
rect 7110 1599 7426 1600
rect 13826 1664 14142 1665
rect 13826 1600 13832 1664
rect 13896 1600 13912 1664
rect 13976 1600 13992 1664
rect 14056 1600 14072 1664
rect 14136 1600 14142 1664
rect 13826 1599 14142 1600
rect 20542 1664 20858 1665
rect 20542 1600 20548 1664
rect 20612 1600 20628 1664
rect 20692 1600 20708 1664
rect 20772 1600 20788 1664
rect 20852 1600 20858 1664
rect 20542 1599 20858 1600
rect 27258 1664 27574 1665
rect 27258 1600 27264 1664
rect 27328 1600 27344 1664
rect 27408 1600 27424 1664
rect 27488 1600 27504 1664
rect 27568 1600 27574 1664
rect 27258 1599 27574 1600
rect 16530 1534 19626 1594
rect 7465 1458 7531 1461
rect 7925 1458 7991 1461
rect 16530 1458 16590 1534
rect 7465 1456 16590 1458
rect 7465 1400 7470 1456
rect 7526 1400 7930 1456
rect 7986 1400 16590 1456
rect 7465 1398 16590 1400
rect 18965 1458 19031 1461
rect 19374 1458 19380 1460
rect 18965 1456 19380 1458
rect 18965 1400 18970 1456
rect 19026 1400 19380 1456
rect 18965 1398 19380 1400
rect 7465 1395 7531 1398
rect 7925 1395 7991 1398
rect 18965 1395 19031 1398
rect 19374 1396 19380 1398
rect 19444 1396 19450 1460
rect 19566 1458 19626 1534
rect 22001 1458 22067 1461
rect 19566 1456 22067 1458
rect 19566 1400 22006 1456
rect 22062 1400 22067 1456
rect 19566 1398 22067 1400
rect 22001 1395 22067 1398
rect 3752 1120 4068 1121
rect 3752 1056 3758 1120
rect 3822 1056 3838 1120
rect 3902 1056 3918 1120
rect 3982 1056 3998 1120
rect 4062 1056 4068 1120
rect 3752 1055 4068 1056
rect 10468 1120 10784 1121
rect 10468 1056 10474 1120
rect 10538 1056 10554 1120
rect 10618 1056 10634 1120
rect 10698 1056 10714 1120
rect 10778 1056 10784 1120
rect 10468 1055 10784 1056
rect 17184 1120 17500 1121
rect 17184 1056 17190 1120
rect 17254 1056 17270 1120
rect 17334 1056 17350 1120
rect 17414 1056 17430 1120
rect 17494 1056 17500 1120
rect 17184 1055 17500 1056
rect 23900 1120 24216 1121
rect 23900 1056 23906 1120
rect 23970 1056 23986 1120
rect 24050 1056 24066 1120
rect 24130 1056 24146 1120
rect 24210 1056 24216 1120
rect 23900 1055 24216 1056
rect 16113 914 16179 917
rect 16246 914 16252 916
rect 16113 912 16252 914
rect 16113 856 16118 912
rect 16174 856 16252 912
rect 16113 854 16252 856
rect 16113 851 16179 854
rect 16246 852 16252 854
rect 16316 852 16322 916
rect 7110 576 7426 577
rect 7110 512 7116 576
rect 7180 512 7196 576
rect 7260 512 7276 576
rect 7340 512 7356 576
rect 7420 512 7426 576
rect 7110 511 7426 512
rect 13826 576 14142 577
rect 13826 512 13832 576
rect 13896 512 13912 576
rect 13976 512 13992 576
rect 14056 512 14072 576
rect 14136 512 14142 576
rect 13826 511 14142 512
rect 20542 576 20858 577
rect 20542 512 20548 576
rect 20612 512 20628 576
rect 20692 512 20708 576
rect 20772 512 20788 576
rect 20852 512 20858 576
rect 20542 511 20858 512
rect 27258 576 27574 577
rect 27258 512 27264 576
rect 27328 512 27344 576
rect 27408 512 27424 576
rect 27488 512 27504 576
rect 27568 512 27574 576
rect 27258 511 27574 512
<< via3 >>
rect 3758 17436 3822 17440
rect 3758 17380 3762 17436
rect 3762 17380 3818 17436
rect 3818 17380 3822 17436
rect 3758 17376 3822 17380
rect 3838 17436 3902 17440
rect 3838 17380 3842 17436
rect 3842 17380 3898 17436
rect 3898 17380 3902 17436
rect 3838 17376 3902 17380
rect 3918 17436 3982 17440
rect 3918 17380 3922 17436
rect 3922 17380 3978 17436
rect 3978 17380 3982 17436
rect 3918 17376 3982 17380
rect 3998 17436 4062 17440
rect 3998 17380 4002 17436
rect 4002 17380 4058 17436
rect 4058 17380 4062 17436
rect 3998 17376 4062 17380
rect 10474 17436 10538 17440
rect 10474 17380 10478 17436
rect 10478 17380 10534 17436
rect 10534 17380 10538 17436
rect 10474 17376 10538 17380
rect 10554 17436 10618 17440
rect 10554 17380 10558 17436
rect 10558 17380 10614 17436
rect 10614 17380 10618 17436
rect 10554 17376 10618 17380
rect 10634 17436 10698 17440
rect 10634 17380 10638 17436
rect 10638 17380 10694 17436
rect 10694 17380 10698 17436
rect 10634 17376 10698 17380
rect 10714 17436 10778 17440
rect 10714 17380 10718 17436
rect 10718 17380 10774 17436
rect 10774 17380 10778 17436
rect 10714 17376 10778 17380
rect 17190 17436 17254 17440
rect 17190 17380 17194 17436
rect 17194 17380 17250 17436
rect 17250 17380 17254 17436
rect 17190 17376 17254 17380
rect 17270 17436 17334 17440
rect 17270 17380 17274 17436
rect 17274 17380 17330 17436
rect 17330 17380 17334 17436
rect 17270 17376 17334 17380
rect 17350 17436 17414 17440
rect 17350 17380 17354 17436
rect 17354 17380 17410 17436
rect 17410 17380 17414 17436
rect 17350 17376 17414 17380
rect 17430 17436 17494 17440
rect 17430 17380 17434 17436
rect 17434 17380 17490 17436
rect 17490 17380 17494 17436
rect 17430 17376 17494 17380
rect 23906 17436 23970 17440
rect 23906 17380 23910 17436
rect 23910 17380 23966 17436
rect 23966 17380 23970 17436
rect 23906 17376 23970 17380
rect 23986 17436 24050 17440
rect 23986 17380 23990 17436
rect 23990 17380 24046 17436
rect 24046 17380 24050 17436
rect 23986 17376 24050 17380
rect 24066 17436 24130 17440
rect 24066 17380 24070 17436
rect 24070 17380 24126 17436
rect 24126 17380 24130 17436
rect 24066 17376 24130 17380
rect 24146 17436 24210 17440
rect 24146 17380 24150 17436
rect 24150 17380 24206 17436
rect 24206 17380 24210 17436
rect 24146 17376 24210 17380
rect 7116 16892 7180 16896
rect 7116 16836 7120 16892
rect 7120 16836 7176 16892
rect 7176 16836 7180 16892
rect 7116 16832 7180 16836
rect 7196 16892 7260 16896
rect 7196 16836 7200 16892
rect 7200 16836 7256 16892
rect 7256 16836 7260 16892
rect 7196 16832 7260 16836
rect 7276 16892 7340 16896
rect 7276 16836 7280 16892
rect 7280 16836 7336 16892
rect 7336 16836 7340 16892
rect 7276 16832 7340 16836
rect 7356 16892 7420 16896
rect 7356 16836 7360 16892
rect 7360 16836 7416 16892
rect 7416 16836 7420 16892
rect 7356 16832 7420 16836
rect 13832 16892 13896 16896
rect 13832 16836 13836 16892
rect 13836 16836 13892 16892
rect 13892 16836 13896 16892
rect 13832 16832 13896 16836
rect 13912 16892 13976 16896
rect 13912 16836 13916 16892
rect 13916 16836 13972 16892
rect 13972 16836 13976 16892
rect 13912 16832 13976 16836
rect 13992 16892 14056 16896
rect 13992 16836 13996 16892
rect 13996 16836 14052 16892
rect 14052 16836 14056 16892
rect 13992 16832 14056 16836
rect 14072 16892 14136 16896
rect 14072 16836 14076 16892
rect 14076 16836 14132 16892
rect 14132 16836 14136 16892
rect 14072 16832 14136 16836
rect 20548 16892 20612 16896
rect 20548 16836 20552 16892
rect 20552 16836 20608 16892
rect 20608 16836 20612 16892
rect 20548 16832 20612 16836
rect 20628 16892 20692 16896
rect 20628 16836 20632 16892
rect 20632 16836 20688 16892
rect 20688 16836 20692 16892
rect 20628 16832 20692 16836
rect 20708 16892 20772 16896
rect 20708 16836 20712 16892
rect 20712 16836 20768 16892
rect 20768 16836 20772 16892
rect 20708 16832 20772 16836
rect 20788 16892 20852 16896
rect 20788 16836 20792 16892
rect 20792 16836 20848 16892
rect 20848 16836 20852 16892
rect 20788 16832 20852 16836
rect 27264 16892 27328 16896
rect 27264 16836 27268 16892
rect 27268 16836 27324 16892
rect 27324 16836 27328 16892
rect 27264 16832 27328 16836
rect 27344 16892 27408 16896
rect 27344 16836 27348 16892
rect 27348 16836 27404 16892
rect 27404 16836 27408 16892
rect 27344 16832 27408 16836
rect 27424 16892 27488 16896
rect 27424 16836 27428 16892
rect 27428 16836 27484 16892
rect 27484 16836 27488 16892
rect 27424 16832 27488 16836
rect 27504 16892 27568 16896
rect 27504 16836 27508 16892
rect 27508 16836 27564 16892
rect 27564 16836 27568 16892
rect 27504 16832 27568 16836
rect 14412 16628 14476 16692
rect 19380 16688 19444 16692
rect 19380 16632 19394 16688
rect 19394 16632 19444 16688
rect 19380 16628 19444 16632
rect 20300 16628 20364 16692
rect 3758 16348 3822 16352
rect 3758 16292 3762 16348
rect 3762 16292 3818 16348
rect 3818 16292 3822 16348
rect 3758 16288 3822 16292
rect 3838 16348 3902 16352
rect 3838 16292 3842 16348
rect 3842 16292 3898 16348
rect 3898 16292 3902 16348
rect 3838 16288 3902 16292
rect 3918 16348 3982 16352
rect 3918 16292 3922 16348
rect 3922 16292 3978 16348
rect 3978 16292 3982 16348
rect 3918 16288 3982 16292
rect 3998 16348 4062 16352
rect 3998 16292 4002 16348
rect 4002 16292 4058 16348
rect 4058 16292 4062 16348
rect 3998 16288 4062 16292
rect 10474 16348 10538 16352
rect 10474 16292 10478 16348
rect 10478 16292 10534 16348
rect 10534 16292 10538 16348
rect 10474 16288 10538 16292
rect 10554 16348 10618 16352
rect 10554 16292 10558 16348
rect 10558 16292 10614 16348
rect 10614 16292 10618 16348
rect 10554 16288 10618 16292
rect 10634 16348 10698 16352
rect 10634 16292 10638 16348
rect 10638 16292 10694 16348
rect 10694 16292 10698 16348
rect 10634 16288 10698 16292
rect 10714 16348 10778 16352
rect 10714 16292 10718 16348
rect 10718 16292 10774 16348
rect 10774 16292 10778 16348
rect 10714 16288 10778 16292
rect 17190 16348 17254 16352
rect 17190 16292 17194 16348
rect 17194 16292 17250 16348
rect 17250 16292 17254 16348
rect 17190 16288 17254 16292
rect 17270 16348 17334 16352
rect 17270 16292 17274 16348
rect 17274 16292 17330 16348
rect 17330 16292 17334 16348
rect 17270 16288 17334 16292
rect 17350 16348 17414 16352
rect 17350 16292 17354 16348
rect 17354 16292 17410 16348
rect 17410 16292 17414 16348
rect 17350 16288 17414 16292
rect 17430 16348 17494 16352
rect 17430 16292 17434 16348
rect 17434 16292 17490 16348
rect 17490 16292 17494 16348
rect 17430 16288 17494 16292
rect 23906 16348 23970 16352
rect 23906 16292 23910 16348
rect 23910 16292 23966 16348
rect 23966 16292 23970 16348
rect 23906 16288 23970 16292
rect 23986 16348 24050 16352
rect 23986 16292 23990 16348
rect 23990 16292 24046 16348
rect 24046 16292 24050 16348
rect 23986 16288 24050 16292
rect 24066 16348 24130 16352
rect 24066 16292 24070 16348
rect 24070 16292 24126 16348
rect 24126 16292 24130 16348
rect 24066 16288 24130 16292
rect 24146 16348 24210 16352
rect 24146 16292 24150 16348
rect 24150 16292 24206 16348
rect 24206 16292 24210 16348
rect 24146 16288 24210 16292
rect 7116 15804 7180 15808
rect 7116 15748 7120 15804
rect 7120 15748 7176 15804
rect 7176 15748 7180 15804
rect 7116 15744 7180 15748
rect 7196 15804 7260 15808
rect 7196 15748 7200 15804
rect 7200 15748 7256 15804
rect 7256 15748 7260 15804
rect 7196 15744 7260 15748
rect 7276 15804 7340 15808
rect 7276 15748 7280 15804
rect 7280 15748 7336 15804
rect 7336 15748 7340 15804
rect 7276 15744 7340 15748
rect 7356 15804 7420 15808
rect 7356 15748 7360 15804
rect 7360 15748 7416 15804
rect 7416 15748 7420 15804
rect 7356 15744 7420 15748
rect 13832 15804 13896 15808
rect 13832 15748 13836 15804
rect 13836 15748 13892 15804
rect 13892 15748 13896 15804
rect 13832 15744 13896 15748
rect 13912 15804 13976 15808
rect 13912 15748 13916 15804
rect 13916 15748 13972 15804
rect 13972 15748 13976 15804
rect 13912 15744 13976 15748
rect 13992 15804 14056 15808
rect 13992 15748 13996 15804
rect 13996 15748 14052 15804
rect 14052 15748 14056 15804
rect 13992 15744 14056 15748
rect 14072 15804 14136 15808
rect 14072 15748 14076 15804
rect 14076 15748 14132 15804
rect 14132 15748 14136 15804
rect 14072 15744 14136 15748
rect 20548 15804 20612 15808
rect 20548 15748 20552 15804
rect 20552 15748 20608 15804
rect 20608 15748 20612 15804
rect 20548 15744 20612 15748
rect 20628 15804 20692 15808
rect 20628 15748 20632 15804
rect 20632 15748 20688 15804
rect 20688 15748 20692 15804
rect 20628 15744 20692 15748
rect 20708 15804 20772 15808
rect 20708 15748 20712 15804
rect 20712 15748 20768 15804
rect 20768 15748 20772 15804
rect 20708 15744 20772 15748
rect 20788 15804 20852 15808
rect 20788 15748 20792 15804
rect 20792 15748 20848 15804
rect 20848 15748 20852 15804
rect 20788 15744 20852 15748
rect 27264 15804 27328 15808
rect 27264 15748 27268 15804
rect 27268 15748 27324 15804
rect 27324 15748 27328 15804
rect 27264 15744 27328 15748
rect 27344 15804 27408 15808
rect 27344 15748 27348 15804
rect 27348 15748 27404 15804
rect 27404 15748 27408 15804
rect 27344 15744 27408 15748
rect 27424 15804 27488 15808
rect 27424 15748 27428 15804
rect 27428 15748 27484 15804
rect 27484 15748 27488 15804
rect 27424 15744 27488 15748
rect 27504 15804 27568 15808
rect 27504 15748 27508 15804
rect 27508 15748 27564 15804
rect 27564 15748 27568 15804
rect 27504 15744 27568 15748
rect 10180 15268 10244 15332
rect 3758 15260 3822 15264
rect 3758 15204 3762 15260
rect 3762 15204 3818 15260
rect 3818 15204 3822 15260
rect 3758 15200 3822 15204
rect 3838 15260 3902 15264
rect 3838 15204 3842 15260
rect 3842 15204 3898 15260
rect 3898 15204 3902 15260
rect 3838 15200 3902 15204
rect 3918 15260 3982 15264
rect 3918 15204 3922 15260
rect 3922 15204 3978 15260
rect 3978 15204 3982 15260
rect 3918 15200 3982 15204
rect 3998 15260 4062 15264
rect 3998 15204 4002 15260
rect 4002 15204 4058 15260
rect 4058 15204 4062 15260
rect 3998 15200 4062 15204
rect 10474 15260 10538 15264
rect 10474 15204 10478 15260
rect 10478 15204 10534 15260
rect 10534 15204 10538 15260
rect 10474 15200 10538 15204
rect 10554 15260 10618 15264
rect 10554 15204 10558 15260
rect 10558 15204 10614 15260
rect 10614 15204 10618 15260
rect 10554 15200 10618 15204
rect 10634 15260 10698 15264
rect 10634 15204 10638 15260
rect 10638 15204 10694 15260
rect 10694 15204 10698 15260
rect 10634 15200 10698 15204
rect 10714 15260 10778 15264
rect 10714 15204 10718 15260
rect 10718 15204 10774 15260
rect 10774 15204 10778 15260
rect 10714 15200 10778 15204
rect 17190 15260 17254 15264
rect 17190 15204 17194 15260
rect 17194 15204 17250 15260
rect 17250 15204 17254 15260
rect 17190 15200 17254 15204
rect 17270 15260 17334 15264
rect 17270 15204 17274 15260
rect 17274 15204 17330 15260
rect 17330 15204 17334 15260
rect 17270 15200 17334 15204
rect 17350 15260 17414 15264
rect 17350 15204 17354 15260
rect 17354 15204 17410 15260
rect 17410 15204 17414 15260
rect 17350 15200 17414 15204
rect 17430 15260 17494 15264
rect 17430 15204 17434 15260
rect 17434 15204 17490 15260
rect 17490 15204 17494 15260
rect 17430 15200 17494 15204
rect 23906 15260 23970 15264
rect 23906 15204 23910 15260
rect 23910 15204 23966 15260
rect 23966 15204 23970 15260
rect 23906 15200 23970 15204
rect 23986 15260 24050 15264
rect 23986 15204 23990 15260
rect 23990 15204 24046 15260
rect 24046 15204 24050 15260
rect 23986 15200 24050 15204
rect 24066 15260 24130 15264
rect 24066 15204 24070 15260
rect 24070 15204 24126 15260
rect 24126 15204 24130 15260
rect 24066 15200 24130 15204
rect 24146 15260 24210 15264
rect 24146 15204 24150 15260
rect 24150 15204 24206 15260
rect 24206 15204 24210 15260
rect 24146 15200 24210 15204
rect 7116 14716 7180 14720
rect 7116 14660 7120 14716
rect 7120 14660 7176 14716
rect 7176 14660 7180 14716
rect 7116 14656 7180 14660
rect 7196 14716 7260 14720
rect 7196 14660 7200 14716
rect 7200 14660 7256 14716
rect 7256 14660 7260 14716
rect 7196 14656 7260 14660
rect 7276 14716 7340 14720
rect 7276 14660 7280 14716
rect 7280 14660 7336 14716
rect 7336 14660 7340 14716
rect 7276 14656 7340 14660
rect 7356 14716 7420 14720
rect 7356 14660 7360 14716
rect 7360 14660 7416 14716
rect 7416 14660 7420 14716
rect 7356 14656 7420 14660
rect 13832 14716 13896 14720
rect 13832 14660 13836 14716
rect 13836 14660 13892 14716
rect 13892 14660 13896 14716
rect 13832 14656 13896 14660
rect 13912 14716 13976 14720
rect 13912 14660 13916 14716
rect 13916 14660 13972 14716
rect 13972 14660 13976 14716
rect 13912 14656 13976 14660
rect 13992 14716 14056 14720
rect 13992 14660 13996 14716
rect 13996 14660 14052 14716
rect 14052 14660 14056 14716
rect 13992 14656 14056 14660
rect 14072 14716 14136 14720
rect 14072 14660 14076 14716
rect 14076 14660 14132 14716
rect 14132 14660 14136 14716
rect 14072 14656 14136 14660
rect 20548 14716 20612 14720
rect 20548 14660 20552 14716
rect 20552 14660 20608 14716
rect 20608 14660 20612 14716
rect 20548 14656 20612 14660
rect 20628 14716 20692 14720
rect 20628 14660 20632 14716
rect 20632 14660 20688 14716
rect 20688 14660 20692 14716
rect 20628 14656 20692 14660
rect 20708 14716 20772 14720
rect 20708 14660 20712 14716
rect 20712 14660 20768 14716
rect 20768 14660 20772 14716
rect 20708 14656 20772 14660
rect 20788 14716 20852 14720
rect 20788 14660 20792 14716
rect 20792 14660 20848 14716
rect 20848 14660 20852 14716
rect 20788 14656 20852 14660
rect 27264 14716 27328 14720
rect 27264 14660 27268 14716
rect 27268 14660 27324 14716
rect 27324 14660 27328 14716
rect 27264 14656 27328 14660
rect 27344 14716 27408 14720
rect 27344 14660 27348 14716
rect 27348 14660 27404 14716
rect 27404 14660 27408 14716
rect 27344 14656 27408 14660
rect 27424 14716 27488 14720
rect 27424 14660 27428 14716
rect 27428 14660 27484 14716
rect 27484 14660 27488 14716
rect 27424 14656 27488 14660
rect 27504 14716 27568 14720
rect 27504 14660 27508 14716
rect 27508 14660 27564 14716
rect 27564 14660 27568 14716
rect 27504 14656 27568 14660
rect 3758 14172 3822 14176
rect 3758 14116 3762 14172
rect 3762 14116 3818 14172
rect 3818 14116 3822 14172
rect 3758 14112 3822 14116
rect 3838 14172 3902 14176
rect 3838 14116 3842 14172
rect 3842 14116 3898 14172
rect 3898 14116 3902 14172
rect 3838 14112 3902 14116
rect 3918 14172 3982 14176
rect 3918 14116 3922 14172
rect 3922 14116 3978 14172
rect 3978 14116 3982 14172
rect 3918 14112 3982 14116
rect 3998 14172 4062 14176
rect 3998 14116 4002 14172
rect 4002 14116 4058 14172
rect 4058 14116 4062 14172
rect 3998 14112 4062 14116
rect 10474 14172 10538 14176
rect 10474 14116 10478 14172
rect 10478 14116 10534 14172
rect 10534 14116 10538 14172
rect 10474 14112 10538 14116
rect 10554 14172 10618 14176
rect 10554 14116 10558 14172
rect 10558 14116 10614 14172
rect 10614 14116 10618 14172
rect 10554 14112 10618 14116
rect 10634 14172 10698 14176
rect 10634 14116 10638 14172
rect 10638 14116 10694 14172
rect 10694 14116 10698 14172
rect 10634 14112 10698 14116
rect 10714 14172 10778 14176
rect 10714 14116 10718 14172
rect 10718 14116 10774 14172
rect 10774 14116 10778 14172
rect 10714 14112 10778 14116
rect 17190 14172 17254 14176
rect 17190 14116 17194 14172
rect 17194 14116 17250 14172
rect 17250 14116 17254 14172
rect 17190 14112 17254 14116
rect 17270 14172 17334 14176
rect 17270 14116 17274 14172
rect 17274 14116 17330 14172
rect 17330 14116 17334 14172
rect 17270 14112 17334 14116
rect 17350 14172 17414 14176
rect 17350 14116 17354 14172
rect 17354 14116 17410 14172
rect 17410 14116 17414 14172
rect 17350 14112 17414 14116
rect 17430 14172 17494 14176
rect 17430 14116 17434 14172
rect 17434 14116 17490 14172
rect 17490 14116 17494 14172
rect 17430 14112 17494 14116
rect 23906 14172 23970 14176
rect 23906 14116 23910 14172
rect 23910 14116 23966 14172
rect 23966 14116 23970 14172
rect 23906 14112 23970 14116
rect 23986 14172 24050 14176
rect 23986 14116 23990 14172
rect 23990 14116 24046 14172
rect 24046 14116 24050 14172
rect 23986 14112 24050 14116
rect 24066 14172 24130 14176
rect 24066 14116 24070 14172
rect 24070 14116 24126 14172
rect 24126 14116 24130 14172
rect 24066 14112 24130 14116
rect 24146 14172 24210 14176
rect 24146 14116 24150 14172
rect 24150 14116 24206 14172
rect 24206 14116 24210 14172
rect 24146 14112 24210 14116
rect 7116 13628 7180 13632
rect 7116 13572 7120 13628
rect 7120 13572 7176 13628
rect 7176 13572 7180 13628
rect 7116 13568 7180 13572
rect 7196 13628 7260 13632
rect 7196 13572 7200 13628
rect 7200 13572 7256 13628
rect 7256 13572 7260 13628
rect 7196 13568 7260 13572
rect 7276 13628 7340 13632
rect 7276 13572 7280 13628
rect 7280 13572 7336 13628
rect 7336 13572 7340 13628
rect 7276 13568 7340 13572
rect 7356 13628 7420 13632
rect 7356 13572 7360 13628
rect 7360 13572 7416 13628
rect 7416 13572 7420 13628
rect 7356 13568 7420 13572
rect 13832 13628 13896 13632
rect 13832 13572 13836 13628
rect 13836 13572 13892 13628
rect 13892 13572 13896 13628
rect 13832 13568 13896 13572
rect 13912 13628 13976 13632
rect 13912 13572 13916 13628
rect 13916 13572 13972 13628
rect 13972 13572 13976 13628
rect 13912 13568 13976 13572
rect 13992 13628 14056 13632
rect 13992 13572 13996 13628
rect 13996 13572 14052 13628
rect 14052 13572 14056 13628
rect 13992 13568 14056 13572
rect 14072 13628 14136 13632
rect 14072 13572 14076 13628
rect 14076 13572 14132 13628
rect 14132 13572 14136 13628
rect 14072 13568 14136 13572
rect 20548 13628 20612 13632
rect 20548 13572 20552 13628
rect 20552 13572 20608 13628
rect 20608 13572 20612 13628
rect 20548 13568 20612 13572
rect 20628 13628 20692 13632
rect 20628 13572 20632 13628
rect 20632 13572 20688 13628
rect 20688 13572 20692 13628
rect 20628 13568 20692 13572
rect 20708 13628 20772 13632
rect 20708 13572 20712 13628
rect 20712 13572 20768 13628
rect 20768 13572 20772 13628
rect 20708 13568 20772 13572
rect 20788 13628 20852 13632
rect 20788 13572 20792 13628
rect 20792 13572 20848 13628
rect 20848 13572 20852 13628
rect 20788 13568 20852 13572
rect 27264 13628 27328 13632
rect 27264 13572 27268 13628
rect 27268 13572 27324 13628
rect 27324 13572 27328 13628
rect 27264 13568 27328 13572
rect 27344 13628 27408 13632
rect 27344 13572 27348 13628
rect 27348 13572 27404 13628
rect 27404 13572 27408 13628
rect 27344 13568 27408 13572
rect 27424 13628 27488 13632
rect 27424 13572 27428 13628
rect 27428 13572 27484 13628
rect 27484 13572 27488 13628
rect 27424 13568 27488 13572
rect 27504 13628 27568 13632
rect 27504 13572 27508 13628
rect 27508 13572 27564 13628
rect 27564 13572 27568 13628
rect 27504 13568 27568 13572
rect 3758 13084 3822 13088
rect 3758 13028 3762 13084
rect 3762 13028 3818 13084
rect 3818 13028 3822 13084
rect 3758 13024 3822 13028
rect 3838 13084 3902 13088
rect 3838 13028 3842 13084
rect 3842 13028 3898 13084
rect 3898 13028 3902 13084
rect 3838 13024 3902 13028
rect 3918 13084 3982 13088
rect 3918 13028 3922 13084
rect 3922 13028 3978 13084
rect 3978 13028 3982 13084
rect 3918 13024 3982 13028
rect 3998 13084 4062 13088
rect 3998 13028 4002 13084
rect 4002 13028 4058 13084
rect 4058 13028 4062 13084
rect 3998 13024 4062 13028
rect 10474 13084 10538 13088
rect 10474 13028 10478 13084
rect 10478 13028 10534 13084
rect 10534 13028 10538 13084
rect 10474 13024 10538 13028
rect 10554 13084 10618 13088
rect 10554 13028 10558 13084
rect 10558 13028 10614 13084
rect 10614 13028 10618 13084
rect 10554 13024 10618 13028
rect 10634 13084 10698 13088
rect 10634 13028 10638 13084
rect 10638 13028 10694 13084
rect 10694 13028 10698 13084
rect 10634 13024 10698 13028
rect 10714 13084 10778 13088
rect 10714 13028 10718 13084
rect 10718 13028 10774 13084
rect 10774 13028 10778 13084
rect 10714 13024 10778 13028
rect 17190 13084 17254 13088
rect 17190 13028 17194 13084
rect 17194 13028 17250 13084
rect 17250 13028 17254 13084
rect 17190 13024 17254 13028
rect 17270 13084 17334 13088
rect 17270 13028 17274 13084
rect 17274 13028 17330 13084
rect 17330 13028 17334 13084
rect 17270 13024 17334 13028
rect 17350 13084 17414 13088
rect 17350 13028 17354 13084
rect 17354 13028 17410 13084
rect 17410 13028 17414 13084
rect 17350 13024 17414 13028
rect 17430 13084 17494 13088
rect 17430 13028 17434 13084
rect 17434 13028 17490 13084
rect 17490 13028 17494 13084
rect 17430 13024 17494 13028
rect 23906 13084 23970 13088
rect 23906 13028 23910 13084
rect 23910 13028 23966 13084
rect 23966 13028 23970 13084
rect 23906 13024 23970 13028
rect 23986 13084 24050 13088
rect 23986 13028 23990 13084
rect 23990 13028 24046 13084
rect 24046 13028 24050 13084
rect 23986 13024 24050 13028
rect 24066 13084 24130 13088
rect 24066 13028 24070 13084
rect 24070 13028 24126 13084
rect 24126 13028 24130 13084
rect 24066 13024 24130 13028
rect 24146 13084 24210 13088
rect 24146 13028 24150 13084
rect 24150 13028 24206 13084
rect 24206 13028 24210 13084
rect 24146 13024 24210 13028
rect 21588 12608 21652 12612
rect 21588 12552 21638 12608
rect 21638 12552 21652 12608
rect 21588 12548 21652 12552
rect 7116 12540 7180 12544
rect 7116 12484 7120 12540
rect 7120 12484 7176 12540
rect 7176 12484 7180 12540
rect 7116 12480 7180 12484
rect 7196 12540 7260 12544
rect 7196 12484 7200 12540
rect 7200 12484 7256 12540
rect 7256 12484 7260 12540
rect 7196 12480 7260 12484
rect 7276 12540 7340 12544
rect 7276 12484 7280 12540
rect 7280 12484 7336 12540
rect 7336 12484 7340 12540
rect 7276 12480 7340 12484
rect 7356 12540 7420 12544
rect 7356 12484 7360 12540
rect 7360 12484 7416 12540
rect 7416 12484 7420 12540
rect 7356 12480 7420 12484
rect 13832 12540 13896 12544
rect 13832 12484 13836 12540
rect 13836 12484 13892 12540
rect 13892 12484 13896 12540
rect 13832 12480 13896 12484
rect 13912 12540 13976 12544
rect 13912 12484 13916 12540
rect 13916 12484 13972 12540
rect 13972 12484 13976 12540
rect 13912 12480 13976 12484
rect 13992 12540 14056 12544
rect 13992 12484 13996 12540
rect 13996 12484 14052 12540
rect 14052 12484 14056 12540
rect 13992 12480 14056 12484
rect 14072 12540 14136 12544
rect 14072 12484 14076 12540
rect 14076 12484 14132 12540
rect 14132 12484 14136 12540
rect 14072 12480 14136 12484
rect 20548 12540 20612 12544
rect 20548 12484 20552 12540
rect 20552 12484 20608 12540
rect 20608 12484 20612 12540
rect 20548 12480 20612 12484
rect 20628 12540 20692 12544
rect 20628 12484 20632 12540
rect 20632 12484 20688 12540
rect 20688 12484 20692 12540
rect 20628 12480 20692 12484
rect 20708 12540 20772 12544
rect 20708 12484 20712 12540
rect 20712 12484 20768 12540
rect 20768 12484 20772 12540
rect 20708 12480 20772 12484
rect 20788 12540 20852 12544
rect 20788 12484 20792 12540
rect 20792 12484 20848 12540
rect 20848 12484 20852 12540
rect 20788 12480 20852 12484
rect 27264 12540 27328 12544
rect 27264 12484 27268 12540
rect 27268 12484 27324 12540
rect 27324 12484 27328 12540
rect 27264 12480 27328 12484
rect 27344 12540 27408 12544
rect 27344 12484 27348 12540
rect 27348 12484 27404 12540
rect 27404 12484 27408 12540
rect 27344 12480 27408 12484
rect 27424 12540 27488 12544
rect 27424 12484 27428 12540
rect 27428 12484 27484 12540
rect 27484 12484 27488 12540
rect 27424 12480 27488 12484
rect 27504 12540 27568 12544
rect 27504 12484 27508 12540
rect 27508 12484 27564 12540
rect 27564 12484 27568 12540
rect 27504 12480 27568 12484
rect 26188 12336 26252 12340
rect 26188 12280 26202 12336
rect 26202 12280 26252 12336
rect 26188 12276 26252 12280
rect 3758 11996 3822 12000
rect 3758 11940 3762 11996
rect 3762 11940 3818 11996
rect 3818 11940 3822 11996
rect 3758 11936 3822 11940
rect 3838 11996 3902 12000
rect 3838 11940 3842 11996
rect 3842 11940 3898 11996
rect 3898 11940 3902 11996
rect 3838 11936 3902 11940
rect 3918 11996 3982 12000
rect 3918 11940 3922 11996
rect 3922 11940 3978 11996
rect 3978 11940 3982 11996
rect 3918 11936 3982 11940
rect 3998 11996 4062 12000
rect 3998 11940 4002 11996
rect 4002 11940 4058 11996
rect 4058 11940 4062 11996
rect 3998 11936 4062 11940
rect 10474 11996 10538 12000
rect 10474 11940 10478 11996
rect 10478 11940 10534 11996
rect 10534 11940 10538 11996
rect 10474 11936 10538 11940
rect 10554 11996 10618 12000
rect 10554 11940 10558 11996
rect 10558 11940 10614 11996
rect 10614 11940 10618 11996
rect 10554 11936 10618 11940
rect 10634 11996 10698 12000
rect 10634 11940 10638 11996
rect 10638 11940 10694 11996
rect 10694 11940 10698 11996
rect 10634 11936 10698 11940
rect 10714 11996 10778 12000
rect 10714 11940 10718 11996
rect 10718 11940 10774 11996
rect 10774 11940 10778 11996
rect 10714 11936 10778 11940
rect 17190 11996 17254 12000
rect 17190 11940 17194 11996
rect 17194 11940 17250 11996
rect 17250 11940 17254 11996
rect 17190 11936 17254 11940
rect 17270 11996 17334 12000
rect 17270 11940 17274 11996
rect 17274 11940 17330 11996
rect 17330 11940 17334 11996
rect 17270 11936 17334 11940
rect 17350 11996 17414 12000
rect 17350 11940 17354 11996
rect 17354 11940 17410 11996
rect 17410 11940 17414 11996
rect 17350 11936 17414 11940
rect 17430 11996 17494 12000
rect 17430 11940 17434 11996
rect 17434 11940 17490 11996
rect 17490 11940 17494 11996
rect 17430 11936 17494 11940
rect 23906 11996 23970 12000
rect 23906 11940 23910 11996
rect 23910 11940 23966 11996
rect 23966 11940 23970 11996
rect 23906 11936 23970 11940
rect 23986 11996 24050 12000
rect 23986 11940 23990 11996
rect 23990 11940 24046 11996
rect 24046 11940 24050 11996
rect 23986 11936 24050 11940
rect 24066 11996 24130 12000
rect 24066 11940 24070 11996
rect 24070 11940 24126 11996
rect 24126 11940 24130 11996
rect 24066 11936 24130 11940
rect 24146 11996 24210 12000
rect 24146 11940 24150 11996
rect 24150 11940 24206 11996
rect 24206 11940 24210 11996
rect 24146 11936 24210 11940
rect 7116 11452 7180 11456
rect 7116 11396 7120 11452
rect 7120 11396 7176 11452
rect 7176 11396 7180 11452
rect 7116 11392 7180 11396
rect 7196 11452 7260 11456
rect 7196 11396 7200 11452
rect 7200 11396 7256 11452
rect 7256 11396 7260 11452
rect 7196 11392 7260 11396
rect 7276 11452 7340 11456
rect 7276 11396 7280 11452
rect 7280 11396 7336 11452
rect 7336 11396 7340 11452
rect 7276 11392 7340 11396
rect 7356 11452 7420 11456
rect 7356 11396 7360 11452
rect 7360 11396 7416 11452
rect 7416 11396 7420 11452
rect 7356 11392 7420 11396
rect 13832 11452 13896 11456
rect 13832 11396 13836 11452
rect 13836 11396 13892 11452
rect 13892 11396 13896 11452
rect 13832 11392 13896 11396
rect 13912 11452 13976 11456
rect 13912 11396 13916 11452
rect 13916 11396 13972 11452
rect 13972 11396 13976 11452
rect 13912 11392 13976 11396
rect 13992 11452 14056 11456
rect 13992 11396 13996 11452
rect 13996 11396 14052 11452
rect 14052 11396 14056 11452
rect 13992 11392 14056 11396
rect 14072 11452 14136 11456
rect 14072 11396 14076 11452
rect 14076 11396 14132 11452
rect 14132 11396 14136 11452
rect 14072 11392 14136 11396
rect 20548 11452 20612 11456
rect 20548 11396 20552 11452
rect 20552 11396 20608 11452
rect 20608 11396 20612 11452
rect 20548 11392 20612 11396
rect 20628 11452 20692 11456
rect 20628 11396 20632 11452
rect 20632 11396 20688 11452
rect 20688 11396 20692 11452
rect 20628 11392 20692 11396
rect 20708 11452 20772 11456
rect 20708 11396 20712 11452
rect 20712 11396 20768 11452
rect 20768 11396 20772 11452
rect 20708 11392 20772 11396
rect 20788 11452 20852 11456
rect 20788 11396 20792 11452
rect 20792 11396 20848 11452
rect 20848 11396 20852 11452
rect 20788 11392 20852 11396
rect 27264 11452 27328 11456
rect 27264 11396 27268 11452
rect 27268 11396 27324 11452
rect 27324 11396 27328 11452
rect 27264 11392 27328 11396
rect 27344 11452 27408 11456
rect 27344 11396 27348 11452
rect 27348 11396 27404 11452
rect 27404 11396 27408 11452
rect 27344 11392 27408 11396
rect 27424 11452 27488 11456
rect 27424 11396 27428 11452
rect 27428 11396 27484 11452
rect 27484 11396 27488 11452
rect 27424 11392 27488 11396
rect 27504 11452 27568 11456
rect 27504 11396 27508 11452
rect 27508 11396 27564 11452
rect 27564 11396 27568 11452
rect 27504 11392 27568 11396
rect 16252 11188 16316 11252
rect 14780 11052 14844 11116
rect 3758 10908 3822 10912
rect 3758 10852 3762 10908
rect 3762 10852 3818 10908
rect 3818 10852 3822 10908
rect 3758 10848 3822 10852
rect 3838 10908 3902 10912
rect 3838 10852 3842 10908
rect 3842 10852 3898 10908
rect 3898 10852 3902 10908
rect 3838 10848 3902 10852
rect 3918 10908 3982 10912
rect 3918 10852 3922 10908
rect 3922 10852 3978 10908
rect 3978 10852 3982 10908
rect 3918 10848 3982 10852
rect 3998 10908 4062 10912
rect 3998 10852 4002 10908
rect 4002 10852 4058 10908
rect 4058 10852 4062 10908
rect 3998 10848 4062 10852
rect 10474 10908 10538 10912
rect 10474 10852 10478 10908
rect 10478 10852 10534 10908
rect 10534 10852 10538 10908
rect 10474 10848 10538 10852
rect 10554 10908 10618 10912
rect 10554 10852 10558 10908
rect 10558 10852 10614 10908
rect 10614 10852 10618 10908
rect 10554 10848 10618 10852
rect 10634 10908 10698 10912
rect 10634 10852 10638 10908
rect 10638 10852 10694 10908
rect 10694 10852 10698 10908
rect 10634 10848 10698 10852
rect 10714 10908 10778 10912
rect 10714 10852 10718 10908
rect 10718 10852 10774 10908
rect 10774 10852 10778 10908
rect 10714 10848 10778 10852
rect 17190 10908 17254 10912
rect 17190 10852 17194 10908
rect 17194 10852 17250 10908
rect 17250 10852 17254 10908
rect 17190 10848 17254 10852
rect 17270 10908 17334 10912
rect 17270 10852 17274 10908
rect 17274 10852 17330 10908
rect 17330 10852 17334 10908
rect 17270 10848 17334 10852
rect 17350 10908 17414 10912
rect 17350 10852 17354 10908
rect 17354 10852 17410 10908
rect 17410 10852 17414 10908
rect 17350 10848 17414 10852
rect 17430 10908 17494 10912
rect 17430 10852 17434 10908
rect 17434 10852 17490 10908
rect 17490 10852 17494 10908
rect 17430 10848 17494 10852
rect 23906 10908 23970 10912
rect 23906 10852 23910 10908
rect 23910 10852 23966 10908
rect 23966 10852 23970 10908
rect 23906 10848 23970 10852
rect 23986 10908 24050 10912
rect 23986 10852 23990 10908
rect 23990 10852 24046 10908
rect 24046 10852 24050 10908
rect 23986 10848 24050 10852
rect 24066 10908 24130 10912
rect 24066 10852 24070 10908
rect 24070 10852 24126 10908
rect 24126 10852 24130 10908
rect 24066 10848 24130 10852
rect 24146 10908 24210 10912
rect 24146 10852 24150 10908
rect 24150 10852 24206 10908
rect 24206 10852 24210 10908
rect 24146 10848 24210 10852
rect 7116 10364 7180 10368
rect 7116 10308 7120 10364
rect 7120 10308 7176 10364
rect 7176 10308 7180 10364
rect 7116 10304 7180 10308
rect 7196 10364 7260 10368
rect 7196 10308 7200 10364
rect 7200 10308 7256 10364
rect 7256 10308 7260 10364
rect 7196 10304 7260 10308
rect 7276 10364 7340 10368
rect 7276 10308 7280 10364
rect 7280 10308 7336 10364
rect 7336 10308 7340 10364
rect 7276 10304 7340 10308
rect 7356 10364 7420 10368
rect 7356 10308 7360 10364
rect 7360 10308 7416 10364
rect 7416 10308 7420 10364
rect 7356 10304 7420 10308
rect 13832 10364 13896 10368
rect 13832 10308 13836 10364
rect 13836 10308 13892 10364
rect 13892 10308 13896 10364
rect 13832 10304 13896 10308
rect 13912 10364 13976 10368
rect 13912 10308 13916 10364
rect 13916 10308 13972 10364
rect 13972 10308 13976 10364
rect 13912 10304 13976 10308
rect 13992 10364 14056 10368
rect 13992 10308 13996 10364
rect 13996 10308 14052 10364
rect 14052 10308 14056 10364
rect 13992 10304 14056 10308
rect 14072 10364 14136 10368
rect 14072 10308 14076 10364
rect 14076 10308 14132 10364
rect 14132 10308 14136 10364
rect 14072 10304 14136 10308
rect 20548 10364 20612 10368
rect 20548 10308 20552 10364
rect 20552 10308 20608 10364
rect 20608 10308 20612 10364
rect 20548 10304 20612 10308
rect 20628 10364 20692 10368
rect 20628 10308 20632 10364
rect 20632 10308 20688 10364
rect 20688 10308 20692 10364
rect 20628 10304 20692 10308
rect 20708 10364 20772 10368
rect 20708 10308 20712 10364
rect 20712 10308 20768 10364
rect 20768 10308 20772 10364
rect 20708 10304 20772 10308
rect 20788 10364 20852 10368
rect 20788 10308 20792 10364
rect 20792 10308 20848 10364
rect 20848 10308 20852 10364
rect 20788 10304 20852 10308
rect 27264 10364 27328 10368
rect 27264 10308 27268 10364
rect 27268 10308 27324 10364
rect 27324 10308 27328 10364
rect 27264 10304 27328 10308
rect 27344 10364 27408 10368
rect 27344 10308 27348 10364
rect 27348 10308 27404 10364
rect 27404 10308 27408 10364
rect 27344 10304 27408 10308
rect 27424 10364 27488 10368
rect 27424 10308 27428 10364
rect 27428 10308 27484 10364
rect 27484 10308 27488 10364
rect 27424 10304 27488 10308
rect 27504 10364 27568 10368
rect 27504 10308 27508 10364
rect 27508 10308 27564 10364
rect 27564 10308 27568 10364
rect 27504 10304 27568 10308
rect 3758 9820 3822 9824
rect 3758 9764 3762 9820
rect 3762 9764 3818 9820
rect 3818 9764 3822 9820
rect 3758 9760 3822 9764
rect 3838 9820 3902 9824
rect 3838 9764 3842 9820
rect 3842 9764 3898 9820
rect 3898 9764 3902 9820
rect 3838 9760 3902 9764
rect 3918 9820 3982 9824
rect 3918 9764 3922 9820
rect 3922 9764 3978 9820
rect 3978 9764 3982 9820
rect 3918 9760 3982 9764
rect 3998 9820 4062 9824
rect 3998 9764 4002 9820
rect 4002 9764 4058 9820
rect 4058 9764 4062 9820
rect 3998 9760 4062 9764
rect 10474 9820 10538 9824
rect 10474 9764 10478 9820
rect 10478 9764 10534 9820
rect 10534 9764 10538 9820
rect 10474 9760 10538 9764
rect 10554 9820 10618 9824
rect 10554 9764 10558 9820
rect 10558 9764 10614 9820
rect 10614 9764 10618 9820
rect 10554 9760 10618 9764
rect 10634 9820 10698 9824
rect 10634 9764 10638 9820
rect 10638 9764 10694 9820
rect 10694 9764 10698 9820
rect 10634 9760 10698 9764
rect 10714 9820 10778 9824
rect 10714 9764 10718 9820
rect 10718 9764 10774 9820
rect 10774 9764 10778 9820
rect 10714 9760 10778 9764
rect 17190 9820 17254 9824
rect 17190 9764 17194 9820
rect 17194 9764 17250 9820
rect 17250 9764 17254 9820
rect 17190 9760 17254 9764
rect 17270 9820 17334 9824
rect 17270 9764 17274 9820
rect 17274 9764 17330 9820
rect 17330 9764 17334 9820
rect 17270 9760 17334 9764
rect 17350 9820 17414 9824
rect 17350 9764 17354 9820
rect 17354 9764 17410 9820
rect 17410 9764 17414 9820
rect 17350 9760 17414 9764
rect 17430 9820 17494 9824
rect 17430 9764 17434 9820
rect 17434 9764 17490 9820
rect 17490 9764 17494 9820
rect 17430 9760 17494 9764
rect 23906 9820 23970 9824
rect 23906 9764 23910 9820
rect 23910 9764 23966 9820
rect 23966 9764 23970 9820
rect 23906 9760 23970 9764
rect 23986 9820 24050 9824
rect 23986 9764 23990 9820
rect 23990 9764 24046 9820
rect 24046 9764 24050 9820
rect 23986 9760 24050 9764
rect 24066 9820 24130 9824
rect 24066 9764 24070 9820
rect 24070 9764 24126 9820
rect 24126 9764 24130 9820
rect 24066 9760 24130 9764
rect 24146 9820 24210 9824
rect 24146 9764 24150 9820
rect 24150 9764 24206 9820
rect 24206 9764 24210 9820
rect 24146 9760 24210 9764
rect 11468 9556 11532 9620
rect 21588 9556 21652 9620
rect 26188 9420 26252 9484
rect 7116 9276 7180 9280
rect 7116 9220 7120 9276
rect 7120 9220 7176 9276
rect 7176 9220 7180 9276
rect 7116 9216 7180 9220
rect 7196 9276 7260 9280
rect 7196 9220 7200 9276
rect 7200 9220 7256 9276
rect 7256 9220 7260 9276
rect 7196 9216 7260 9220
rect 7276 9276 7340 9280
rect 7276 9220 7280 9276
rect 7280 9220 7336 9276
rect 7336 9220 7340 9276
rect 7276 9216 7340 9220
rect 7356 9276 7420 9280
rect 7356 9220 7360 9276
rect 7360 9220 7416 9276
rect 7416 9220 7420 9276
rect 7356 9216 7420 9220
rect 13832 9276 13896 9280
rect 13832 9220 13836 9276
rect 13836 9220 13892 9276
rect 13892 9220 13896 9276
rect 13832 9216 13896 9220
rect 13912 9276 13976 9280
rect 13912 9220 13916 9276
rect 13916 9220 13972 9276
rect 13972 9220 13976 9276
rect 13912 9216 13976 9220
rect 13992 9276 14056 9280
rect 13992 9220 13996 9276
rect 13996 9220 14052 9276
rect 14052 9220 14056 9276
rect 13992 9216 14056 9220
rect 14072 9276 14136 9280
rect 14072 9220 14076 9276
rect 14076 9220 14132 9276
rect 14132 9220 14136 9276
rect 14072 9216 14136 9220
rect 20548 9276 20612 9280
rect 20548 9220 20552 9276
rect 20552 9220 20608 9276
rect 20608 9220 20612 9276
rect 20548 9216 20612 9220
rect 20628 9276 20692 9280
rect 20628 9220 20632 9276
rect 20632 9220 20688 9276
rect 20688 9220 20692 9276
rect 20628 9216 20692 9220
rect 20708 9276 20772 9280
rect 20708 9220 20712 9276
rect 20712 9220 20768 9276
rect 20768 9220 20772 9276
rect 20708 9216 20772 9220
rect 20788 9276 20852 9280
rect 20788 9220 20792 9276
rect 20792 9220 20848 9276
rect 20848 9220 20852 9276
rect 20788 9216 20852 9220
rect 27264 9276 27328 9280
rect 27264 9220 27268 9276
rect 27268 9220 27324 9276
rect 27324 9220 27328 9276
rect 27264 9216 27328 9220
rect 27344 9276 27408 9280
rect 27344 9220 27348 9276
rect 27348 9220 27404 9276
rect 27404 9220 27408 9276
rect 27344 9216 27408 9220
rect 27424 9276 27488 9280
rect 27424 9220 27428 9276
rect 27428 9220 27484 9276
rect 27484 9220 27488 9276
rect 27424 9216 27488 9220
rect 27504 9276 27568 9280
rect 27504 9220 27508 9276
rect 27508 9220 27564 9276
rect 27564 9220 27568 9276
rect 27504 9216 27568 9220
rect 10180 9012 10244 9076
rect 3758 8732 3822 8736
rect 3758 8676 3762 8732
rect 3762 8676 3818 8732
rect 3818 8676 3822 8732
rect 3758 8672 3822 8676
rect 3838 8732 3902 8736
rect 3838 8676 3842 8732
rect 3842 8676 3898 8732
rect 3898 8676 3902 8732
rect 3838 8672 3902 8676
rect 3918 8732 3982 8736
rect 3918 8676 3922 8732
rect 3922 8676 3978 8732
rect 3978 8676 3982 8732
rect 3918 8672 3982 8676
rect 3998 8732 4062 8736
rect 3998 8676 4002 8732
rect 4002 8676 4058 8732
rect 4058 8676 4062 8732
rect 3998 8672 4062 8676
rect 10474 8732 10538 8736
rect 10474 8676 10478 8732
rect 10478 8676 10534 8732
rect 10534 8676 10538 8732
rect 10474 8672 10538 8676
rect 10554 8732 10618 8736
rect 10554 8676 10558 8732
rect 10558 8676 10614 8732
rect 10614 8676 10618 8732
rect 10554 8672 10618 8676
rect 10634 8732 10698 8736
rect 10634 8676 10638 8732
rect 10638 8676 10694 8732
rect 10694 8676 10698 8732
rect 10634 8672 10698 8676
rect 10714 8732 10778 8736
rect 10714 8676 10718 8732
rect 10718 8676 10774 8732
rect 10774 8676 10778 8732
rect 10714 8672 10778 8676
rect 17190 8732 17254 8736
rect 17190 8676 17194 8732
rect 17194 8676 17250 8732
rect 17250 8676 17254 8732
rect 17190 8672 17254 8676
rect 17270 8732 17334 8736
rect 17270 8676 17274 8732
rect 17274 8676 17330 8732
rect 17330 8676 17334 8732
rect 17270 8672 17334 8676
rect 17350 8732 17414 8736
rect 17350 8676 17354 8732
rect 17354 8676 17410 8732
rect 17410 8676 17414 8732
rect 17350 8672 17414 8676
rect 17430 8732 17494 8736
rect 17430 8676 17434 8732
rect 17434 8676 17490 8732
rect 17490 8676 17494 8732
rect 17430 8672 17494 8676
rect 23906 8732 23970 8736
rect 23906 8676 23910 8732
rect 23910 8676 23966 8732
rect 23966 8676 23970 8732
rect 23906 8672 23970 8676
rect 23986 8732 24050 8736
rect 23986 8676 23990 8732
rect 23990 8676 24046 8732
rect 24046 8676 24050 8732
rect 23986 8672 24050 8676
rect 24066 8732 24130 8736
rect 24066 8676 24070 8732
rect 24070 8676 24126 8732
rect 24126 8676 24130 8732
rect 24066 8672 24130 8676
rect 24146 8732 24210 8736
rect 24146 8676 24150 8732
rect 24150 8676 24206 8732
rect 24206 8676 24210 8732
rect 24146 8672 24210 8676
rect 7116 8188 7180 8192
rect 7116 8132 7120 8188
rect 7120 8132 7176 8188
rect 7176 8132 7180 8188
rect 7116 8128 7180 8132
rect 7196 8188 7260 8192
rect 7196 8132 7200 8188
rect 7200 8132 7256 8188
rect 7256 8132 7260 8188
rect 7196 8128 7260 8132
rect 7276 8188 7340 8192
rect 7276 8132 7280 8188
rect 7280 8132 7336 8188
rect 7336 8132 7340 8188
rect 7276 8128 7340 8132
rect 7356 8188 7420 8192
rect 7356 8132 7360 8188
rect 7360 8132 7416 8188
rect 7416 8132 7420 8188
rect 7356 8128 7420 8132
rect 13832 8188 13896 8192
rect 13832 8132 13836 8188
rect 13836 8132 13892 8188
rect 13892 8132 13896 8188
rect 13832 8128 13896 8132
rect 13912 8188 13976 8192
rect 13912 8132 13916 8188
rect 13916 8132 13972 8188
rect 13972 8132 13976 8188
rect 13912 8128 13976 8132
rect 13992 8188 14056 8192
rect 13992 8132 13996 8188
rect 13996 8132 14052 8188
rect 14052 8132 14056 8188
rect 13992 8128 14056 8132
rect 14072 8188 14136 8192
rect 14072 8132 14076 8188
rect 14076 8132 14132 8188
rect 14132 8132 14136 8188
rect 14072 8128 14136 8132
rect 20548 8188 20612 8192
rect 20548 8132 20552 8188
rect 20552 8132 20608 8188
rect 20608 8132 20612 8188
rect 20548 8128 20612 8132
rect 20628 8188 20692 8192
rect 20628 8132 20632 8188
rect 20632 8132 20688 8188
rect 20688 8132 20692 8188
rect 20628 8128 20692 8132
rect 20708 8188 20772 8192
rect 20708 8132 20712 8188
rect 20712 8132 20768 8188
rect 20768 8132 20772 8188
rect 20708 8128 20772 8132
rect 20788 8188 20852 8192
rect 20788 8132 20792 8188
rect 20792 8132 20848 8188
rect 20848 8132 20852 8188
rect 20788 8128 20852 8132
rect 27264 8188 27328 8192
rect 27264 8132 27268 8188
rect 27268 8132 27324 8188
rect 27324 8132 27328 8188
rect 27264 8128 27328 8132
rect 27344 8188 27408 8192
rect 27344 8132 27348 8188
rect 27348 8132 27404 8188
rect 27404 8132 27408 8188
rect 27344 8128 27408 8132
rect 27424 8188 27488 8192
rect 27424 8132 27428 8188
rect 27428 8132 27484 8188
rect 27484 8132 27488 8188
rect 27424 8128 27488 8132
rect 27504 8188 27568 8192
rect 27504 8132 27508 8188
rect 27508 8132 27564 8188
rect 27564 8132 27568 8188
rect 27504 8128 27568 8132
rect 3758 7644 3822 7648
rect 3758 7588 3762 7644
rect 3762 7588 3818 7644
rect 3818 7588 3822 7644
rect 3758 7584 3822 7588
rect 3838 7644 3902 7648
rect 3838 7588 3842 7644
rect 3842 7588 3898 7644
rect 3898 7588 3902 7644
rect 3838 7584 3902 7588
rect 3918 7644 3982 7648
rect 3918 7588 3922 7644
rect 3922 7588 3978 7644
rect 3978 7588 3982 7644
rect 3918 7584 3982 7588
rect 3998 7644 4062 7648
rect 3998 7588 4002 7644
rect 4002 7588 4058 7644
rect 4058 7588 4062 7644
rect 3998 7584 4062 7588
rect 10474 7644 10538 7648
rect 10474 7588 10478 7644
rect 10478 7588 10534 7644
rect 10534 7588 10538 7644
rect 10474 7584 10538 7588
rect 10554 7644 10618 7648
rect 10554 7588 10558 7644
rect 10558 7588 10614 7644
rect 10614 7588 10618 7644
rect 10554 7584 10618 7588
rect 10634 7644 10698 7648
rect 10634 7588 10638 7644
rect 10638 7588 10694 7644
rect 10694 7588 10698 7644
rect 10634 7584 10698 7588
rect 10714 7644 10778 7648
rect 10714 7588 10718 7644
rect 10718 7588 10774 7644
rect 10774 7588 10778 7644
rect 10714 7584 10778 7588
rect 17190 7644 17254 7648
rect 17190 7588 17194 7644
rect 17194 7588 17250 7644
rect 17250 7588 17254 7644
rect 17190 7584 17254 7588
rect 17270 7644 17334 7648
rect 17270 7588 17274 7644
rect 17274 7588 17330 7644
rect 17330 7588 17334 7644
rect 17270 7584 17334 7588
rect 17350 7644 17414 7648
rect 17350 7588 17354 7644
rect 17354 7588 17410 7644
rect 17410 7588 17414 7644
rect 17350 7584 17414 7588
rect 17430 7644 17494 7648
rect 17430 7588 17434 7644
rect 17434 7588 17490 7644
rect 17490 7588 17494 7644
rect 17430 7584 17494 7588
rect 23906 7644 23970 7648
rect 23906 7588 23910 7644
rect 23910 7588 23966 7644
rect 23966 7588 23970 7644
rect 23906 7584 23970 7588
rect 23986 7644 24050 7648
rect 23986 7588 23990 7644
rect 23990 7588 24046 7644
rect 24046 7588 24050 7644
rect 23986 7584 24050 7588
rect 24066 7644 24130 7648
rect 24066 7588 24070 7644
rect 24070 7588 24126 7644
rect 24126 7588 24130 7644
rect 24066 7584 24130 7588
rect 24146 7644 24210 7648
rect 24146 7588 24150 7644
rect 24150 7588 24206 7644
rect 24206 7588 24210 7644
rect 24146 7584 24210 7588
rect 21588 7380 21652 7444
rect 7116 7100 7180 7104
rect 7116 7044 7120 7100
rect 7120 7044 7176 7100
rect 7176 7044 7180 7100
rect 7116 7040 7180 7044
rect 7196 7100 7260 7104
rect 7196 7044 7200 7100
rect 7200 7044 7256 7100
rect 7256 7044 7260 7100
rect 7196 7040 7260 7044
rect 7276 7100 7340 7104
rect 7276 7044 7280 7100
rect 7280 7044 7336 7100
rect 7336 7044 7340 7100
rect 7276 7040 7340 7044
rect 7356 7100 7420 7104
rect 7356 7044 7360 7100
rect 7360 7044 7416 7100
rect 7416 7044 7420 7100
rect 7356 7040 7420 7044
rect 13832 7100 13896 7104
rect 13832 7044 13836 7100
rect 13836 7044 13892 7100
rect 13892 7044 13896 7100
rect 13832 7040 13896 7044
rect 13912 7100 13976 7104
rect 13912 7044 13916 7100
rect 13916 7044 13972 7100
rect 13972 7044 13976 7100
rect 13912 7040 13976 7044
rect 13992 7100 14056 7104
rect 13992 7044 13996 7100
rect 13996 7044 14052 7100
rect 14052 7044 14056 7100
rect 13992 7040 14056 7044
rect 14072 7100 14136 7104
rect 14072 7044 14076 7100
rect 14076 7044 14132 7100
rect 14132 7044 14136 7100
rect 14072 7040 14136 7044
rect 20548 7100 20612 7104
rect 20548 7044 20552 7100
rect 20552 7044 20608 7100
rect 20608 7044 20612 7100
rect 20548 7040 20612 7044
rect 20628 7100 20692 7104
rect 20628 7044 20632 7100
rect 20632 7044 20688 7100
rect 20688 7044 20692 7100
rect 20628 7040 20692 7044
rect 20708 7100 20772 7104
rect 20708 7044 20712 7100
rect 20712 7044 20768 7100
rect 20768 7044 20772 7100
rect 20708 7040 20772 7044
rect 20788 7100 20852 7104
rect 20788 7044 20792 7100
rect 20792 7044 20848 7100
rect 20848 7044 20852 7100
rect 20788 7040 20852 7044
rect 27264 7100 27328 7104
rect 27264 7044 27268 7100
rect 27268 7044 27324 7100
rect 27324 7044 27328 7100
rect 27264 7040 27328 7044
rect 27344 7100 27408 7104
rect 27344 7044 27348 7100
rect 27348 7044 27404 7100
rect 27404 7044 27408 7100
rect 27344 7040 27408 7044
rect 27424 7100 27488 7104
rect 27424 7044 27428 7100
rect 27428 7044 27484 7100
rect 27484 7044 27488 7100
rect 27424 7040 27488 7044
rect 27504 7100 27568 7104
rect 27504 7044 27508 7100
rect 27508 7044 27564 7100
rect 27564 7044 27568 7100
rect 27504 7040 27568 7044
rect 14412 6896 14476 6900
rect 14412 6840 14462 6896
rect 14462 6840 14476 6896
rect 14412 6836 14476 6840
rect 3758 6556 3822 6560
rect 3758 6500 3762 6556
rect 3762 6500 3818 6556
rect 3818 6500 3822 6556
rect 3758 6496 3822 6500
rect 3838 6556 3902 6560
rect 3838 6500 3842 6556
rect 3842 6500 3898 6556
rect 3898 6500 3902 6556
rect 3838 6496 3902 6500
rect 3918 6556 3982 6560
rect 3918 6500 3922 6556
rect 3922 6500 3978 6556
rect 3978 6500 3982 6556
rect 3918 6496 3982 6500
rect 3998 6556 4062 6560
rect 3998 6500 4002 6556
rect 4002 6500 4058 6556
rect 4058 6500 4062 6556
rect 3998 6496 4062 6500
rect 10474 6556 10538 6560
rect 10474 6500 10478 6556
rect 10478 6500 10534 6556
rect 10534 6500 10538 6556
rect 10474 6496 10538 6500
rect 10554 6556 10618 6560
rect 10554 6500 10558 6556
rect 10558 6500 10614 6556
rect 10614 6500 10618 6556
rect 10554 6496 10618 6500
rect 10634 6556 10698 6560
rect 10634 6500 10638 6556
rect 10638 6500 10694 6556
rect 10694 6500 10698 6556
rect 10634 6496 10698 6500
rect 10714 6556 10778 6560
rect 10714 6500 10718 6556
rect 10718 6500 10774 6556
rect 10774 6500 10778 6556
rect 10714 6496 10778 6500
rect 17190 6556 17254 6560
rect 17190 6500 17194 6556
rect 17194 6500 17250 6556
rect 17250 6500 17254 6556
rect 17190 6496 17254 6500
rect 17270 6556 17334 6560
rect 17270 6500 17274 6556
rect 17274 6500 17330 6556
rect 17330 6500 17334 6556
rect 17270 6496 17334 6500
rect 17350 6556 17414 6560
rect 17350 6500 17354 6556
rect 17354 6500 17410 6556
rect 17410 6500 17414 6556
rect 17350 6496 17414 6500
rect 17430 6556 17494 6560
rect 17430 6500 17434 6556
rect 17434 6500 17490 6556
rect 17490 6500 17494 6556
rect 17430 6496 17494 6500
rect 23906 6556 23970 6560
rect 23906 6500 23910 6556
rect 23910 6500 23966 6556
rect 23966 6500 23970 6556
rect 23906 6496 23970 6500
rect 23986 6556 24050 6560
rect 23986 6500 23990 6556
rect 23990 6500 24046 6556
rect 24046 6500 24050 6556
rect 23986 6496 24050 6500
rect 24066 6556 24130 6560
rect 24066 6500 24070 6556
rect 24070 6500 24126 6556
rect 24126 6500 24130 6556
rect 24066 6496 24130 6500
rect 24146 6556 24210 6560
rect 24146 6500 24150 6556
rect 24150 6500 24206 6556
rect 24206 6500 24210 6556
rect 24146 6496 24210 6500
rect 11468 6156 11532 6220
rect 7116 6012 7180 6016
rect 7116 5956 7120 6012
rect 7120 5956 7176 6012
rect 7176 5956 7180 6012
rect 7116 5952 7180 5956
rect 7196 6012 7260 6016
rect 7196 5956 7200 6012
rect 7200 5956 7256 6012
rect 7256 5956 7260 6012
rect 7196 5952 7260 5956
rect 7276 6012 7340 6016
rect 7276 5956 7280 6012
rect 7280 5956 7336 6012
rect 7336 5956 7340 6012
rect 7276 5952 7340 5956
rect 7356 6012 7420 6016
rect 7356 5956 7360 6012
rect 7360 5956 7416 6012
rect 7416 5956 7420 6012
rect 7356 5952 7420 5956
rect 13832 6012 13896 6016
rect 13832 5956 13836 6012
rect 13836 5956 13892 6012
rect 13892 5956 13896 6012
rect 13832 5952 13896 5956
rect 13912 6012 13976 6016
rect 13912 5956 13916 6012
rect 13916 5956 13972 6012
rect 13972 5956 13976 6012
rect 13912 5952 13976 5956
rect 13992 6012 14056 6016
rect 13992 5956 13996 6012
rect 13996 5956 14052 6012
rect 14052 5956 14056 6012
rect 13992 5952 14056 5956
rect 14072 6012 14136 6016
rect 14072 5956 14076 6012
rect 14076 5956 14132 6012
rect 14132 5956 14136 6012
rect 14072 5952 14136 5956
rect 20548 6012 20612 6016
rect 20548 5956 20552 6012
rect 20552 5956 20608 6012
rect 20608 5956 20612 6012
rect 20548 5952 20612 5956
rect 20628 6012 20692 6016
rect 20628 5956 20632 6012
rect 20632 5956 20688 6012
rect 20688 5956 20692 6012
rect 20628 5952 20692 5956
rect 20708 6012 20772 6016
rect 20708 5956 20712 6012
rect 20712 5956 20768 6012
rect 20768 5956 20772 6012
rect 20708 5952 20772 5956
rect 20788 6012 20852 6016
rect 20788 5956 20792 6012
rect 20792 5956 20848 6012
rect 20848 5956 20852 6012
rect 20788 5952 20852 5956
rect 27264 6012 27328 6016
rect 27264 5956 27268 6012
rect 27268 5956 27324 6012
rect 27324 5956 27328 6012
rect 27264 5952 27328 5956
rect 27344 6012 27408 6016
rect 27344 5956 27348 6012
rect 27348 5956 27404 6012
rect 27404 5956 27408 6012
rect 27344 5952 27408 5956
rect 27424 6012 27488 6016
rect 27424 5956 27428 6012
rect 27428 5956 27484 6012
rect 27484 5956 27488 6012
rect 27424 5952 27488 5956
rect 27504 6012 27568 6016
rect 27504 5956 27508 6012
rect 27508 5956 27564 6012
rect 27564 5956 27568 6012
rect 27504 5952 27568 5956
rect 3758 5468 3822 5472
rect 3758 5412 3762 5468
rect 3762 5412 3818 5468
rect 3818 5412 3822 5468
rect 3758 5408 3822 5412
rect 3838 5468 3902 5472
rect 3838 5412 3842 5468
rect 3842 5412 3898 5468
rect 3898 5412 3902 5468
rect 3838 5408 3902 5412
rect 3918 5468 3982 5472
rect 3918 5412 3922 5468
rect 3922 5412 3978 5468
rect 3978 5412 3982 5468
rect 3918 5408 3982 5412
rect 3998 5468 4062 5472
rect 3998 5412 4002 5468
rect 4002 5412 4058 5468
rect 4058 5412 4062 5468
rect 3998 5408 4062 5412
rect 10474 5468 10538 5472
rect 10474 5412 10478 5468
rect 10478 5412 10534 5468
rect 10534 5412 10538 5468
rect 10474 5408 10538 5412
rect 10554 5468 10618 5472
rect 10554 5412 10558 5468
rect 10558 5412 10614 5468
rect 10614 5412 10618 5468
rect 10554 5408 10618 5412
rect 10634 5468 10698 5472
rect 10634 5412 10638 5468
rect 10638 5412 10694 5468
rect 10694 5412 10698 5468
rect 10634 5408 10698 5412
rect 10714 5468 10778 5472
rect 10714 5412 10718 5468
rect 10718 5412 10774 5468
rect 10774 5412 10778 5468
rect 10714 5408 10778 5412
rect 17190 5468 17254 5472
rect 17190 5412 17194 5468
rect 17194 5412 17250 5468
rect 17250 5412 17254 5468
rect 17190 5408 17254 5412
rect 17270 5468 17334 5472
rect 17270 5412 17274 5468
rect 17274 5412 17330 5468
rect 17330 5412 17334 5468
rect 17270 5408 17334 5412
rect 17350 5468 17414 5472
rect 17350 5412 17354 5468
rect 17354 5412 17410 5468
rect 17410 5412 17414 5468
rect 17350 5408 17414 5412
rect 17430 5468 17494 5472
rect 17430 5412 17434 5468
rect 17434 5412 17490 5468
rect 17490 5412 17494 5468
rect 17430 5408 17494 5412
rect 23906 5468 23970 5472
rect 23906 5412 23910 5468
rect 23910 5412 23966 5468
rect 23966 5412 23970 5468
rect 23906 5408 23970 5412
rect 23986 5468 24050 5472
rect 23986 5412 23990 5468
rect 23990 5412 24046 5468
rect 24046 5412 24050 5468
rect 23986 5408 24050 5412
rect 24066 5468 24130 5472
rect 24066 5412 24070 5468
rect 24070 5412 24126 5468
rect 24126 5412 24130 5468
rect 24066 5408 24130 5412
rect 24146 5468 24210 5472
rect 24146 5412 24150 5468
rect 24150 5412 24206 5468
rect 24206 5412 24210 5468
rect 24146 5408 24210 5412
rect 11468 5264 11532 5268
rect 11468 5208 11482 5264
rect 11482 5208 11532 5264
rect 11468 5204 11532 5208
rect 7116 4924 7180 4928
rect 7116 4868 7120 4924
rect 7120 4868 7176 4924
rect 7176 4868 7180 4924
rect 7116 4864 7180 4868
rect 7196 4924 7260 4928
rect 7196 4868 7200 4924
rect 7200 4868 7256 4924
rect 7256 4868 7260 4924
rect 7196 4864 7260 4868
rect 7276 4924 7340 4928
rect 7276 4868 7280 4924
rect 7280 4868 7336 4924
rect 7336 4868 7340 4924
rect 7276 4864 7340 4868
rect 7356 4924 7420 4928
rect 7356 4868 7360 4924
rect 7360 4868 7416 4924
rect 7416 4868 7420 4924
rect 7356 4864 7420 4868
rect 13832 4924 13896 4928
rect 13832 4868 13836 4924
rect 13836 4868 13892 4924
rect 13892 4868 13896 4924
rect 13832 4864 13896 4868
rect 13912 4924 13976 4928
rect 13912 4868 13916 4924
rect 13916 4868 13972 4924
rect 13972 4868 13976 4924
rect 13912 4864 13976 4868
rect 13992 4924 14056 4928
rect 13992 4868 13996 4924
rect 13996 4868 14052 4924
rect 14052 4868 14056 4924
rect 13992 4864 14056 4868
rect 14072 4924 14136 4928
rect 14072 4868 14076 4924
rect 14076 4868 14132 4924
rect 14132 4868 14136 4924
rect 14072 4864 14136 4868
rect 20548 4924 20612 4928
rect 20548 4868 20552 4924
rect 20552 4868 20608 4924
rect 20608 4868 20612 4924
rect 20548 4864 20612 4868
rect 20628 4924 20692 4928
rect 20628 4868 20632 4924
rect 20632 4868 20688 4924
rect 20688 4868 20692 4924
rect 20628 4864 20692 4868
rect 20708 4924 20772 4928
rect 20708 4868 20712 4924
rect 20712 4868 20768 4924
rect 20768 4868 20772 4924
rect 20708 4864 20772 4868
rect 20788 4924 20852 4928
rect 20788 4868 20792 4924
rect 20792 4868 20848 4924
rect 20848 4868 20852 4924
rect 20788 4864 20852 4868
rect 27264 4924 27328 4928
rect 27264 4868 27268 4924
rect 27268 4868 27324 4924
rect 27324 4868 27328 4924
rect 27264 4864 27328 4868
rect 27344 4924 27408 4928
rect 27344 4868 27348 4924
rect 27348 4868 27404 4924
rect 27404 4868 27408 4924
rect 27344 4864 27408 4868
rect 27424 4924 27488 4928
rect 27424 4868 27428 4924
rect 27428 4868 27484 4924
rect 27484 4868 27488 4924
rect 27424 4864 27488 4868
rect 27504 4924 27568 4928
rect 27504 4868 27508 4924
rect 27508 4868 27564 4924
rect 27564 4868 27568 4924
rect 27504 4864 27568 4868
rect 3758 4380 3822 4384
rect 3758 4324 3762 4380
rect 3762 4324 3818 4380
rect 3818 4324 3822 4380
rect 3758 4320 3822 4324
rect 3838 4380 3902 4384
rect 3838 4324 3842 4380
rect 3842 4324 3898 4380
rect 3898 4324 3902 4380
rect 3838 4320 3902 4324
rect 3918 4380 3982 4384
rect 3918 4324 3922 4380
rect 3922 4324 3978 4380
rect 3978 4324 3982 4380
rect 3918 4320 3982 4324
rect 3998 4380 4062 4384
rect 3998 4324 4002 4380
rect 4002 4324 4058 4380
rect 4058 4324 4062 4380
rect 3998 4320 4062 4324
rect 10474 4380 10538 4384
rect 10474 4324 10478 4380
rect 10478 4324 10534 4380
rect 10534 4324 10538 4380
rect 10474 4320 10538 4324
rect 10554 4380 10618 4384
rect 10554 4324 10558 4380
rect 10558 4324 10614 4380
rect 10614 4324 10618 4380
rect 10554 4320 10618 4324
rect 10634 4380 10698 4384
rect 10634 4324 10638 4380
rect 10638 4324 10694 4380
rect 10694 4324 10698 4380
rect 10634 4320 10698 4324
rect 10714 4380 10778 4384
rect 10714 4324 10718 4380
rect 10718 4324 10774 4380
rect 10774 4324 10778 4380
rect 10714 4320 10778 4324
rect 17190 4380 17254 4384
rect 17190 4324 17194 4380
rect 17194 4324 17250 4380
rect 17250 4324 17254 4380
rect 17190 4320 17254 4324
rect 17270 4380 17334 4384
rect 17270 4324 17274 4380
rect 17274 4324 17330 4380
rect 17330 4324 17334 4380
rect 17270 4320 17334 4324
rect 17350 4380 17414 4384
rect 17350 4324 17354 4380
rect 17354 4324 17410 4380
rect 17410 4324 17414 4380
rect 17350 4320 17414 4324
rect 17430 4380 17494 4384
rect 17430 4324 17434 4380
rect 17434 4324 17490 4380
rect 17490 4324 17494 4380
rect 17430 4320 17494 4324
rect 23906 4380 23970 4384
rect 23906 4324 23910 4380
rect 23910 4324 23966 4380
rect 23966 4324 23970 4380
rect 23906 4320 23970 4324
rect 23986 4380 24050 4384
rect 23986 4324 23990 4380
rect 23990 4324 24046 4380
rect 24046 4324 24050 4380
rect 23986 4320 24050 4324
rect 24066 4380 24130 4384
rect 24066 4324 24070 4380
rect 24070 4324 24126 4380
rect 24126 4324 24130 4380
rect 24066 4320 24130 4324
rect 24146 4380 24210 4384
rect 24146 4324 24150 4380
rect 24150 4324 24206 4380
rect 24206 4324 24210 4380
rect 24146 4320 24210 4324
rect 7116 3836 7180 3840
rect 7116 3780 7120 3836
rect 7120 3780 7176 3836
rect 7176 3780 7180 3836
rect 7116 3776 7180 3780
rect 7196 3836 7260 3840
rect 7196 3780 7200 3836
rect 7200 3780 7256 3836
rect 7256 3780 7260 3836
rect 7196 3776 7260 3780
rect 7276 3836 7340 3840
rect 7276 3780 7280 3836
rect 7280 3780 7336 3836
rect 7336 3780 7340 3836
rect 7276 3776 7340 3780
rect 7356 3836 7420 3840
rect 7356 3780 7360 3836
rect 7360 3780 7416 3836
rect 7416 3780 7420 3836
rect 7356 3776 7420 3780
rect 13832 3836 13896 3840
rect 13832 3780 13836 3836
rect 13836 3780 13892 3836
rect 13892 3780 13896 3836
rect 13832 3776 13896 3780
rect 13912 3836 13976 3840
rect 13912 3780 13916 3836
rect 13916 3780 13972 3836
rect 13972 3780 13976 3836
rect 13912 3776 13976 3780
rect 13992 3836 14056 3840
rect 13992 3780 13996 3836
rect 13996 3780 14052 3836
rect 14052 3780 14056 3836
rect 13992 3776 14056 3780
rect 14072 3836 14136 3840
rect 14072 3780 14076 3836
rect 14076 3780 14132 3836
rect 14132 3780 14136 3836
rect 14072 3776 14136 3780
rect 20548 3836 20612 3840
rect 20548 3780 20552 3836
rect 20552 3780 20608 3836
rect 20608 3780 20612 3836
rect 20548 3776 20612 3780
rect 20628 3836 20692 3840
rect 20628 3780 20632 3836
rect 20632 3780 20688 3836
rect 20688 3780 20692 3836
rect 20628 3776 20692 3780
rect 20708 3836 20772 3840
rect 20708 3780 20712 3836
rect 20712 3780 20768 3836
rect 20768 3780 20772 3836
rect 20708 3776 20772 3780
rect 20788 3836 20852 3840
rect 20788 3780 20792 3836
rect 20792 3780 20848 3836
rect 20848 3780 20852 3836
rect 20788 3776 20852 3780
rect 27264 3836 27328 3840
rect 27264 3780 27268 3836
rect 27268 3780 27324 3836
rect 27324 3780 27328 3836
rect 27264 3776 27328 3780
rect 27344 3836 27408 3840
rect 27344 3780 27348 3836
rect 27348 3780 27404 3836
rect 27404 3780 27408 3836
rect 27344 3776 27408 3780
rect 27424 3836 27488 3840
rect 27424 3780 27428 3836
rect 27428 3780 27484 3836
rect 27484 3780 27488 3836
rect 27424 3776 27488 3780
rect 27504 3836 27568 3840
rect 27504 3780 27508 3836
rect 27508 3780 27564 3836
rect 27564 3780 27568 3836
rect 27504 3776 27568 3780
rect 3758 3292 3822 3296
rect 3758 3236 3762 3292
rect 3762 3236 3818 3292
rect 3818 3236 3822 3292
rect 3758 3232 3822 3236
rect 3838 3292 3902 3296
rect 3838 3236 3842 3292
rect 3842 3236 3898 3292
rect 3898 3236 3902 3292
rect 3838 3232 3902 3236
rect 3918 3292 3982 3296
rect 3918 3236 3922 3292
rect 3922 3236 3978 3292
rect 3978 3236 3982 3292
rect 3918 3232 3982 3236
rect 3998 3292 4062 3296
rect 3998 3236 4002 3292
rect 4002 3236 4058 3292
rect 4058 3236 4062 3292
rect 3998 3232 4062 3236
rect 10474 3292 10538 3296
rect 10474 3236 10478 3292
rect 10478 3236 10534 3292
rect 10534 3236 10538 3292
rect 10474 3232 10538 3236
rect 10554 3292 10618 3296
rect 10554 3236 10558 3292
rect 10558 3236 10614 3292
rect 10614 3236 10618 3292
rect 10554 3232 10618 3236
rect 10634 3292 10698 3296
rect 10634 3236 10638 3292
rect 10638 3236 10694 3292
rect 10694 3236 10698 3292
rect 10634 3232 10698 3236
rect 10714 3292 10778 3296
rect 10714 3236 10718 3292
rect 10718 3236 10774 3292
rect 10774 3236 10778 3292
rect 10714 3232 10778 3236
rect 17190 3292 17254 3296
rect 17190 3236 17194 3292
rect 17194 3236 17250 3292
rect 17250 3236 17254 3292
rect 17190 3232 17254 3236
rect 17270 3292 17334 3296
rect 17270 3236 17274 3292
rect 17274 3236 17330 3292
rect 17330 3236 17334 3292
rect 17270 3232 17334 3236
rect 17350 3292 17414 3296
rect 17350 3236 17354 3292
rect 17354 3236 17410 3292
rect 17410 3236 17414 3292
rect 17350 3232 17414 3236
rect 17430 3292 17494 3296
rect 17430 3236 17434 3292
rect 17434 3236 17490 3292
rect 17490 3236 17494 3292
rect 17430 3232 17494 3236
rect 23906 3292 23970 3296
rect 23906 3236 23910 3292
rect 23910 3236 23966 3292
rect 23966 3236 23970 3292
rect 23906 3232 23970 3236
rect 23986 3292 24050 3296
rect 23986 3236 23990 3292
rect 23990 3236 24046 3292
rect 24046 3236 24050 3292
rect 23986 3232 24050 3236
rect 24066 3292 24130 3296
rect 24066 3236 24070 3292
rect 24070 3236 24126 3292
rect 24126 3236 24130 3292
rect 24066 3232 24130 3236
rect 24146 3292 24210 3296
rect 24146 3236 24150 3292
rect 24150 3236 24206 3292
rect 24206 3236 24210 3292
rect 24146 3232 24210 3236
rect 7116 2748 7180 2752
rect 7116 2692 7120 2748
rect 7120 2692 7176 2748
rect 7176 2692 7180 2748
rect 7116 2688 7180 2692
rect 7196 2748 7260 2752
rect 7196 2692 7200 2748
rect 7200 2692 7256 2748
rect 7256 2692 7260 2748
rect 7196 2688 7260 2692
rect 7276 2748 7340 2752
rect 7276 2692 7280 2748
rect 7280 2692 7336 2748
rect 7336 2692 7340 2748
rect 7276 2688 7340 2692
rect 7356 2748 7420 2752
rect 7356 2692 7360 2748
rect 7360 2692 7416 2748
rect 7416 2692 7420 2748
rect 7356 2688 7420 2692
rect 13832 2748 13896 2752
rect 13832 2692 13836 2748
rect 13836 2692 13892 2748
rect 13892 2692 13896 2748
rect 13832 2688 13896 2692
rect 13912 2748 13976 2752
rect 13912 2692 13916 2748
rect 13916 2692 13972 2748
rect 13972 2692 13976 2748
rect 13912 2688 13976 2692
rect 13992 2748 14056 2752
rect 13992 2692 13996 2748
rect 13996 2692 14052 2748
rect 14052 2692 14056 2748
rect 13992 2688 14056 2692
rect 14072 2748 14136 2752
rect 14072 2692 14076 2748
rect 14076 2692 14132 2748
rect 14132 2692 14136 2748
rect 14072 2688 14136 2692
rect 20548 2748 20612 2752
rect 20548 2692 20552 2748
rect 20552 2692 20608 2748
rect 20608 2692 20612 2748
rect 20548 2688 20612 2692
rect 20628 2748 20692 2752
rect 20628 2692 20632 2748
rect 20632 2692 20688 2748
rect 20688 2692 20692 2748
rect 20628 2688 20692 2692
rect 20708 2748 20772 2752
rect 20708 2692 20712 2748
rect 20712 2692 20768 2748
rect 20768 2692 20772 2748
rect 20708 2688 20772 2692
rect 20788 2748 20852 2752
rect 20788 2692 20792 2748
rect 20792 2692 20848 2748
rect 20848 2692 20852 2748
rect 20788 2688 20852 2692
rect 27264 2748 27328 2752
rect 27264 2692 27268 2748
rect 27268 2692 27324 2748
rect 27324 2692 27328 2748
rect 27264 2688 27328 2692
rect 27344 2748 27408 2752
rect 27344 2692 27348 2748
rect 27348 2692 27404 2748
rect 27404 2692 27408 2748
rect 27344 2688 27408 2692
rect 27424 2748 27488 2752
rect 27424 2692 27428 2748
rect 27428 2692 27484 2748
rect 27484 2692 27488 2748
rect 27424 2688 27488 2692
rect 27504 2748 27568 2752
rect 27504 2692 27508 2748
rect 27508 2692 27564 2748
rect 27564 2692 27568 2748
rect 27504 2688 27568 2692
rect 14780 2620 14844 2684
rect 19380 2484 19444 2548
rect 20300 2348 20364 2412
rect 3758 2204 3822 2208
rect 3758 2148 3762 2204
rect 3762 2148 3818 2204
rect 3818 2148 3822 2204
rect 3758 2144 3822 2148
rect 3838 2204 3902 2208
rect 3838 2148 3842 2204
rect 3842 2148 3898 2204
rect 3898 2148 3902 2204
rect 3838 2144 3902 2148
rect 3918 2204 3982 2208
rect 3918 2148 3922 2204
rect 3922 2148 3978 2204
rect 3978 2148 3982 2204
rect 3918 2144 3982 2148
rect 3998 2204 4062 2208
rect 3998 2148 4002 2204
rect 4002 2148 4058 2204
rect 4058 2148 4062 2204
rect 3998 2144 4062 2148
rect 10474 2204 10538 2208
rect 10474 2148 10478 2204
rect 10478 2148 10534 2204
rect 10534 2148 10538 2204
rect 10474 2144 10538 2148
rect 10554 2204 10618 2208
rect 10554 2148 10558 2204
rect 10558 2148 10614 2204
rect 10614 2148 10618 2204
rect 10554 2144 10618 2148
rect 10634 2204 10698 2208
rect 10634 2148 10638 2204
rect 10638 2148 10694 2204
rect 10694 2148 10698 2204
rect 10634 2144 10698 2148
rect 10714 2204 10778 2208
rect 10714 2148 10718 2204
rect 10718 2148 10774 2204
rect 10774 2148 10778 2204
rect 10714 2144 10778 2148
rect 17190 2204 17254 2208
rect 17190 2148 17194 2204
rect 17194 2148 17250 2204
rect 17250 2148 17254 2204
rect 17190 2144 17254 2148
rect 17270 2204 17334 2208
rect 17270 2148 17274 2204
rect 17274 2148 17330 2204
rect 17330 2148 17334 2204
rect 17270 2144 17334 2148
rect 17350 2204 17414 2208
rect 17350 2148 17354 2204
rect 17354 2148 17410 2204
rect 17410 2148 17414 2204
rect 17350 2144 17414 2148
rect 17430 2204 17494 2208
rect 17430 2148 17434 2204
rect 17434 2148 17490 2204
rect 17490 2148 17494 2204
rect 17430 2144 17494 2148
rect 23906 2204 23970 2208
rect 23906 2148 23910 2204
rect 23910 2148 23966 2204
rect 23966 2148 23970 2204
rect 23906 2144 23970 2148
rect 23986 2204 24050 2208
rect 23986 2148 23990 2204
rect 23990 2148 24046 2204
rect 24046 2148 24050 2204
rect 23986 2144 24050 2148
rect 24066 2204 24130 2208
rect 24066 2148 24070 2204
rect 24070 2148 24126 2204
rect 24126 2148 24130 2204
rect 24066 2144 24130 2148
rect 24146 2204 24210 2208
rect 24146 2148 24150 2204
rect 24150 2148 24206 2204
rect 24206 2148 24210 2204
rect 24146 2144 24210 2148
rect 20300 2000 20364 2004
rect 20300 1944 20314 2000
rect 20314 1944 20364 2000
rect 20300 1940 20364 1944
rect 7116 1660 7180 1664
rect 7116 1604 7120 1660
rect 7120 1604 7176 1660
rect 7176 1604 7180 1660
rect 7116 1600 7180 1604
rect 7196 1660 7260 1664
rect 7196 1604 7200 1660
rect 7200 1604 7256 1660
rect 7256 1604 7260 1660
rect 7196 1600 7260 1604
rect 7276 1660 7340 1664
rect 7276 1604 7280 1660
rect 7280 1604 7336 1660
rect 7336 1604 7340 1660
rect 7276 1600 7340 1604
rect 7356 1660 7420 1664
rect 7356 1604 7360 1660
rect 7360 1604 7416 1660
rect 7416 1604 7420 1660
rect 7356 1600 7420 1604
rect 13832 1660 13896 1664
rect 13832 1604 13836 1660
rect 13836 1604 13892 1660
rect 13892 1604 13896 1660
rect 13832 1600 13896 1604
rect 13912 1660 13976 1664
rect 13912 1604 13916 1660
rect 13916 1604 13972 1660
rect 13972 1604 13976 1660
rect 13912 1600 13976 1604
rect 13992 1660 14056 1664
rect 13992 1604 13996 1660
rect 13996 1604 14052 1660
rect 14052 1604 14056 1660
rect 13992 1600 14056 1604
rect 14072 1660 14136 1664
rect 14072 1604 14076 1660
rect 14076 1604 14132 1660
rect 14132 1604 14136 1660
rect 14072 1600 14136 1604
rect 20548 1660 20612 1664
rect 20548 1604 20552 1660
rect 20552 1604 20608 1660
rect 20608 1604 20612 1660
rect 20548 1600 20612 1604
rect 20628 1660 20692 1664
rect 20628 1604 20632 1660
rect 20632 1604 20688 1660
rect 20688 1604 20692 1660
rect 20628 1600 20692 1604
rect 20708 1660 20772 1664
rect 20708 1604 20712 1660
rect 20712 1604 20768 1660
rect 20768 1604 20772 1660
rect 20708 1600 20772 1604
rect 20788 1660 20852 1664
rect 20788 1604 20792 1660
rect 20792 1604 20848 1660
rect 20848 1604 20852 1660
rect 20788 1600 20852 1604
rect 27264 1660 27328 1664
rect 27264 1604 27268 1660
rect 27268 1604 27324 1660
rect 27324 1604 27328 1660
rect 27264 1600 27328 1604
rect 27344 1660 27408 1664
rect 27344 1604 27348 1660
rect 27348 1604 27404 1660
rect 27404 1604 27408 1660
rect 27344 1600 27408 1604
rect 27424 1660 27488 1664
rect 27424 1604 27428 1660
rect 27428 1604 27484 1660
rect 27484 1604 27488 1660
rect 27424 1600 27488 1604
rect 27504 1660 27568 1664
rect 27504 1604 27508 1660
rect 27508 1604 27564 1660
rect 27564 1604 27568 1660
rect 27504 1600 27568 1604
rect 19380 1396 19444 1460
rect 3758 1116 3822 1120
rect 3758 1060 3762 1116
rect 3762 1060 3818 1116
rect 3818 1060 3822 1116
rect 3758 1056 3822 1060
rect 3838 1116 3902 1120
rect 3838 1060 3842 1116
rect 3842 1060 3898 1116
rect 3898 1060 3902 1116
rect 3838 1056 3902 1060
rect 3918 1116 3982 1120
rect 3918 1060 3922 1116
rect 3922 1060 3978 1116
rect 3978 1060 3982 1116
rect 3918 1056 3982 1060
rect 3998 1116 4062 1120
rect 3998 1060 4002 1116
rect 4002 1060 4058 1116
rect 4058 1060 4062 1116
rect 3998 1056 4062 1060
rect 10474 1116 10538 1120
rect 10474 1060 10478 1116
rect 10478 1060 10534 1116
rect 10534 1060 10538 1116
rect 10474 1056 10538 1060
rect 10554 1116 10618 1120
rect 10554 1060 10558 1116
rect 10558 1060 10614 1116
rect 10614 1060 10618 1116
rect 10554 1056 10618 1060
rect 10634 1116 10698 1120
rect 10634 1060 10638 1116
rect 10638 1060 10694 1116
rect 10694 1060 10698 1116
rect 10634 1056 10698 1060
rect 10714 1116 10778 1120
rect 10714 1060 10718 1116
rect 10718 1060 10774 1116
rect 10774 1060 10778 1116
rect 10714 1056 10778 1060
rect 17190 1116 17254 1120
rect 17190 1060 17194 1116
rect 17194 1060 17250 1116
rect 17250 1060 17254 1116
rect 17190 1056 17254 1060
rect 17270 1116 17334 1120
rect 17270 1060 17274 1116
rect 17274 1060 17330 1116
rect 17330 1060 17334 1116
rect 17270 1056 17334 1060
rect 17350 1116 17414 1120
rect 17350 1060 17354 1116
rect 17354 1060 17410 1116
rect 17410 1060 17414 1116
rect 17350 1056 17414 1060
rect 17430 1116 17494 1120
rect 17430 1060 17434 1116
rect 17434 1060 17490 1116
rect 17490 1060 17494 1116
rect 17430 1056 17494 1060
rect 23906 1116 23970 1120
rect 23906 1060 23910 1116
rect 23910 1060 23966 1116
rect 23966 1060 23970 1116
rect 23906 1056 23970 1060
rect 23986 1116 24050 1120
rect 23986 1060 23990 1116
rect 23990 1060 24046 1116
rect 24046 1060 24050 1116
rect 23986 1056 24050 1060
rect 24066 1116 24130 1120
rect 24066 1060 24070 1116
rect 24070 1060 24126 1116
rect 24126 1060 24130 1116
rect 24066 1056 24130 1060
rect 24146 1116 24210 1120
rect 24146 1060 24150 1116
rect 24150 1060 24206 1116
rect 24206 1060 24210 1116
rect 24146 1056 24210 1060
rect 16252 852 16316 916
rect 7116 572 7180 576
rect 7116 516 7120 572
rect 7120 516 7176 572
rect 7176 516 7180 572
rect 7116 512 7180 516
rect 7196 572 7260 576
rect 7196 516 7200 572
rect 7200 516 7256 572
rect 7256 516 7260 572
rect 7196 512 7260 516
rect 7276 572 7340 576
rect 7276 516 7280 572
rect 7280 516 7336 572
rect 7336 516 7340 572
rect 7276 512 7340 516
rect 7356 572 7420 576
rect 7356 516 7360 572
rect 7360 516 7416 572
rect 7416 516 7420 572
rect 7356 512 7420 516
rect 13832 572 13896 576
rect 13832 516 13836 572
rect 13836 516 13892 572
rect 13892 516 13896 572
rect 13832 512 13896 516
rect 13912 572 13976 576
rect 13912 516 13916 572
rect 13916 516 13972 572
rect 13972 516 13976 572
rect 13912 512 13976 516
rect 13992 572 14056 576
rect 13992 516 13996 572
rect 13996 516 14052 572
rect 14052 516 14056 572
rect 13992 512 14056 516
rect 14072 572 14136 576
rect 14072 516 14076 572
rect 14076 516 14132 572
rect 14132 516 14136 572
rect 14072 512 14136 516
rect 20548 572 20612 576
rect 20548 516 20552 572
rect 20552 516 20608 572
rect 20608 516 20612 572
rect 20548 512 20612 516
rect 20628 572 20692 576
rect 20628 516 20632 572
rect 20632 516 20688 572
rect 20688 516 20692 572
rect 20628 512 20692 516
rect 20708 572 20772 576
rect 20708 516 20712 572
rect 20712 516 20768 572
rect 20768 516 20772 572
rect 20708 512 20772 516
rect 20788 572 20852 576
rect 20788 516 20792 572
rect 20792 516 20848 572
rect 20848 516 20852 572
rect 20788 512 20852 516
rect 27264 572 27328 576
rect 27264 516 27268 572
rect 27268 516 27324 572
rect 27324 516 27328 572
rect 27264 512 27328 516
rect 27344 572 27408 576
rect 27344 516 27348 572
rect 27348 516 27404 572
rect 27404 516 27408 572
rect 27344 512 27408 516
rect 27424 572 27488 576
rect 27424 516 27428 572
rect 27428 516 27484 572
rect 27484 516 27488 572
rect 27424 512 27488 516
rect 27504 572 27568 576
rect 27504 516 27508 572
rect 27508 516 27564 572
rect 27564 516 27568 572
rect 27504 512 27568 516
<< metal4 >>
rect 3750 17440 4070 17456
rect 3750 17376 3758 17440
rect 3822 17376 3838 17440
rect 3902 17376 3918 17440
rect 3982 17376 3998 17440
rect 4062 17376 4070 17440
rect 3750 16352 4070 17376
rect 3750 16288 3758 16352
rect 3822 16288 3838 16352
rect 3902 16288 3918 16352
rect 3982 16288 3998 16352
rect 4062 16288 4070 16352
rect 3750 15264 4070 16288
rect 3750 15200 3758 15264
rect 3822 15200 3838 15264
rect 3902 15200 3918 15264
rect 3982 15200 3998 15264
rect 4062 15200 4070 15264
rect 3750 14176 4070 15200
rect 3750 14112 3758 14176
rect 3822 14112 3838 14176
rect 3902 14112 3918 14176
rect 3982 14112 3998 14176
rect 4062 14112 4070 14176
rect 3750 13088 4070 14112
rect 3750 13024 3758 13088
rect 3822 13024 3838 13088
rect 3902 13024 3918 13088
rect 3982 13024 3998 13088
rect 4062 13024 4070 13088
rect 3750 12000 4070 13024
rect 3750 11936 3758 12000
rect 3822 11936 3838 12000
rect 3902 11936 3918 12000
rect 3982 11936 3998 12000
rect 4062 11936 4070 12000
rect 3750 10912 4070 11936
rect 3750 10848 3758 10912
rect 3822 10848 3838 10912
rect 3902 10848 3918 10912
rect 3982 10848 3998 10912
rect 4062 10848 4070 10912
rect 3750 9824 4070 10848
rect 3750 9760 3758 9824
rect 3822 9760 3838 9824
rect 3902 9760 3918 9824
rect 3982 9760 3998 9824
rect 4062 9760 4070 9824
rect 3750 8736 4070 9760
rect 3750 8672 3758 8736
rect 3822 8672 3838 8736
rect 3902 8672 3918 8736
rect 3982 8672 3998 8736
rect 4062 8672 4070 8736
rect 3750 7648 4070 8672
rect 3750 7584 3758 7648
rect 3822 7584 3838 7648
rect 3902 7584 3918 7648
rect 3982 7584 3998 7648
rect 4062 7584 4070 7648
rect 3750 6560 4070 7584
rect 3750 6496 3758 6560
rect 3822 6496 3838 6560
rect 3902 6496 3918 6560
rect 3982 6496 3998 6560
rect 4062 6496 4070 6560
rect 3750 5472 4070 6496
rect 3750 5408 3758 5472
rect 3822 5408 3838 5472
rect 3902 5408 3918 5472
rect 3982 5408 3998 5472
rect 4062 5408 4070 5472
rect 3750 4384 4070 5408
rect 3750 4320 3758 4384
rect 3822 4320 3838 4384
rect 3902 4320 3918 4384
rect 3982 4320 3998 4384
rect 4062 4320 4070 4384
rect 3750 3296 4070 4320
rect 3750 3232 3758 3296
rect 3822 3232 3838 3296
rect 3902 3232 3918 3296
rect 3982 3232 3998 3296
rect 4062 3232 4070 3296
rect 3750 2208 4070 3232
rect 3750 2144 3758 2208
rect 3822 2144 3838 2208
rect 3902 2144 3918 2208
rect 3982 2144 3998 2208
rect 4062 2144 4070 2208
rect 3750 1120 4070 2144
rect 3750 1056 3758 1120
rect 3822 1056 3838 1120
rect 3902 1056 3918 1120
rect 3982 1056 3998 1120
rect 4062 1056 4070 1120
rect 3750 496 4070 1056
rect 7108 16896 7428 17456
rect 7108 16832 7116 16896
rect 7180 16832 7196 16896
rect 7260 16832 7276 16896
rect 7340 16832 7356 16896
rect 7420 16832 7428 16896
rect 7108 15808 7428 16832
rect 7108 15744 7116 15808
rect 7180 15744 7196 15808
rect 7260 15744 7276 15808
rect 7340 15744 7356 15808
rect 7420 15744 7428 15808
rect 7108 14720 7428 15744
rect 10466 17440 10786 17456
rect 10466 17376 10474 17440
rect 10538 17376 10554 17440
rect 10618 17376 10634 17440
rect 10698 17376 10714 17440
rect 10778 17376 10786 17440
rect 10466 16352 10786 17376
rect 10466 16288 10474 16352
rect 10538 16288 10554 16352
rect 10618 16288 10634 16352
rect 10698 16288 10714 16352
rect 10778 16288 10786 16352
rect 10179 15332 10245 15333
rect 10179 15268 10180 15332
rect 10244 15268 10245 15332
rect 10179 15267 10245 15268
rect 7108 14656 7116 14720
rect 7180 14656 7196 14720
rect 7260 14656 7276 14720
rect 7340 14656 7356 14720
rect 7420 14656 7428 14720
rect 7108 13632 7428 14656
rect 7108 13568 7116 13632
rect 7180 13568 7196 13632
rect 7260 13568 7276 13632
rect 7340 13568 7356 13632
rect 7420 13568 7428 13632
rect 7108 12544 7428 13568
rect 7108 12480 7116 12544
rect 7180 12480 7196 12544
rect 7260 12480 7276 12544
rect 7340 12480 7356 12544
rect 7420 12480 7428 12544
rect 7108 11456 7428 12480
rect 7108 11392 7116 11456
rect 7180 11392 7196 11456
rect 7260 11392 7276 11456
rect 7340 11392 7356 11456
rect 7420 11392 7428 11456
rect 7108 10368 7428 11392
rect 7108 10304 7116 10368
rect 7180 10304 7196 10368
rect 7260 10304 7276 10368
rect 7340 10304 7356 10368
rect 7420 10304 7428 10368
rect 7108 9280 7428 10304
rect 7108 9216 7116 9280
rect 7180 9216 7196 9280
rect 7260 9216 7276 9280
rect 7340 9216 7356 9280
rect 7420 9216 7428 9280
rect 7108 8192 7428 9216
rect 10182 9077 10242 15267
rect 10466 15264 10786 16288
rect 10466 15200 10474 15264
rect 10538 15200 10554 15264
rect 10618 15200 10634 15264
rect 10698 15200 10714 15264
rect 10778 15200 10786 15264
rect 10466 14176 10786 15200
rect 10466 14112 10474 14176
rect 10538 14112 10554 14176
rect 10618 14112 10634 14176
rect 10698 14112 10714 14176
rect 10778 14112 10786 14176
rect 10466 13088 10786 14112
rect 10466 13024 10474 13088
rect 10538 13024 10554 13088
rect 10618 13024 10634 13088
rect 10698 13024 10714 13088
rect 10778 13024 10786 13088
rect 10466 12000 10786 13024
rect 10466 11936 10474 12000
rect 10538 11936 10554 12000
rect 10618 11936 10634 12000
rect 10698 11936 10714 12000
rect 10778 11936 10786 12000
rect 10466 10912 10786 11936
rect 10466 10848 10474 10912
rect 10538 10848 10554 10912
rect 10618 10848 10634 10912
rect 10698 10848 10714 10912
rect 10778 10848 10786 10912
rect 10466 9824 10786 10848
rect 10466 9760 10474 9824
rect 10538 9760 10554 9824
rect 10618 9760 10634 9824
rect 10698 9760 10714 9824
rect 10778 9760 10786 9824
rect 10179 9076 10245 9077
rect 10179 9012 10180 9076
rect 10244 9012 10245 9076
rect 10179 9011 10245 9012
rect 7108 8128 7116 8192
rect 7180 8128 7196 8192
rect 7260 8128 7276 8192
rect 7340 8128 7356 8192
rect 7420 8128 7428 8192
rect 7108 7104 7428 8128
rect 7108 7040 7116 7104
rect 7180 7040 7196 7104
rect 7260 7040 7276 7104
rect 7340 7040 7356 7104
rect 7420 7040 7428 7104
rect 7108 6016 7428 7040
rect 7108 5952 7116 6016
rect 7180 5952 7196 6016
rect 7260 5952 7276 6016
rect 7340 5952 7356 6016
rect 7420 5952 7428 6016
rect 7108 4928 7428 5952
rect 7108 4864 7116 4928
rect 7180 4864 7196 4928
rect 7260 4864 7276 4928
rect 7340 4864 7356 4928
rect 7420 4864 7428 4928
rect 7108 3840 7428 4864
rect 7108 3776 7116 3840
rect 7180 3776 7196 3840
rect 7260 3776 7276 3840
rect 7340 3776 7356 3840
rect 7420 3776 7428 3840
rect 7108 2752 7428 3776
rect 7108 2688 7116 2752
rect 7180 2688 7196 2752
rect 7260 2688 7276 2752
rect 7340 2688 7356 2752
rect 7420 2688 7428 2752
rect 7108 1664 7428 2688
rect 7108 1600 7116 1664
rect 7180 1600 7196 1664
rect 7260 1600 7276 1664
rect 7340 1600 7356 1664
rect 7420 1600 7428 1664
rect 7108 576 7428 1600
rect 7108 512 7116 576
rect 7180 512 7196 576
rect 7260 512 7276 576
rect 7340 512 7356 576
rect 7420 512 7428 576
rect 7108 496 7428 512
rect 10466 8736 10786 9760
rect 13824 16896 14144 17456
rect 13824 16832 13832 16896
rect 13896 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14144 16896
rect 13824 15808 14144 16832
rect 17182 17440 17502 17456
rect 17182 17376 17190 17440
rect 17254 17376 17270 17440
rect 17334 17376 17350 17440
rect 17414 17376 17430 17440
rect 17494 17376 17502 17440
rect 14411 16692 14477 16693
rect 14411 16628 14412 16692
rect 14476 16628 14477 16692
rect 14411 16627 14477 16628
rect 13824 15744 13832 15808
rect 13896 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14144 15808
rect 13824 14720 14144 15744
rect 13824 14656 13832 14720
rect 13896 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14144 14720
rect 13824 13632 14144 14656
rect 13824 13568 13832 13632
rect 13896 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14144 13632
rect 13824 12544 14144 13568
rect 13824 12480 13832 12544
rect 13896 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14144 12544
rect 13824 11456 14144 12480
rect 13824 11392 13832 11456
rect 13896 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14144 11456
rect 13824 10368 14144 11392
rect 13824 10304 13832 10368
rect 13896 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14144 10368
rect 11467 9620 11533 9621
rect 11467 9556 11468 9620
rect 11532 9556 11533 9620
rect 11467 9555 11533 9556
rect 10466 8672 10474 8736
rect 10538 8672 10554 8736
rect 10618 8672 10634 8736
rect 10698 8672 10714 8736
rect 10778 8672 10786 8736
rect 10466 7648 10786 8672
rect 10466 7584 10474 7648
rect 10538 7584 10554 7648
rect 10618 7584 10634 7648
rect 10698 7584 10714 7648
rect 10778 7584 10786 7648
rect 10466 6560 10786 7584
rect 10466 6496 10474 6560
rect 10538 6496 10554 6560
rect 10618 6496 10634 6560
rect 10698 6496 10714 6560
rect 10778 6496 10786 6560
rect 10466 5472 10786 6496
rect 11470 6221 11530 9555
rect 13824 9280 14144 10304
rect 13824 9216 13832 9280
rect 13896 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14144 9280
rect 13824 8192 14144 9216
rect 13824 8128 13832 8192
rect 13896 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14144 8192
rect 13824 7104 14144 8128
rect 13824 7040 13832 7104
rect 13896 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14144 7104
rect 11467 6220 11533 6221
rect 11467 6156 11468 6220
rect 11532 6156 11533 6220
rect 11467 6155 11533 6156
rect 10466 5408 10474 5472
rect 10538 5408 10554 5472
rect 10618 5408 10634 5472
rect 10698 5408 10714 5472
rect 10778 5408 10786 5472
rect 10466 4384 10786 5408
rect 11470 5269 11530 6155
rect 13824 6016 14144 7040
rect 14414 6901 14474 16627
rect 17182 16352 17502 17376
rect 20540 16896 20860 17456
rect 20540 16832 20548 16896
rect 20612 16832 20628 16896
rect 20692 16832 20708 16896
rect 20772 16832 20788 16896
rect 20852 16832 20860 16896
rect 19379 16692 19445 16693
rect 19379 16628 19380 16692
rect 19444 16628 19445 16692
rect 19379 16627 19445 16628
rect 20299 16692 20365 16693
rect 20299 16628 20300 16692
rect 20364 16628 20365 16692
rect 20299 16627 20365 16628
rect 17182 16288 17190 16352
rect 17254 16288 17270 16352
rect 17334 16288 17350 16352
rect 17414 16288 17430 16352
rect 17494 16288 17502 16352
rect 17182 15264 17502 16288
rect 17182 15200 17190 15264
rect 17254 15200 17270 15264
rect 17334 15200 17350 15264
rect 17414 15200 17430 15264
rect 17494 15200 17502 15264
rect 17182 14176 17502 15200
rect 17182 14112 17190 14176
rect 17254 14112 17270 14176
rect 17334 14112 17350 14176
rect 17414 14112 17430 14176
rect 17494 14112 17502 14176
rect 17182 13088 17502 14112
rect 17182 13024 17190 13088
rect 17254 13024 17270 13088
rect 17334 13024 17350 13088
rect 17414 13024 17430 13088
rect 17494 13024 17502 13088
rect 17182 12000 17502 13024
rect 17182 11936 17190 12000
rect 17254 11936 17270 12000
rect 17334 11936 17350 12000
rect 17414 11936 17430 12000
rect 17494 11936 17502 12000
rect 16251 11252 16317 11253
rect 16251 11188 16252 11252
rect 16316 11188 16317 11252
rect 16251 11187 16317 11188
rect 14779 11116 14845 11117
rect 14779 11052 14780 11116
rect 14844 11052 14845 11116
rect 14779 11051 14845 11052
rect 14411 6900 14477 6901
rect 14411 6836 14412 6900
rect 14476 6836 14477 6900
rect 14411 6835 14477 6836
rect 13824 5952 13832 6016
rect 13896 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14144 6016
rect 11467 5268 11533 5269
rect 11467 5204 11468 5268
rect 11532 5204 11533 5268
rect 11467 5203 11533 5204
rect 10466 4320 10474 4384
rect 10538 4320 10554 4384
rect 10618 4320 10634 4384
rect 10698 4320 10714 4384
rect 10778 4320 10786 4384
rect 10466 3296 10786 4320
rect 10466 3232 10474 3296
rect 10538 3232 10554 3296
rect 10618 3232 10634 3296
rect 10698 3232 10714 3296
rect 10778 3232 10786 3296
rect 10466 2208 10786 3232
rect 10466 2144 10474 2208
rect 10538 2144 10554 2208
rect 10618 2144 10634 2208
rect 10698 2144 10714 2208
rect 10778 2144 10786 2208
rect 10466 1120 10786 2144
rect 10466 1056 10474 1120
rect 10538 1056 10554 1120
rect 10618 1056 10634 1120
rect 10698 1056 10714 1120
rect 10778 1056 10786 1120
rect 10466 496 10786 1056
rect 13824 4928 14144 5952
rect 13824 4864 13832 4928
rect 13896 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14144 4928
rect 13824 3840 14144 4864
rect 13824 3776 13832 3840
rect 13896 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14144 3840
rect 13824 2752 14144 3776
rect 13824 2688 13832 2752
rect 13896 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14144 2752
rect 13824 1664 14144 2688
rect 14782 2685 14842 11051
rect 14779 2684 14845 2685
rect 14779 2620 14780 2684
rect 14844 2620 14845 2684
rect 14779 2619 14845 2620
rect 13824 1600 13832 1664
rect 13896 1600 13912 1664
rect 13976 1600 13992 1664
rect 14056 1600 14072 1664
rect 14136 1600 14144 1664
rect 13824 576 14144 1600
rect 16254 917 16314 11187
rect 17182 10912 17502 11936
rect 17182 10848 17190 10912
rect 17254 10848 17270 10912
rect 17334 10848 17350 10912
rect 17414 10848 17430 10912
rect 17494 10848 17502 10912
rect 17182 9824 17502 10848
rect 17182 9760 17190 9824
rect 17254 9760 17270 9824
rect 17334 9760 17350 9824
rect 17414 9760 17430 9824
rect 17494 9760 17502 9824
rect 17182 8736 17502 9760
rect 17182 8672 17190 8736
rect 17254 8672 17270 8736
rect 17334 8672 17350 8736
rect 17414 8672 17430 8736
rect 17494 8672 17502 8736
rect 17182 7648 17502 8672
rect 17182 7584 17190 7648
rect 17254 7584 17270 7648
rect 17334 7584 17350 7648
rect 17414 7584 17430 7648
rect 17494 7584 17502 7648
rect 17182 6560 17502 7584
rect 17182 6496 17190 6560
rect 17254 6496 17270 6560
rect 17334 6496 17350 6560
rect 17414 6496 17430 6560
rect 17494 6496 17502 6560
rect 17182 5472 17502 6496
rect 17182 5408 17190 5472
rect 17254 5408 17270 5472
rect 17334 5408 17350 5472
rect 17414 5408 17430 5472
rect 17494 5408 17502 5472
rect 17182 4384 17502 5408
rect 17182 4320 17190 4384
rect 17254 4320 17270 4384
rect 17334 4320 17350 4384
rect 17414 4320 17430 4384
rect 17494 4320 17502 4384
rect 17182 3296 17502 4320
rect 17182 3232 17190 3296
rect 17254 3232 17270 3296
rect 17334 3232 17350 3296
rect 17414 3232 17430 3296
rect 17494 3232 17502 3296
rect 17182 2208 17502 3232
rect 19382 2549 19442 16627
rect 19379 2548 19445 2549
rect 19379 2484 19380 2548
rect 19444 2484 19445 2548
rect 19379 2483 19445 2484
rect 17182 2144 17190 2208
rect 17254 2144 17270 2208
rect 17334 2144 17350 2208
rect 17414 2144 17430 2208
rect 17494 2144 17502 2208
rect 17182 1120 17502 2144
rect 19382 1461 19442 2483
rect 20302 2413 20362 16627
rect 20540 15808 20860 16832
rect 20540 15744 20548 15808
rect 20612 15744 20628 15808
rect 20692 15744 20708 15808
rect 20772 15744 20788 15808
rect 20852 15744 20860 15808
rect 20540 14720 20860 15744
rect 20540 14656 20548 14720
rect 20612 14656 20628 14720
rect 20692 14656 20708 14720
rect 20772 14656 20788 14720
rect 20852 14656 20860 14720
rect 20540 13632 20860 14656
rect 20540 13568 20548 13632
rect 20612 13568 20628 13632
rect 20692 13568 20708 13632
rect 20772 13568 20788 13632
rect 20852 13568 20860 13632
rect 20540 12544 20860 13568
rect 23898 17440 24218 17456
rect 23898 17376 23906 17440
rect 23970 17376 23986 17440
rect 24050 17376 24066 17440
rect 24130 17376 24146 17440
rect 24210 17376 24218 17440
rect 23898 16352 24218 17376
rect 23898 16288 23906 16352
rect 23970 16288 23986 16352
rect 24050 16288 24066 16352
rect 24130 16288 24146 16352
rect 24210 16288 24218 16352
rect 23898 15264 24218 16288
rect 23898 15200 23906 15264
rect 23970 15200 23986 15264
rect 24050 15200 24066 15264
rect 24130 15200 24146 15264
rect 24210 15200 24218 15264
rect 23898 14176 24218 15200
rect 23898 14112 23906 14176
rect 23970 14112 23986 14176
rect 24050 14112 24066 14176
rect 24130 14112 24146 14176
rect 24210 14112 24218 14176
rect 23898 13088 24218 14112
rect 23898 13024 23906 13088
rect 23970 13024 23986 13088
rect 24050 13024 24066 13088
rect 24130 13024 24146 13088
rect 24210 13024 24218 13088
rect 21587 12612 21653 12613
rect 21587 12548 21588 12612
rect 21652 12548 21653 12612
rect 21587 12547 21653 12548
rect 20540 12480 20548 12544
rect 20612 12480 20628 12544
rect 20692 12480 20708 12544
rect 20772 12480 20788 12544
rect 20852 12480 20860 12544
rect 20540 11456 20860 12480
rect 20540 11392 20548 11456
rect 20612 11392 20628 11456
rect 20692 11392 20708 11456
rect 20772 11392 20788 11456
rect 20852 11392 20860 11456
rect 20540 10368 20860 11392
rect 20540 10304 20548 10368
rect 20612 10304 20628 10368
rect 20692 10304 20708 10368
rect 20772 10304 20788 10368
rect 20852 10304 20860 10368
rect 20540 9280 20860 10304
rect 21590 9621 21650 12547
rect 23898 12000 24218 13024
rect 27256 16896 27576 17456
rect 27256 16832 27264 16896
rect 27328 16832 27344 16896
rect 27408 16832 27424 16896
rect 27488 16832 27504 16896
rect 27568 16832 27576 16896
rect 27256 15808 27576 16832
rect 27256 15744 27264 15808
rect 27328 15744 27344 15808
rect 27408 15744 27424 15808
rect 27488 15744 27504 15808
rect 27568 15744 27576 15808
rect 27256 14720 27576 15744
rect 27256 14656 27264 14720
rect 27328 14656 27344 14720
rect 27408 14656 27424 14720
rect 27488 14656 27504 14720
rect 27568 14656 27576 14720
rect 27256 13632 27576 14656
rect 27256 13568 27264 13632
rect 27328 13568 27344 13632
rect 27408 13568 27424 13632
rect 27488 13568 27504 13632
rect 27568 13568 27576 13632
rect 27256 12544 27576 13568
rect 27256 12480 27264 12544
rect 27328 12480 27344 12544
rect 27408 12480 27424 12544
rect 27488 12480 27504 12544
rect 27568 12480 27576 12544
rect 26187 12340 26253 12341
rect 26187 12276 26188 12340
rect 26252 12276 26253 12340
rect 26187 12275 26253 12276
rect 23898 11936 23906 12000
rect 23970 11936 23986 12000
rect 24050 11936 24066 12000
rect 24130 11936 24146 12000
rect 24210 11936 24218 12000
rect 23898 10912 24218 11936
rect 23898 10848 23906 10912
rect 23970 10848 23986 10912
rect 24050 10848 24066 10912
rect 24130 10848 24146 10912
rect 24210 10848 24218 10912
rect 23898 9824 24218 10848
rect 23898 9760 23906 9824
rect 23970 9760 23986 9824
rect 24050 9760 24066 9824
rect 24130 9760 24146 9824
rect 24210 9760 24218 9824
rect 21587 9620 21653 9621
rect 21587 9556 21588 9620
rect 21652 9556 21653 9620
rect 21587 9555 21653 9556
rect 20540 9216 20548 9280
rect 20612 9216 20628 9280
rect 20692 9216 20708 9280
rect 20772 9216 20788 9280
rect 20852 9216 20860 9280
rect 20540 8192 20860 9216
rect 20540 8128 20548 8192
rect 20612 8128 20628 8192
rect 20692 8128 20708 8192
rect 20772 8128 20788 8192
rect 20852 8128 20860 8192
rect 20540 7104 20860 8128
rect 21590 7445 21650 9555
rect 23898 8736 24218 9760
rect 26190 9485 26250 12275
rect 27256 11456 27576 12480
rect 27256 11392 27264 11456
rect 27328 11392 27344 11456
rect 27408 11392 27424 11456
rect 27488 11392 27504 11456
rect 27568 11392 27576 11456
rect 27256 10368 27576 11392
rect 27256 10304 27264 10368
rect 27328 10304 27344 10368
rect 27408 10304 27424 10368
rect 27488 10304 27504 10368
rect 27568 10304 27576 10368
rect 26187 9484 26253 9485
rect 26187 9420 26188 9484
rect 26252 9420 26253 9484
rect 26187 9419 26253 9420
rect 23898 8672 23906 8736
rect 23970 8672 23986 8736
rect 24050 8672 24066 8736
rect 24130 8672 24146 8736
rect 24210 8672 24218 8736
rect 23898 7648 24218 8672
rect 23898 7584 23906 7648
rect 23970 7584 23986 7648
rect 24050 7584 24066 7648
rect 24130 7584 24146 7648
rect 24210 7584 24218 7648
rect 21587 7444 21653 7445
rect 21587 7380 21588 7444
rect 21652 7380 21653 7444
rect 21587 7379 21653 7380
rect 20540 7040 20548 7104
rect 20612 7040 20628 7104
rect 20692 7040 20708 7104
rect 20772 7040 20788 7104
rect 20852 7040 20860 7104
rect 20540 6016 20860 7040
rect 20540 5952 20548 6016
rect 20612 5952 20628 6016
rect 20692 5952 20708 6016
rect 20772 5952 20788 6016
rect 20852 5952 20860 6016
rect 20540 4928 20860 5952
rect 20540 4864 20548 4928
rect 20612 4864 20628 4928
rect 20692 4864 20708 4928
rect 20772 4864 20788 4928
rect 20852 4864 20860 4928
rect 20540 3840 20860 4864
rect 20540 3776 20548 3840
rect 20612 3776 20628 3840
rect 20692 3776 20708 3840
rect 20772 3776 20788 3840
rect 20852 3776 20860 3840
rect 20540 2752 20860 3776
rect 20540 2688 20548 2752
rect 20612 2688 20628 2752
rect 20692 2688 20708 2752
rect 20772 2688 20788 2752
rect 20852 2688 20860 2752
rect 20299 2412 20365 2413
rect 20299 2348 20300 2412
rect 20364 2348 20365 2412
rect 20299 2347 20365 2348
rect 20302 2005 20362 2347
rect 20299 2004 20365 2005
rect 20299 1940 20300 2004
rect 20364 1940 20365 2004
rect 20299 1939 20365 1940
rect 20540 1664 20860 2688
rect 20540 1600 20548 1664
rect 20612 1600 20628 1664
rect 20692 1600 20708 1664
rect 20772 1600 20788 1664
rect 20852 1600 20860 1664
rect 19379 1460 19445 1461
rect 19379 1396 19380 1460
rect 19444 1396 19445 1460
rect 19379 1395 19445 1396
rect 17182 1056 17190 1120
rect 17254 1056 17270 1120
rect 17334 1056 17350 1120
rect 17414 1056 17430 1120
rect 17494 1056 17502 1120
rect 16251 916 16317 917
rect 16251 852 16252 916
rect 16316 852 16317 916
rect 16251 851 16317 852
rect 13824 512 13832 576
rect 13896 512 13912 576
rect 13976 512 13992 576
rect 14056 512 14072 576
rect 14136 512 14144 576
rect 13824 496 14144 512
rect 17182 496 17502 1056
rect 20540 576 20860 1600
rect 20540 512 20548 576
rect 20612 512 20628 576
rect 20692 512 20708 576
rect 20772 512 20788 576
rect 20852 512 20860 576
rect 20540 496 20860 512
rect 23898 6560 24218 7584
rect 23898 6496 23906 6560
rect 23970 6496 23986 6560
rect 24050 6496 24066 6560
rect 24130 6496 24146 6560
rect 24210 6496 24218 6560
rect 23898 5472 24218 6496
rect 23898 5408 23906 5472
rect 23970 5408 23986 5472
rect 24050 5408 24066 5472
rect 24130 5408 24146 5472
rect 24210 5408 24218 5472
rect 23898 4384 24218 5408
rect 23898 4320 23906 4384
rect 23970 4320 23986 4384
rect 24050 4320 24066 4384
rect 24130 4320 24146 4384
rect 24210 4320 24218 4384
rect 23898 3296 24218 4320
rect 23898 3232 23906 3296
rect 23970 3232 23986 3296
rect 24050 3232 24066 3296
rect 24130 3232 24146 3296
rect 24210 3232 24218 3296
rect 23898 2208 24218 3232
rect 23898 2144 23906 2208
rect 23970 2144 23986 2208
rect 24050 2144 24066 2208
rect 24130 2144 24146 2208
rect 24210 2144 24218 2208
rect 23898 1120 24218 2144
rect 23898 1056 23906 1120
rect 23970 1056 23986 1120
rect 24050 1056 24066 1120
rect 24130 1056 24146 1120
rect 24210 1056 24218 1120
rect 23898 496 24218 1056
rect 27256 9280 27576 10304
rect 27256 9216 27264 9280
rect 27328 9216 27344 9280
rect 27408 9216 27424 9280
rect 27488 9216 27504 9280
rect 27568 9216 27576 9280
rect 27256 8192 27576 9216
rect 27256 8128 27264 8192
rect 27328 8128 27344 8192
rect 27408 8128 27424 8192
rect 27488 8128 27504 8192
rect 27568 8128 27576 8192
rect 27256 7104 27576 8128
rect 27256 7040 27264 7104
rect 27328 7040 27344 7104
rect 27408 7040 27424 7104
rect 27488 7040 27504 7104
rect 27568 7040 27576 7104
rect 27256 6016 27576 7040
rect 27256 5952 27264 6016
rect 27328 5952 27344 6016
rect 27408 5952 27424 6016
rect 27488 5952 27504 6016
rect 27568 5952 27576 6016
rect 27256 4928 27576 5952
rect 27256 4864 27264 4928
rect 27328 4864 27344 4928
rect 27408 4864 27424 4928
rect 27488 4864 27504 4928
rect 27568 4864 27576 4928
rect 27256 3840 27576 4864
rect 27256 3776 27264 3840
rect 27328 3776 27344 3840
rect 27408 3776 27424 3840
rect 27488 3776 27504 3840
rect 27568 3776 27576 3840
rect 27256 2752 27576 3776
rect 27256 2688 27264 2752
rect 27328 2688 27344 2752
rect 27408 2688 27424 2752
rect 27488 2688 27504 2752
rect 27568 2688 27576 2752
rect 27256 1664 27576 2688
rect 27256 1600 27264 1664
rect 27328 1600 27344 1664
rect 27408 1600 27424 1664
rect 27488 1600 27504 1664
rect 27568 1600 27576 1664
rect 27256 576 27576 1600
rect 27256 512 27264 576
rect 27328 512 27344 576
rect 27408 512 27424 576
rect 27488 512 27504 576
rect 27568 512 27576 576
rect 27256 496 27576 512
use sky130_fd_sc_hd__buf_2  _381_
timestamp -7200
transform 1 0 15088 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp -7200
transform -1 0 14076 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _383_
timestamp -7200
transform 1 0 14076 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _384_
timestamp -7200
transform -1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _385_
timestamp -7200
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _386_
timestamp -7200
transform 1 0 20608 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp -7200
transform 1 0 10580 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp -7200
transform -1 0 11408 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _389_
timestamp -7200
transform 1 0 14444 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _390_
timestamp -7200
transform -1 0 11500 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _391_
timestamp -7200
transform 1 0 11592 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _392_
timestamp -7200
transform 1 0 3956 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _393_
timestamp -7200
transform 1 0 3956 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _394_
timestamp -7200
transform -1 0 6072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _395_
timestamp -7200
transform -1 0 7728 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _396_
timestamp -7200
transform -1 0 8004 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _397_
timestamp -7200
transform -1 0 6900 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _398_
timestamp -7200
transform 1 0 5152 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _399_
timestamp -7200
transform -1 0 6808 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _400_
timestamp -7200
transform 1 0 7268 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _401_
timestamp -7200
transform -1 0 11408 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _402_
timestamp -7200
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _403_
timestamp -7200
transform 1 0 7360 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _404_
timestamp -7200
transform 1 0 10856 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _405_
timestamp -7200
transform 1 0 8648 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _406_
timestamp -7200
transform -1 0 10028 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _407_
timestamp -7200
transform 1 0 9844 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _408_
timestamp -7200
transform 1 0 10120 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _409_
timestamp -7200
transform -1 0 10856 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _410_
timestamp -7200
transform -1 0 11132 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _411_
timestamp -7200
transform 1 0 6348 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp -7200
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _413_
timestamp -7200
transform -1 0 13616 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _414_
timestamp -7200
transform -1 0 16744 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _415_
timestamp -7200
transform -1 0 16008 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_4  _416_
timestamp -7200
transform 1 0 14168 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp -7200
transform -1 0 14352 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _418_
timestamp -7200
transform -1 0 17020 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _419_
timestamp -7200
transform 1 0 5796 0 -1 1632
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_2  _420_
timestamp -7200
transform -1 0 19228 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _421_
timestamp -7200
transform 1 0 4416 0 -1 1632
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_2  _422_
timestamp -7200
transform -1 0 19780 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _423_
timestamp -7200
transform -1 0 6532 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _424_
timestamp -7200
transform 1 0 21804 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _425_
timestamp -7200
transform 1 0 7452 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _426_
timestamp -7200
transform -1 0 20332 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _427_
timestamp -7200
transform 1 0 9016 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _428_
timestamp -7200
transform -1 0 21804 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _429_
timestamp -7200
transform -1 0 11868 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _430_
timestamp -7200
transform -1 0 20884 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _431_
timestamp -7200
transform 1 0 12512 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _432_
timestamp -7200
transform 1 0 14352 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  _433_
timestamp -7200
transform 1 0 13708 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _434_
timestamp -7200
transform 1 0 15456 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _435_
timestamp -7200
transform 1 0 16100 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _436_
timestamp -7200
transform -1 0 18952 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _437_
timestamp -7200
transform 1 0 18952 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _438_
timestamp -7200
transform -1 0 22540 0 -1 1632
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _439_
timestamp -7200
transform -1 0 21068 0 1 1632
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _440_
timestamp -7200
transform -1 0 20976 0 -1 1632
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _441_
timestamp -7200
transform -1 0 20976 0 1 544
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _442_
timestamp -7200
transform 1 0 14628 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _443_
timestamp -7200
transform -1 0 15180 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _444_
timestamp -7200
transform 1 0 15640 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _445_
timestamp -7200
transform -1 0 16008 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _446_
timestamp -7200
transform 1 0 15180 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _447_
timestamp -7200
transform -1 0 14720 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _448_
timestamp -7200
transform 1 0 14720 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _449_
timestamp -7200
transform -1 0 14904 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _450_
timestamp -7200
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _451_
timestamp -7200
transform 1 0 14352 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _452_
timestamp -7200
transform 1 0 14168 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _453_
timestamp -7200
transform -1 0 14444 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _454_
timestamp -7200
transform 1 0 13892 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _455_
timestamp -7200
transform 1 0 13340 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _456_
timestamp -7200
transform -1 0 13064 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _457_
timestamp -7200
transform 1 0 13524 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _458_
timestamp -7200
transform -1 0 13892 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _459_
timestamp -7200
transform 1 0 12512 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _460_
timestamp -7200
transform -1 0 12328 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _461_
timestamp -7200
transform 1 0 12604 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp -7200
transform 1 0 11684 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _463_
timestamp -7200
transform 1 0 11868 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _464_
timestamp -7200
transform 1 0 13524 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _465_
timestamp -7200
transform 1 0 11776 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _466_
timestamp -7200
transform -1 0 11776 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _467_
timestamp -7200
transform -1 0 14812 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _468_
timestamp -7200
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp -7200
transform 1 0 23368 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _470_
timestamp -7200
transform -1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _471_
timestamp -7200
transform 1 0 3864 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _472_
timestamp -7200
transform -1 0 4968 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _473_
timestamp -7200
transform -1 0 4876 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _474_
timestamp -7200
transform 1 0 3956 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _475_
timestamp -7200
transform 1 0 1748 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _476_
timestamp -7200
transform 1 0 2852 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _477_
timestamp -7200
transform -1 0 26220 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _478_
timestamp -7200
transform 1 0 1932 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _479_
timestamp -7200
transform 1 0 1564 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _480_
timestamp -7200
transform -1 0 4692 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _481_
timestamp -7200
transform 1 0 3404 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _482_
timestamp -7200
transform -1 0 3864 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _483_
timestamp -7200
transform -1 0 2668 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _484_
timestamp -7200
transform -1 0 3128 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _485_
timestamp -7200
transform -1 0 2668 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _486_
timestamp -7200
transform 1 0 2024 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _487_
timestamp -7200
transform 1 0 3864 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _488_
timestamp -7200
transform -1 0 4232 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _489_
timestamp -7200
transform 1 0 4232 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _490_
timestamp -7200
transform -1 0 5704 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _491_
timestamp -7200
transform -1 0 5336 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _492_
timestamp -7200
transform 1 0 5336 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _493_
timestamp -7200
transform -1 0 18124 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _494_
timestamp -7200
transform -1 0 17664 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _495_
timestamp -7200
transform -1 0 17112 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _496_
timestamp -7200
transform -1 0 23184 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _497_
timestamp -7200
transform 1 0 20516 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _498_
timestamp -7200
transform 1 0 20608 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _499_
timestamp -7200
transform -1 0 21712 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _500_
timestamp -7200
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _501_
timestamp -7200
transform 1 0 21712 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _502_
timestamp -7200
transform -1 0 20608 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_1  _503_
timestamp -7200
transform 1 0 18768 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _504_
timestamp -7200
transform 1 0 19044 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _505_
timestamp -7200
transform 1 0 18400 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _506_
timestamp -7200
transform 1 0 17756 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _507_
timestamp -7200
transform 1 0 18676 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _508_
timestamp -7200
transform -1 0 23276 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _509_
timestamp -7200
transform -1 0 23184 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _510_
timestamp -7200
transform -1 0 22632 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _511_
timestamp -7200
transform 1 0 22356 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _512_
timestamp -7200
transform 1 0 23828 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _513_
timestamp -7200
transform 1 0 23276 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _514_
timestamp -7200
transform 1 0 22816 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _515_
timestamp -7200
transform -1 0 24564 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _516_
timestamp -7200
transform -1 0 25760 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _517_
timestamp -7200
transform 1 0 24564 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _518_
timestamp -7200
transform 1 0 24104 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _519_
timestamp -7200
transform -1 0 24564 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _520_
timestamp -7200
transform -1 0 26128 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _521_
timestamp -7200
transform -1 0 25852 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _522_
timestamp -7200
transform 1 0 24196 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _523_
timestamp -7200
transform 1 0 24932 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _524_
timestamp -7200
transform -1 0 24196 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _525_
timestamp -7200
transform 1 0 25300 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _526_
timestamp -7200
transform 1 0 23920 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _527_
timestamp -7200
transform 1 0 25484 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _528_
timestamp -7200
transform 1 0 22172 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _529_
timestamp -7200
transform -1 0 23552 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _530_
timestamp -7200
transform -1 0 22448 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _531_
timestamp -7200
transform -1 0 21712 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _532_
timestamp -7200
transform -1 0 23736 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _533_
timestamp -7200
transform 1 0 22816 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _534_
timestamp -7200
transform 1 0 22356 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _535_
timestamp -7200
transform -1 0 24012 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _536_
timestamp -7200
transform 1 0 22448 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _537_
timestamp -7200
transform 1 0 21252 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _538_
timestamp -7200
transform -1 0 22264 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _539_
timestamp -7200
transform 1 0 21344 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _540_
timestamp -7200
transform 1 0 20700 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _541_
timestamp -7200
transform 1 0 19504 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _542_
timestamp -7200
transform 1 0 19596 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _543_
timestamp -7200
transform -1 0 17664 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _544_
timestamp -7200
transform 1 0 17112 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _545_
timestamp -7200
transform -1 0 17388 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _546_
timestamp -7200
transform 1 0 16652 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _547_
timestamp -7200
transform -1 0 16008 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _548_
timestamp -7200
transform 1 0 10212 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _549_
timestamp -7200
transform -1 0 12144 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _550_
timestamp -7200
transform 1 0 7820 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _551_
timestamp -7200
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _552_
timestamp -7200
transform 1 0 11500 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _553_
timestamp -7200
transform 1 0 9200 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _554_
timestamp -7200
transform 1 0 8464 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _555_
timestamp -7200
transform -1 0 13432 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _556_
timestamp -7200
transform -1 0 10856 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _557_
timestamp -7200
transform 1 0 7912 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _558_
timestamp -7200
transform 1 0 13340 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _559_
timestamp -7200
transform 1 0 15548 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _560_
timestamp -7200
transform -1 0 10856 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _561_
timestamp -7200
transform -1 0 10120 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _562_
timestamp -7200
transform 1 0 10856 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _563_
timestamp -7200
transform 1 0 6164 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _564_
timestamp -7200
transform -1 0 10396 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _565_
timestamp -7200
transform -1 0 8280 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _566_
timestamp -7200
transform 1 0 9844 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _567_
timestamp -7200
transform 1 0 9292 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _568_
timestamp -7200
transform -1 0 8004 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _569_
timestamp -7200
transform -1 0 6164 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _570_
timestamp -7200
transform -1 0 4968 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _571_
timestamp -7200
transform -1 0 5244 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _572_
timestamp -7200
transform 1 0 3220 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _573_
timestamp -7200
transform 1 0 2576 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _574_
timestamp -7200
transform -1 0 6164 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _575_
timestamp -7200
transform -1 0 2024 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _576_
timestamp -7200
transform 1 0 1840 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _577_
timestamp -7200
transform 1 0 2852 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _578_
timestamp -7200
transform -1 0 4048 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _579_
timestamp -7200
transform 1 0 2024 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _580_
timestamp -7200
transform -1 0 4784 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _581_
timestamp -7200
transform -1 0 4324 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _582_
timestamp -7200
transform 1 0 3220 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _583_
timestamp -7200
transform 1 0 3312 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _584_
timestamp -7200
transform 1 0 2300 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _585_
timestamp -7200
transform 1 0 12144 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _586_
timestamp -7200
transform -1 0 5612 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _587_
timestamp -7200
transform 1 0 4968 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _588_
timestamp -7200
transform 1 0 4784 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _589_
timestamp -7200
transform 1 0 5244 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _590_
timestamp -7200
transform 1 0 8740 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _591_
timestamp -7200
transform -1 0 10028 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _592_
timestamp -7200
transform 1 0 11040 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _593_
timestamp -7200
transform 1 0 8280 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _594_
timestamp -7200
transform 1 0 9200 0 -1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _595_
timestamp -7200
transform 1 0 10948 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _596_
timestamp -7200
transform -1 0 12144 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _597_
timestamp -7200
transform 1 0 8372 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _598_
timestamp -7200
transform -1 0 10212 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _599_
timestamp -7200
transform -1 0 9016 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _600_
timestamp -7200
transform 1 0 4600 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _601_
timestamp -7200
transform 1 0 8924 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _602_
timestamp -7200
transform 1 0 10212 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _603_
timestamp -7200
transform -1 0 9660 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _604_
timestamp -7200
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _605_
timestamp -7200
transform -1 0 9568 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _606_
timestamp -7200
transform 1 0 7544 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _607_
timestamp -7200
transform -1 0 9200 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _608_
timestamp -7200
transform 1 0 8648 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _609_
timestamp -7200
transform -1 0 9660 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _610_
timestamp -7200
transform 1 0 9384 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _611_
timestamp -7200
transform -1 0 12788 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _612_
timestamp -7200
transform 1 0 9292 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _613_
timestamp -7200
transform -1 0 10856 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _614_
timestamp -7200
transform 1 0 11132 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _615_
timestamp -7200
transform -1 0 13340 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _616_
timestamp -7200
transform -1 0 14076 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _617_
timestamp -7200
transform 1 0 11868 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _618_
timestamp -7200
transform 1 0 12144 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _619_
timestamp -7200
transform 1 0 12420 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _620_
timestamp -7200
transform 1 0 20516 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _621_
timestamp -7200
transform 1 0 18676 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _622_
timestamp -7200
transform 1 0 23276 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _623_
timestamp -7200
transform 1 0 19412 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _624_
timestamp -7200
transform 1 0 18216 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _625_
timestamp -7200
transform 1 0 19412 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _626_
timestamp -7200
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _627_
timestamp -7200
transform 1 0 16836 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _628_
timestamp -7200
transform 1 0 18400 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _629_
timestamp -7200
transform 1 0 20884 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _630_
timestamp -7200
transform -1 0 22816 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _631_
timestamp -7200
transform 1 0 23828 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _632_
timestamp -7200
transform -1 0 25300 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _633_
timestamp -7200
transform 1 0 25576 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _634_
timestamp -7200
transform 1 0 25484 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _635_
timestamp -7200
transform 1 0 26312 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _636_
timestamp -7200
transform -1 0 26404 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _637_
timestamp -7200
transform 1 0 26404 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _638_
timestamp -7200
transform 1 0 26404 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _639_
timestamp -7200
transform -1 0 24748 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _640_
timestamp -7200
transform -1 0 24840 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _641_
timestamp -7200
transform -1 0 23276 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _642_
timestamp -7200
transform 1 0 22172 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _643_
timestamp -7200
transform -1 0 22816 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _644_
timestamp -7200
transform 1 0 19228 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _645_
timestamp -7200
transform -1 0 20884 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _646_
timestamp -7200
transform 1 0 20332 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _647_
timestamp -7200
transform -1 0 19412 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _648_
timestamp -7200
transform 1 0 17572 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _649_
timestamp -7200
transform 1 0 18676 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _650_
timestamp -7200
transform -1 0 17112 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _651_
timestamp -7200
transform -1 0 15272 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _652_
timestamp -7200
transform -1 0 16192 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _653_
timestamp -7200
transform 1 0 13800 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _654_
timestamp -7200
transform 1 0 23552 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _655_
timestamp -7200
transform 1 0 16100 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _656_
timestamp -7200
transform 1 0 14536 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _657_
timestamp -7200
transform 1 0 5244 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _658_
timestamp -7200
transform -1 0 7268 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _659_
timestamp -7200
transform 1 0 7268 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _660_
timestamp -7200
transform 1 0 4784 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _661_
timestamp -7200
transform -1 0 8464 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _662_
timestamp -7200
transform 1 0 5704 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _663_
timestamp -7200
transform 1 0 5244 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _664_
timestamp -7200
transform -1 0 7268 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _665_
timestamp -7200
transform 1 0 5980 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _666_
timestamp -7200
transform 1 0 5520 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _667_
timestamp -7200
transform -1 0 8648 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _668_
timestamp -7200
transform 1 0 6900 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _669_
timestamp -7200
transform 1 0 5520 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _670_
timestamp -7200
transform -1 0 8188 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _671_
timestamp -7200
transform -1 0 6900 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _672_
timestamp -7200
transform 1 0 5980 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _673_
timestamp -7200
transform 1 0 8372 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _674_
timestamp -7200
transform 1 0 8372 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _675_
timestamp -7200
transform 1 0 8924 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _676_
timestamp -7200
transform 1 0 12144 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _677_
timestamp -7200
transform 1 0 10948 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _678_
timestamp -7200
transform 1 0 15916 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _679_
timestamp -7200
transform 1 0 15824 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _680_
timestamp -7200
transform 1 0 15364 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _681_
timestamp -7200
transform -1 0 15732 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _682_
timestamp -7200
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _683_
timestamp -7200
transform 1 0 20148 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _684_
timestamp -7200
transform 1 0 19688 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _685_
timestamp -7200
transform 1 0 18952 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _686_
timestamp -7200
transform -1 0 19228 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _687_
timestamp -7200
transform -1 0 19320 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _688_
timestamp -7200
transform 1 0 21988 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _689_
timestamp -7200
transform 1 0 21252 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _690_
timestamp -7200
transform 1 0 24564 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _691_
timestamp -7200
transform 1 0 22080 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _692_
timestamp -7200
transform -1 0 23644 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _693_
timestamp -7200
transform -1 0 24748 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _694_
timestamp -7200
transform -1 0 25484 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _695_
timestamp -7200
transform 1 0 25484 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _696_
timestamp -7200
transform -1 0 25484 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _697_
timestamp -7200
transform 1 0 24840 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _698_
timestamp -7200
transform -1 0 24748 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _699_
timestamp -7200
transform 1 0 22908 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _700_
timestamp -7200
transform -1 0 23552 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _701_
timestamp -7200
transform -1 0 22540 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _702_
timestamp -7200
transform 1 0 22724 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _703_
timestamp -7200
transform -1 0 21988 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _704_
timestamp -7200
transform -1 0 22356 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _705_
timestamp -7200
transform -1 0 18584 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _706_
timestamp -7200
transform 1 0 20148 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _707_
timestamp -7200
transform -1 0 18308 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _708_
timestamp -7200
transform 1 0 17664 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _709_
timestamp -7200
transform -1 0 17480 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _710_
timestamp -7200
transform 1 0 16928 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _711_
timestamp -7200
transform 1 0 16008 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _712_
timestamp -7200
transform -1 0 13432 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _713_
timestamp -7200
transform 1 0 13432 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _714_
timestamp -7200
transform -1 0 15456 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _715_
timestamp -7200
transform 1 0 15088 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _716_
timestamp -7200
transform 1 0 15824 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _717_
timestamp -7200
transform -1 0 15088 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _718_
timestamp -7200
transform -1 0 10304 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _719_
timestamp -7200
transform -1 0 14444 0 -1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_2  _720_
timestamp -7200
transform 1 0 7820 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _721_
timestamp -7200
transform -1 0 9844 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _722_
timestamp -7200
transform 1 0 10028 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _723_
timestamp -7200
transform 1 0 9016 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _724_
timestamp -7200
transform 1 0 4876 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _725_
timestamp -7200
transform 1 0 7268 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _726_
timestamp -7200
transform 1 0 3404 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _727_
timestamp -7200
transform 1 0 8372 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _728_
timestamp -7200
transform 1 0 6532 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _729_
timestamp -7200
transform 1 0 7912 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _730_
timestamp -7200
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _731_
timestamp -7200
transform -1 0 9200 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _732_
timestamp -7200
transform 1 0 8556 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _733_
timestamp -7200
transform -1 0 10856 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _734_
timestamp -7200
transform -1 0 11684 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _735_
timestamp -7200
transform -1 0 10948 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _736_
timestamp -7200
transform -1 0 11684 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _737_
timestamp -7200
transform -1 0 9200 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _738_
timestamp -7200
transform -1 0 8740 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _739_
timestamp -7200
transform -1 0 10396 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _740_
timestamp -7200
transform -1 0 9936 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _741_
timestamp -7200
transform -1 0 9476 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _742_
timestamp -7200
transform -1 0 5704 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _743_
timestamp -7200
transform 1 0 5244 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _744_
timestamp -7200
transform 1 0 6256 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _745_
timestamp -7200
transform 1 0 5704 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _746_
timestamp -7200
transform -1 0 6256 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _747_
timestamp -7200
transform 1 0 4324 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _748_
timestamp -7200
transform -1 0 7176 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _749_
timestamp -7200
transform -1 0 4048 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _750_
timestamp -7200
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _751_
timestamp -7200
transform -1 0 7912 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _752_
timestamp -7200
transform 1 0 7360 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _753_
timestamp -7200
transform 1 0 7452 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _754_
timestamp -7200
transform -1 0 9752 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _755_
timestamp -7200
transform 1 0 8648 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _756_
timestamp -7200
transform -1 0 9200 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _757_
timestamp -7200
transform -1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _758_
timestamp -7200
transform 1 0 12052 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _759_
timestamp -7200
transform 1 0 12236 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _760_
timestamp -7200
transform -1 0 12972 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _761_
timestamp -7200
transform 1 0 12144 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _762_
timestamp -7200
transform 1 0 12512 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _763_
timestamp -7200
transform 1 0 12696 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _764_
timestamp -7200
transform -1 0 14628 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _765_
timestamp -7200
transform 1 0 13708 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _766_
timestamp -7200
transform 1 0 15640 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _767_
timestamp -7200
transform 1 0 16008 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _768_
timestamp -7200
transform 1 0 16652 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _769_
timestamp -7200
transform -1 0 17020 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _770_
timestamp -7200
transform 1 0 16100 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _771_
timestamp -7200
transform -1 0 17572 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _772_
timestamp -7200
transform 1 0 17020 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _773_
timestamp -7200
transform 1 0 16100 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _774_
timestamp -7200
transform 1 0 16744 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _775_
timestamp -7200
transform -1 0 17388 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _776_
timestamp -7200
transform 1 0 15916 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _777_
timestamp -7200
transform -1 0 19136 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _778_
timestamp -7200
transform -1 0 18768 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _779_
timestamp -7200
transform 1 0 15272 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _780_
timestamp -7200
transform 1 0 17940 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _781_
timestamp -7200
transform -1 0 19044 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _782_
timestamp -7200
transform 1 0 14628 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _783_
timestamp -7200
transform 1 0 17756 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _784_
timestamp -7200
transform -1 0 18584 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _785_
timestamp -7200
transform 1 0 15456 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _786_
timestamp -7200
transform 1 0 17204 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _787_
timestamp -7200
transform -1 0 18308 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _788_
timestamp -7200
transform 1 0 1564 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _789_
timestamp -7200
transform 1 0 2392 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _790_
timestamp -7200
transform 1 0 1380 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _791_
timestamp -7200
transform 1 0 2668 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _792_
timestamp -7200
transform 1 0 1472 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _793_
timestamp -7200
transform 1 0 3404 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _794_
timestamp -7200
transform 1 0 4876 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _795_
timestamp -7200
transform 1 0 17112 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _796_
timestamp -7200
transform -1 0 21344 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _797_
timestamp -7200
transform 1 0 19412 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _798_
timestamp -7200
transform 1 0 17112 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _799_
timestamp -7200
transform 1 0 22632 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _800_
timestamp -7200
transform 1 0 22540 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _801_
timestamp -7200
transform -1 0 26036 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _802_
timestamp -7200
transform 1 0 25116 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _803_
timestamp -7200
transform -1 0 26128 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _804_
timestamp -7200
transform 1 0 25116 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _805_
timestamp -7200
transform 1 0 21804 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _806_
timestamp -7200
transform -1 0 25484 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _807_
timestamp -7200
transform -1 0 22816 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _808_
timestamp -7200
transform 1 0 19228 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _809_
timestamp -7200
transform 1 0 16468 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _810_
timestamp -7200
transform 1 0 15824 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _811_
timestamp -7200
transform 1 0 11960 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _812_
timestamp -7200
transform 1 0 5796 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _813_
timestamp -7200
transform 1 0 10580 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _814_
timestamp -7200
transform 1 0 6900 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _815_
timestamp -7200
transform 1 0 5060 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _816_
timestamp -7200
transform 1 0 12512 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _817_
timestamp -7200
transform 1 0 8188 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _818_
timestamp -7200
transform 1 0 6440 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _819_
timestamp -7200
transform -1 0 12420 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _820_
timestamp -7200
transform 1 0 2392 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _821_
timestamp -7200
transform 1 0 1472 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _822_
timestamp -7200
transform 1 0 1380 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _823_
timestamp -7200
transform 1 0 1656 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _824_
timestamp -7200
transform 1 0 4876 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _825_
timestamp -7200
transform 1 0 11408 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _826_
timestamp -7200
transform 1 0 9200 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _827_
timestamp -7200
transform 1 0 9568 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _828_
timestamp -7200
transform 1 0 9016 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _829_
timestamp -7200
transform 1 0 9660 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _830_
timestamp -7200
transform 1 0 13524 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _831_
timestamp -7200
transform 1 0 11040 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _832_
timestamp -7200
transform 1 0 12788 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _833_
timestamp -7200
transform 1 0 11592 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _834_
timestamp -7200
transform 1 0 12328 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _835_
timestamp -7200
transform 1 0 18584 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _836_
timestamp -7200
transform 1 0 19688 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _837_
timestamp -7200
transform 1 0 21620 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _838_
timestamp -7200
transform 1 0 23460 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _839_
timestamp -7200
transform 1 0 25300 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _840_
timestamp -7200
transform 1 0 24840 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _841_
timestamp -7200
transform 1 0 24840 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _842_
timestamp -7200
transform -1 0 25300 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _843_
timestamp -7200
transform 1 0 21068 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _844_
timestamp -7200
transform 1 0 18676 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _845_
timestamp -7200
transform 1 0 17204 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _846_
timestamp -7200
transform 1 0 15640 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _847_
timestamp -7200
transform 1 0 13984 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _848_
timestamp -7200
transform 1 0 14076 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _849_
timestamp -7200
transform 1 0 14076 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _850_
timestamp -7200
transform 1 0 5796 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _851_
timestamp -7200
transform 1 0 4324 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _852_
timestamp -7200
transform 1 0 5796 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _853_
timestamp -7200
transform 1 0 6716 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _854_
timestamp -7200
transform 1 0 6532 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _855_
timestamp -7200
transform 1 0 7452 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _856_
timestamp -7200
transform 1 0 9568 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _857_
timestamp -7200
transform -1 0 16376 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _858_
timestamp -7200
transform -1 0 15824 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _859_
timestamp -7200
transform 1 0 18860 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _860_
timestamp -7200
transform 1 0 18676 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _861_
timestamp -7200
transform 1 0 21068 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _862_
timestamp -7200
transform 1 0 22724 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _863_
timestamp -7200
transform 1 0 24840 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _864_
timestamp -7200
transform 1 0 24840 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _865_
timestamp -7200
transform 1 0 25208 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _866_
timestamp -7200
transform 1 0 23828 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _867_
timestamp -7200
transform 1 0 21160 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _868_
timestamp -7200
transform -1 0 22724 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _869_
timestamp -7200
transform 1 0 18308 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _870_
timestamp -7200
transform 1 0 17112 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _871_
timestamp -7200
transform -1 0 18032 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _872_
timestamp -7200
transform 1 0 13340 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _873_
timestamp -7200
transform -1 0 15824 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _874_
timestamp -7200
transform 1 0 8740 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _875_
timestamp -7200
transform 1 0 4048 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _876_
timestamp -7200
transform 1 0 3772 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _877_
timestamp -7200
transform 1 0 4232 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _878_
timestamp -7200
transform 1 0 6440 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _879_
timestamp -7200
transform 1 0 8280 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _880_
timestamp -7200
transform 1 0 11040 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _881_
timestamp -7200
transform 1 0 10948 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _882_
timestamp -7200
transform 1 0 8372 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _883_
timestamp -7200
transform 1 0 9936 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _884_
timestamp -7200
transform -1 0 6440 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _885_
timestamp -7200
transform 1 0 3772 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _886_
timestamp -7200
transform 1 0 3312 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _887_
timestamp -7200
transform 1 0 7268 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _888_
timestamp -7200
transform 1 0 9292 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _889_
timestamp -7200
transform -1 0 13524 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _890_
timestamp -7200
transform 1 0 11868 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _891_
timestamp -7200
transform -1 0 15548 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _892_
timestamp -7200
transform -1 0 17480 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _893_
timestamp -7200
transform 1 0 16744 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _894_
timestamp -7200
transform 1 0 17388 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _895_
timestamp -7200
transform 1 0 19412 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _896_
timestamp -7200
transform 1 0 19044 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _897_
timestamp -7200
transform 1 0 18676 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _898_
timestamp -7200
transform 1 0 18860 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _909_
timestamp -7200
transform -1 0 10856 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _910_
timestamp -7200
transform -1 0 10028 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _911_
timestamp -7200
transform 1 0 7912 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _912_
timestamp -7200
transform 1 0 6900 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -7200
transform -1 0 15824 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp -7200
transform 1 0 6348 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp -7200
transform -1 0 11500 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp -7200
transform -1 0 8096 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp -7200
transform 1 0 9568 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp -7200
transform -1 0 20516 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp -7200
transform 1 0 21712 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp -7200
transform -1 0 20516 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp -7200
transform 1 0 21620 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  digital_top_14
timestamp -7200
transform -1 0 4324 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_15
timestamp -7200
transform -1 0 1748 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_16
timestamp -7200
transform -1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_17
timestamp -7200
transform -1 0 9476 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_18
timestamp -7200
transform -1 0 6900 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_19
timestamp -7200
transform -1 0 6256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_20
timestamp -7200
transform 1 0 5336 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_21
timestamp -7200
transform 1 0 4692 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_22
timestamp -7200
transform 1 0 3404 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  digital_top_23
timestamp -7200
transform 1 0 2760 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp -7200
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp -7200
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp -7200
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp -7200
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp -7200
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp -7200
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_65
timestamp -7200
transform 1 0 6532 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_73
timestamp -7200
transform 1 0 7268 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp -7200
transform 1 0 8188 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_85
timestamp -7200
transform 1 0 8372 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_91
timestamp -7200
transform 1 0 8924 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_100
timestamp -7200
transform 1 0 9752 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp -7200
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_125
timestamp -7200
transform 1 0 12052 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_129
timestamp -7200
transform 1 0 12420 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138
timestamp -7200
transform 1 0 13248 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_141
timestamp -7200
transform 1 0 13524 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_163
timestamp -7200
transform 1 0 15548 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp -7200
transform 1 0 15916 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_177
timestamp -7200
transform 1 0 16836 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_189
timestamp -7200
transform 1 0 17940 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp -7200
transform 1 0 18492 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_197
timestamp -7200
transform 1 0 18676 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_205
timestamp -7200
transform 1 0 19412 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_222
timestamp -7200
transform 1 0 20976 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp -7200
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp -7200
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp -7200
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp -7200
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp -7200
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp -7200
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_281
timestamp -7200
transform 1 0 26404 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp -7200
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp -7200
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp -7200
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_39
timestamp -7200
transform 1 0 4140 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_71
timestamp -7200
transform 1 0 7084 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_89
timestamp -7200
transform 1 0 8740 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp -7200
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp -7200
transform 1 0 10948 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_123
timestamp -7200
transform 1 0 11868 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_141
timestamp -7200
transform 1 0 13524 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp -7200
transform 1 0 15824 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_169
timestamp -7200
transform 1 0 16100 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_175
timestamp -7200
transform 1 0 16652 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_222
timestamp -7200
transform 1 0 20976 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_239
timestamp -7200
transform 1 0 22540 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_251
timestamp -7200
transform 1 0 23644 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_263
timestamp -7200
transform 1 0 24748 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_275
timestamp -7200
transform 1 0 25852 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp -7200
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_281
timestamp -7200
transform 1 0 26404 0 -1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp -7200
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp -7200
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp -7200
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp -7200
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_44
timestamp -7200
transform 1 0 4600 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_64
timestamp -7200
transform 1 0 6440 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_72
timestamp -7200
transform 1 0 7176 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_78
timestamp -7200
transform 1 0 7728 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_85
timestamp -7200
transform 1 0 8372 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_118
timestamp -7200
transform 1 0 11408 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_126
timestamp -7200
transform 1 0 12144 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_135
timestamp -7200
transform 1 0 12972 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp -7200
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_141
timestamp -7200
transform 1 0 13524 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_167
timestamp -7200
transform 1 0 15916 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_184
timestamp -7200
transform 1 0 17480 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp -7200
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_223
timestamp -7200
transform 1 0 21068 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_235
timestamp -7200
transform 1 0 22172 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_247
timestamp -7200
transform 1 0 23276 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp -7200
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp -7200
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp -7200
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp -7200
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp -7200
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp -7200
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_27
timestamp -7200
transform 1 0 3036 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_65
timestamp -7200
transform 1 0 6532 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_73
timestamp -7200
transform 1 0 7268 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_79
timestamp -7200
transform 1 0 7820 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_87
timestamp -7200
transform 1 0 8556 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_107
timestamp -7200
transform 1 0 10396 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp -7200
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_113
timestamp -7200
transform 1 0 10948 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_121
timestamp -7200
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_139
timestamp -7200
transform 1 0 13340 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_145
timestamp -7200
transform 1 0 13892 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_162
timestamp -7200
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_169
timestamp -7200
transform 1 0 16100 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_182
timestamp -7200
transform 1 0 17296 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_194
timestamp -7200
transform 1 0 18400 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_206
timestamp -7200
transform 1 0 19504 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_218
timestamp -7200
transform 1 0 20608 0 -1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp -7200
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp -7200
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp -7200
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp -7200
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp -7200
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp -7200
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_281
timestamp -7200
transform 1 0 26404 0 -1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp -7200
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp -7200
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp -7200
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_29
timestamp -7200
transform 1 0 3220 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_46
timestamp -7200
transform 1 0 4784 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_63
timestamp -7200
transform 1 0 6348 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_71
timestamp -7200
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_80
timestamp -7200
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_85
timestamp -7200
transform 1 0 8372 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_105
timestamp -7200
transform 1 0 10212 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_117
timestamp -7200
transform 1 0 11316 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_135
timestamp -7200
transform 1 0 12972 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp -7200
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp -7200
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_153
timestamp -7200
transform 1 0 14628 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_185
timestamp -7200
transform 1 0 17572 0 1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_213
timestamp -7200
transform 1 0 20148 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_225
timestamp -7200
transform 1 0 21252 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_237
timestamp -7200
transform 1 0 22356 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_249
timestamp -7200
transform 1 0 23460 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp -7200
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp -7200
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp -7200
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp -7200
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp -7200
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_27
timestamp -7200
transform 1 0 3036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_31
timestamp -7200
transform 1 0 3404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp -7200
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp -7200
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_57
timestamp -7200
transform 1 0 5796 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_63
timestamp -7200
transform 1 0 6348 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_80
timestamp -7200
transform 1 0 7912 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_100
timestamp -7200
transform 1 0 9752 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp -7200
transform 1 0 10948 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_135
timestamp -7200
transform 1 0 12972 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_143
timestamp -7200
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_163
timestamp -7200
transform 1 0 15548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp -7200
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_176
timestamp -7200
transform 1 0 16744 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_184
timestamp -7200
transform 1 0 17480 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_192
timestamp -7200
transform 1 0 18216 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp -7200
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp -7200
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp -7200
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp -7200
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp -7200
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp -7200
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp -7200
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp -7200
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_281
timestamp -7200
transform 1 0 26404 0 -1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp -7200
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp -7200
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp -7200
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_29
timestamp -7200
transform 1 0 3220 0 1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_54
timestamp -7200
transform 1 0 5520 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_66
timestamp -7200
transform 1 0 6624 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp -7200
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_111
timestamp -7200
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_121
timestamp -7200
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_150
timestamp -7200
transform 1 0 14352 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_174
timestamp -7200
transform 1 0 16560 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_186
timestamp -7200
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp -7200
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_202
timestamp -7200
transform 1 0 19136 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp -7200
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_233
timestamp -7200
transform 1 0 21988 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_241
timestamp -7200
transform 1 0 22724 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp -7200
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp -7200
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp -7200
transform 1 0 23828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp -7200
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp -7200
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp -7200
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp -7200
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_27
timestamp -7200
transform 1 0 3036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp -7200
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_72
timestamp -7200
transform 1 0 7176 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_101
timestamp -7200
transform 1 0 9844 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_121
timestamp -7200
transform 1 0 11684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_125
timestamp -7200
transform 1 0 12052 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_133
timestamp -7200
transform 1 0 12788 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_145
timestamp -7200
transform 1 0 13892 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_157
timestamp -7200
transform 1 0 14996 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_162
timestamp -7200
transform 1 0 15456 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_169
timestamp -7200
transform 1 0 16100 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_177
timestamp -7200
transform 1 0 16836 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_215
timestamp -7200
transform 1 0 20332 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp -7200
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp -7200
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_237
timestamp -7200
transform 1 0 22356 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_255
timestamp -7200
transform 1 0 24012 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_267
timestamp -7200
transform 1 0 25116 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp -7200
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_281
timestamp -7200
transform 1 0 26404 0 -1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp -7200
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp -7200
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp -7200
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp -7200
transform 1 0 3220 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_37
timestamp -7200
transform 1 0 3956 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_56
timestamp -7200
transform 1 0 5704 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_73
timestamp -7200
transform 1 0 7268 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_119
timestamp -7200
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp -7200
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_159
timestamp -7200
transform 1 0 15180 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_186
timestamp -7200
transform 1 0 17664 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp -7200
transform 1 0 18308 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_197
timestamp -7200
transform 1 0 18676 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_205
timestamp -7200
transform 1 0 19412 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_209
timestamp -7200
transform 1 0 19780 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_226
timestamp -7200
transform 1 0 21344 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_234
timestamp -7200
transform 1 0 22080 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_262
timestamp -7200
transform 1 0 24656 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_266
timestamp -7200
transform 1 0 25024 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_275
timestamp -7200
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_287
timestamp -7200
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp -7200
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp -7200
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp -7200
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp -7200
transform 1 0 4140 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_47
timestamp -7200
transform 1 0 4876 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp -7200
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_65
timestamp -7200
transform 1 0 6532 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_77
timestamp -7200
transform 1 0 7636 0 -1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_94
timestamp -7200
transform 1 0 9200 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_106
timestamp -7200
transform 1 0 10304 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_158
timestamp -7200
transform 1 0 15088 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp -7200
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp -7200
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_181
timestamp -7200
transform 1 0 17204 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_199
timestamp -7200
transform 1 0 18860 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_230
timestamp -7200
transform 1 0 21712 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_236
timestamp -7200
transform 1 0 22264 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_256
timestamp -7200
transform 1 0 24104 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_277
timestamp -7200
transform 1 0 26036 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_281
timestamp -7200
transform 1 0 26404 0 -1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp -7200
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_15
timestamp -7200
transform 1 0 1932 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29
timestamp -7200
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp -7200
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_101
timestamp -7200
transform 1 0 9844 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_121
timestamp -7200
transform 1 0 11684 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_131
timestamp -7200
transform 1 0 12604 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp -7200
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_145
timestamp -7200
transform 1 0 13892 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_149
timestamp -7200
transform 1 0 14260 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_170
timestamp -7200
transform 1 0 16192 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_176
timestamp -7200
transform 1 0 16744 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_238
timestamp -7200
transform 1 0 22448 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_246
timestamp -7200
transform 1 0 23184 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_266
timestamp -7200
transform 1 0 25024 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_283
timestamp -7200
transform 1 0 26588 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_3
timestamp -7200
transform 1 0 828 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_9
timestamp -7200
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_34
timestamp -7200
transform 1 0 3680 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp -7200
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_69
timestamp -7200
transform 1 0 6900 0 -1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_96
timestamp -7200
transform 1 0 9384 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_108
timestamp -7200
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_113
timestamp -7200
transform 1 0 10948 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_117
timestamp -7200
transform 1 0 11316 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_131
timestamp -7200
transform 1 0 12604 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_139
timestamp -7200
transform 1 0 13340 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp -7200
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_181
timestamp -7200
transform 1 0 17204 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_201
timestamp -7200
transform 1 0 19044 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_221
timestamp -7200
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_225
timestamp -7200
transform 1 0 21252 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_247
timestamp -7200
transform 1 0 23276 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_253
timestamp -7200
transform 1 0 23828 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_278
timestamp -7200
transform 1 0 26128 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp -7200
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp -7200
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp -7200
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_47
timestamp -7200
transform 1 0 4876 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_53
timestamp -7200
transform 1 0 5428 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_64
timestamp -7200
transform 1 0 6440 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp -7200
transform 1 0 8004 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_93
timestamp -7200
transform 1 0 9108 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_97
timestamp -7200
transform 1 0 9476 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_130
timestamp -7200
transform 1 0 12512 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp -7200
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_157
timestamp -7200
transform 1 0 14996 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_173
timestamp -7200
transform 1 0 16468 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_179
timestamp -7200
transform 1 0 17020 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_200
timestamp -7200
transform 1 0 18952 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_208
timestamp -7200
transform 1 0 19688 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_220
timestamp -7200
transform 1 0 20792 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_226
timestamp -7200
transform 1 0 21344 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp -7200
transform 1 0 23552 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp -7200
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_275
timestamp -7200
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_287
timestamp -7200
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp -7200
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_15
timestamp -7200
transform 1 0 1932 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_19
timestamp -7200
transform 1 0 2300 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp -7200
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp -7200
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp -7200
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_57
timestamp -7200
transform 1 0 5796 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_77
timestamp -7200
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_87
timestamp -7200
transform 1 0 8556 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp -7200
transform 1 0 10948 0 -1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp -7200
transform 1 0 14260 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp -7200
transform 1 0 15364 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp -7200
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp -7200
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp -7200
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp -7200
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_205
timestamp -7200
transform 1 0 19412 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_213
timestamp -7200
transform 1 0 20148 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_217
timestamp -7200
transform 1 0 20516 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_225
timestamp -7200
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_233
timestamp -7200
transform 1 0 21988 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_250
timestamp -7200
transform 1 0 23552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_278
timestamp -7200
transform 1 0 26128 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp -7200
transform 1 0 828 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp -7200
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp -7200
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_45
timestamp -7200
transform 1 0 4692 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_53
timestamp -7200
transform 1 0 5428 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_59
timestamp -7200
transform 1 0 5980 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_67
timestamp -7200
transform 1 0 6716 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp -7200
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_90
timestamp -7200
transform 1 0 8832 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_94
timestamp -7200
transform 1 0 9200 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_103
timestamp -7200
transform 1 0 10028 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp -7200
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp -7200
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_153
timestamp -7200
transform 1 0 14628 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_184
timestamp -7200
transform 1 0 17480 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp -7200
transform 1 0 17940 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp -7200
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_197
timestamp -7200
transform 1 0 18676 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_226
timestamp -7200
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_236
timestamp -7200
transform 1 0 22264 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_244
timestamp -7200
transform 1 0 23000 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_253
timestamp -7200
transform 1 0 23828 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_266
timestamp -7200
transform 1 0 25024 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_283
timestamp -7200
transform 1 0 26588 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp -7200
transform 1 0 828 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_27
timestamp -7200
transform 1 0 3036 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp -7200
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp -7200
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp -7200
transform 1 0 5796 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_65
timestamp -7200
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_96
timestamp -7200
transform 1 0 9384 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_108
timestamp -7200
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_113
timestamp -7200
transform 1 0 10948 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_121
timestamp -7200
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_147
timestamp -7200
transform 1 0 14076 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_166
timestamp -7200
transform 1 0 15824 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_169
timestamp -7200
transform 1 0 16100 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_203
timestamp -7200
transform 1 0 19228 0 -1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_210
timestamp -7200
transform 1 0 19872 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp -7200
transform 1 0 20976 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_228
timestamp -7200
transform 1 0 21528 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp -7200
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_281
timestamp -7200
transform 1 0 26404 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_3
timestamp -7200
transform 1 0 828 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_48
timestamp -7200
transform 1 0 4968 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_64
timestamp -7200
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_85
timestamp -7200
transform 1 0 8372 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_115
timestamp -7200
transform 1 0 11132 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_119
timestamp -7200
transform 1 0 11500 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp -7200
transform 1 0 13064 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_141
timestamp -7200
transform 1 0 13524 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_145
timestamp -7200
transform 1 0 13892 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_174
timestamp -7200
transform 1 0 16560 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_186
timestamp -7200
transform 1 0 17664 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp -7200
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_197
timestamp -7200
transform 1 0 18676 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_214
timestamp -7200
transform 1 0 20240 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_219
timestamp -7200
transform 1 0 20700 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_225
timestamp -7200
transform 1 0 21252 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_249
timestamp -7200
transform 1 0 23460 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_253
timestamp -7200
transform 1 0 23828 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_263
timestamp -7200
transform 1 0 24748 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_270
timestamp -7200
transform 1 0 25392 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_282
timestamp -7200
transform 1 0 26496 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_288
timestamp -7200
transform 1 0 27048 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp -7200
transform 1 0 828 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_11
timestamp -7200
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_36
timestamp -7200
transform 1 0 3864 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_44
timestamp -7200
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp -7200
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_67
timestamp -7200
transform 1 0 6716 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_81
timestamp -7200
transform 1 0 8004 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_108
timestamp -7200
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp -7200
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_125
timestamp -7200
transform 1 0 12052 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_134
timestamp -7200
transform 1 0 12880 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_138
timestamp -7200
transform 1 0 13248 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_177
timestamp -7200
transform 1 0 16836 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp -7200
transform 1 0 21068 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_225
timestamp -7200
transform 1 0 21252 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_239
timestamp -7200
transform 1 0 22540 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_249
timestamp -7200
transform 1 0 23460 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_277
timestamp -7200
transform 1 0 26036 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp -7200
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp -7200
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp -7200
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp -7200
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_73
timestamp -7200
transform 1 0 7268 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp -7200
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_89
timestamp -7200
transform 1 0 8740 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_114
timestamp -7200
transform 1 0 11040 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_126
timestamp -7200
transform 1 0 12144 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp -7200
transform 1 0 13156 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_141
timestamp -7200
transform 1 0 13524 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_156
timestamp -7200
transform 1 0 14904 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_165
timestamp -7200
transform 1 0 15732 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_190
timestamp -7200
transform 1 0 18032 0 1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_217
timestamp -7200
transform 1 0 20516 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_229
timestamp -7200
transform 1 0 21620 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_239
timestamp -7200
transform 1 0 22540 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp -7200
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_267
timestamp -7200
transform 1 0 25116 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_284
timestamp -7200
transform 1 0 26680 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_288
timestamp -7200
transform 1 0 27048 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp -7200
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp -7200
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_27
timestamp -7200
transform 1 0 3036 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_34
timestamp -7200
transform 1 0 3680 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_42
timestamp -7200
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_48
timestamp -7200
transform 1 0 4968 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp -7200
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_113
timestamp -7200
transform 1 0 10948 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_119
timestamp -7200
transform 1 0 11500 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_164
timestamp -7200
transform 1 0 15640 0 -1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp -7200
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_181
timestamp -7200
transform 1 0 17204 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_220
timestamp -7200
transform 1 0 20792 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_233
timestamp -7200
transform 1 0 21988 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_238
timestamp -7200
transform 1 0 22448 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_257
timestamp -7200
transform 1 0 24196 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_263
timestamp -7200
transform 1 0 24748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp -7200
transform 1 0 828 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_11
timestamp -7200
transform 1 0 1564 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp -7200
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp -7200
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_53
timestamp -7200
transform 1 0 5428 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_61
timestamp -7200
transform 1 0 6164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp -7200
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_92
timestamp -7200
transform 1 0 9016 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_130
timestamp -7200
transform 1 0 12512 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_149
timestamp -7200
transform 1 0 14260 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_174
timestamp -7200
transform 1 0 16560 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_184
timestamp -7200
transform 1 0 17480 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_193
timestamp -7200
transform 1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_213
timestamp -7200
transform 1 0 20148 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_221
timestamp -7200
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp -7200
transform 1 0 23644 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_261
timestamp -7200
transform 1 0 24564 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_288
timestamp -7200
transform 1 0 27048 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp -7200
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_15
timestamp -7200
transform 1 0 1932 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_41
timestamp -7200
transform 1 0 4324 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_45
timestamp -7200
transform 1 0 4692 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp -7200
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_57
timestamp -7200
transform 1 0 5796 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_65
timestamp -7200
transform 1 0 6532 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_89
timestamp -7200
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_109
timestamp -7200
transform 1 0 10580 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_134
timestamp -7200
transform 1 0 12880 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_138
timestamp -7200
transform 1 0 13248 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_172
timestamp -7200
transform 1 0 16376 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_186
timestamp -7200
transform 1 0 17664 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_194
timestamp -7200
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_220
timestamp -7200
transform 1 0 20792 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_225
timestamp -7200
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_254
timestamp -7200
transform 1 0 23920 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_262
timestamp -7200
transform 1 0 24656 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp -7200
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_3
timestamp -7200
transform 1 0 828 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_46
timestamp -7200
transform 1 0 4784 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_63
timestamp -7200
transform 1 0 6348 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_71
timestamp -7200
transform 1 0 7084 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp -7200
transform 1 0 8004 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_89
timestamp -7200
transform 1 0 8740 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_103
timestamp -7200
transform 1 0 10028 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_111
timestamp -7200
transform 1 0 10764 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_116
timestamp -7200
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_128
timestamp -7200
transform 1 0 12328 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_141
timestamp -7200
transform 1 0 13524 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_169
timestamp -7200
transform 1 0 16100 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_173
timestamp -7200
transform 1 0 16468 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_190
timestamp -7200
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_225
timestamp -7200
transform 1 0 21252 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp -7200
transform 1 0 23460 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_285
timestamp -7200
transform 1 0 26772 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp -7200
transform 1 0 828 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_11
timestamp -7200
transform 1 0 1564 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_38
timestamp -7200
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_46
timestamp -7200
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_60
timestamp -7200
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_68
timestamp -7200
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_91
timestamp -7200
transform 1 0 8924 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_103
timestamp -7200
transform 1 0 10028 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_113
timestamp -7200
transform 1 0 10948 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_122
timestamp -7200
transform 1 0 11776 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_130
timestamp -7200
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_140
timestamp -7200
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_150
timestamp -7200
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_177
timestamp -7200
transform 1 0 16836 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_198
timestamp -7200
transform 1 0 18768 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_225
timestamp -7200
transform 1 0 21252 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_245
timestamp -7200
transform 1 0 23092 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp -7200
transform 1 0 25668 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp -7200
transform 1 0 26220 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_3
timestamp -7200
transform 1 0 828 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_9
timestamp -7200
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp -7200
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_42
timestamp -7200
transform 1 0 4416 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_48
timestamp -7200
transform 1 0 4968 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_55
timestamp -7200
transform 1 0 5612 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_64
timestamp -7200
transform 1 0 6440 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_72
timestamp -7200
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_85
timestamp -7200
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_94
timestamp -7200
transform 1 0 9200 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_100
timestamp -7200
transform 1 0 9752 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_125
timestamp -7200
transform 1 0 12052 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp -7200
transform 1 0 13156 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_141
timestamp -7200
transform 1 0 13524 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_145
timestamp -7200
transform 1 0 13892 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_170
timestamp -7200
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp -7200
transform 1 0 23092 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp -7200
transform 1 0 23644 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_253
timestamp -7200
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_263
timestamp -7200
transform 1 0 24748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_288
timestamp -7200
transform 1 0 27048 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_3
timestamp -7200
transform 1 0 828 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_11
timestamp -7200
transform 1 0 1564 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp -7200
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp -7200
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_61
timestamp -7200
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_70
timestamp -7200
transform 1 0 6992 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_78
timestamp -7200
transform 1 0 7728 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_107
timestamp -7200
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_118
timestamp -7200
transform 1 0 11408 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_128
timestamp -7200
transform 1 0 12328 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_136
timestamp -7200
transform 1 0 13064 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_181
timestamp -7200
transform 1 0 17204 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_192
timestamp -7200
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_221
timestamp -7200
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_257
timestamp -7200
transform 1 0 24196 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_263
timestamp -7200
transform 1 0 24748 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp -7200
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_15
timestamp -7200
transform 1 0 1932 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_21
timestamp -7200
transform 1 0 2484 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_37
timestamp -7200
transform 1 0 3956 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp -7200
transform 1 0 8372 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_93
timestamp -7200
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_118
timestamp -7200
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_123
timestamp -7200
transform 1 0 11868 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_141
timestamp -7200
transform 1 0 13524 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_163
timestamp -7200
transform 1 0 15548 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_180
timestamp -7200
transform 1 0 17112 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_184
timestamp -7200
transform 1 0 17480 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp -7200
transform 1 0 18308 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_221
timestamp -7200
transform 1 0 20884 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_248
timestamp -7200
transform 1 0 23368 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_269
timestamp -7200
transform 1 0 25300 0 1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp -7200
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp -7200
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp -7200
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_39
timestamp -7200
transform 1 0 4140 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_47
timestamp -7200
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_74
timestamp -7200
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_86
timestamp -7200
transform 1 0 8464 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_90
timestamp -7200
transform 1 0 8832 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_102
timestamp -7200
transform 1 0 9936 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_108
timestamp -7200
transform 1 0 10488 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_126
timestamp -7200
transform 1 0 12144 0 -1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_155
timestamp -7200
transform 1 0 14812 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp -7200
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp -7200
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_221
timestamp -7200
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_225
timestamp -7200
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_258
timestamp -7200
transform 1 0 24288 0 -1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp -7200
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp -7200
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp -7200
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp -7200
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp -7200
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_53
timestamp -7200
transform 1 0 5428 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_61
timestamp -7200
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_73
timestamp -7200
transform 1 0 7268 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp -7200
transform 1 0 8004 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_85
timestamp -7200
transform 1 0 8372 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_116
timestamp -7200
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_122
timestamp -7200
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_128
timestamp -7200
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_149
timestamp -7200
transform 1 0 14260 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_154
timestamp -7200
transform 1 0 14720 0 1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_162
timestamp -7200
transform 1 0 15456 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_174
timestamp -7200
transform 1 0 16560 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_180
timestamp -7200
transform 1 0 17112 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp -7200
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp -7200
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_221
timestamp -7200
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_247
timestamp -7200
transform 1 0 23276 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp -7200
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_277
timestamp -7200
transform 1 0 26036 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_286
timestamp -7200
transform 1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp -7200
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp -7200
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp -7200
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp -7200
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp -7200
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp -7200
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_57
timestamp -7200
transform 1 0 5796 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_63
timestamp -7200
transform 1 0 6348 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_103
timestamp -7200
transform 1 0 10028 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_129
timestamp -7200
transform 1 0 12420 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_169
timestamp -7200
transform 1 0 16100 0 -1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_179
timestamp -7200
transform 1 0 17020 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_191
timestamp -7200
transform 1 0 18124 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_202
timestamp -7200
transform 1 0 19136 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_219
timestamp -7200
transform 1 0 20700 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp -7200
transform 1 0 21068 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_225
timestamp -7200
transform 1 0 21252 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_251
timestamp -7200
transform 1 0 23644 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_255
timestamp -7200
transform 1 0 24012 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_264
timestamp -7200
transform 1 0 24840 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_273
timestamp -7200
transform 1 0 25668 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_6
timestamp -7200
transform 1 0 1104 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_13
timestamp -7200
transform 1 0 1748 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_21
timestamp -7200
transform 1 0 2484 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp -7200
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_29
timestamp -7200
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_34
timestamp -7200
transform 1 0 3680 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_41
timestamp -7200
transform 1 0 4324 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_48
timestamp -7200
transform 1 0 4968 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_55
timestamp -7200
transform 1 0 5612 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_57
timestamp -7200
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_62
timestamp -7200
transform 1 0 6256 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_69
timestamp -7200
transform 1 0 6900 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_77
timestamp -7200
transform 1 0 7636 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_85
timestamp -7200
transform 1 0 8372 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_93
timestamp -7200
transform 1 0 9108 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_97
timestamp -7200
transform 1 0 9476 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_106
timestamp -7200
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_113
timestamp -7200
transform 1 0 10948 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_121
timestamp -7200
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_127
timestamp -7200
transform 1 0 12236 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp -7200
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_141
timestamp -7200
transform 1 0 13524 0 1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_151
timestamp -7200
transform 1 0 14444 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_163
timestamp -7200
transform 1 0 15548 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_167
timestamp -7200
transform 1 0 15916 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_169
timestamp -7200
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_174
timestamp -7200
transform 1 0 16560 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_182
timestamp -7200
transform 1 0 17296 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_188
timestamp -7200
transform 1 0 17848 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_192
timestamp -7200
transform 1 0 18216 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_240
timestamp -7200
transform 1 0 22632 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_244
timestamp -7200
transform 1 0 23000 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp -7200
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_253
timestamp -7200
transform 1 0 23828 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_258
timestamp -7200
transform 1 0 24288 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_265
timestamp -7200
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp -7200
transform 1 0 10120 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp -7200
transform -1 0 13340 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp -7200
transform -1 0 12604 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp -7200
transform -1 0 19412 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp -7200
transform -1 0 18216 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp -7200
transform -1 0 10028 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp -7200
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp -7200
transform 1 0 20148 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp -7200
transform -1 0 20148 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp -7200
transform -1 0 12604 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp -7200
transform 1 0 18400 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp -7200
transform -1 0 20148 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp -7200
transform -1 0 8280 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp -7200
transform -1 0 20700 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp -7200
transform -1 0 20884 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp -7200
transform -1 0 16836 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp -7200
transform -1 0 16008 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp -7200
transform 1 0 17204 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp -7200
transform 1 0 24840 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp -7200
transform -1 0 25668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp -7200
transform -1 0 20792 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp -7200
transform -1 0 20056 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp -7200
transform -1 0 13156 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp -7200
transform -1 0 23644 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp -7200
transform -1 0 22172 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp -7200
transform -1 0 25300 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp -7200
transform 1 0 25116 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp -7200
transform -1 0 14812 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp -7200
transform 1 0 16928 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp -7200
transform -1 0 6532 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp -7200
transform -1 0 23276 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp -7200
transform -1 0 22080 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp -7200
transform -1 0 20516 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp -7200
transform -1 0 19688 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp -7200
transform -1 0 26036 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp -7200
transform -1 0 25668 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp -7200
transform 1 0 26128 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp -7200
transform -1 0 27140 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp -7200
transform 1 0 21344 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp -7200
transform -1 0 23368 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp -7200
transform -1 0 24288 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp -7200
transform -1 0 21068 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp -7200
transform 1 0 18124 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp -7200
transform -1 0 24196 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp -7200
transform -1 0 27140 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp -7200
transform -1 0 24564 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp -7200
transform -1 0 24564 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp -7200
transform -1 0 27140 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp -7200
transform -1 0 15548 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp -7200
transform -1 0 14352 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp -7200
transform -1 0 23552 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp -7200
transform -1 0 23092 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp -7200
transform -1 0 4876 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp -7200
transform -1 0 3956 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp -7200
transform -1 0 21252 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp -7200
transform 1 0 26404 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp -7200
transform 1 0 14996 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp -7200
transform -1 0 16836 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp -7200
transform -1 0 16008 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp -7200
transform -1 0 17112 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp -7200
transform 1 0 20976 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp -7200
transform 1 0 19412 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp -7200
transform -1 0 7268 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp -7200
transform -1 0 18032 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp -7200
transform -1 0 18032 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp -7200
transform -1 0 27048 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp -7200
transform -1 0 27140 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp -7200
transform -1 0 18676 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp -7200
transform -1 0 27140 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp -7200
transform -1 0 3772 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp -7200
transform -1 0 10856 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp -7200
transform -1 0 14260 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp -7200
transform 1 0 11592 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp -7200
transform 1 0 5796 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp -7200
transform -1 0 27140 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp -7200
transform -1 0 10304 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp -7200
transform -1 0 5060 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp -7200
transform -1 0 22448 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp -7200
transform -1 0 4600 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp -7200
transform 1 0 3128 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp -7200
transform -1 0 3036 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp -7200
transform -1 0 27140 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp -7200
transform -1 0 3680 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp -7200
transform -1 0 3956 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp -7200
transform 1 0 7268 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp -7200
transform 1 0 7544 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp -7200
transform -1 0 7728 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp -7200
transform 1 0 11408 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp -7200
transform 1 0 7820 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp -7200
transform -1 0 14260 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp -7200
transform 1 0 12420 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp -7200
transform 1 0 8648 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp -7200
transform -1 0 3496 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp -7200
transform 1 0 8004 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp -7200
transform -1 0 24564 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp -7200
transform -1 0 18860 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp -7200
transform -1 0 12052 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp -7200
transform 1 0 7268 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp -7200
transform -1 0 25024 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp -7200
transform -1 0 18124 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp -7200
transform -1 0 16836 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp -7200
transform -1 0 13432 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp -7200
transform 1 0 26404 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp -7200
transform -1 0 26312 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp -7200
transform 1 0 25392 0 1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp -7200
transform 1 0 25116 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -7200
transform 1 0 24656 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp -7200
transform 1 0 24012 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp -7200
transform 1 0 23368 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp -7200
transform 1 0 22724 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp -7200
transform 1 0 22356 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp -7200
transform 1 0 20884 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp -7200
transform -1 0 18584 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp -7200
transform 1 0 17572 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input12
timestamp -7200
transform 1 0 16928 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input13
timestamp -7200
transform -1 0 16560 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_31
timestamp -7200
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -7200
transform -1 0 27416 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_32
timestamp -7200
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -7200
transform -1 0 27416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_33
timestamp -7200
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -7200
transform -1 0 27416 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_34
timestamp -7200
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -7200
transform -1 0 27416 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_35
timestamp -7200
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -7200
transform -1 0 27416 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_36
timestamp -7200
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -7200
transform -1 0 27416 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_37
timestamp -7200
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -7200
transform -1 0 27416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_38
timestamp -7200
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -7200
transform -1 0 27416 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_39
timestamp -7200
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -7200
transform -1 0 27416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_40
timestamp -7200
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -7200
transform -1 0 27416 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_41
timestamp -7200
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -7200
transform -1 0 27416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_42
timestamp -7200
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -7200
transform -1 0 27416 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_43
timestamp -7200
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -7200
transform -1 0 27416 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_44
timestamp -7200
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -7200
transform -1 0 27416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_45
timestamp -7200
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -7200
transform -1 0 27416 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_46
timestamp -7200
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -7200
transform -1 0 27416 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_47
timestamp -7200
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -7200
transform -1 0 27416 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_48
timestamp -7200
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -7200
transform -1 0 27416 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_49
timestamp -7200
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -7200
transform -1 0 27416 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_50
timestamp -7200
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -7200
transform -1 0 27416 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_51
timestamp -7200
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -7200
transform -1 0 27416 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_52
timestamp -7200
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -7200
transform -1 0 27416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_53
timestamp -7200
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -7200
transform -1 0 27416 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_54
timestamp -7200
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -7200
transform -1 0 27416 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_55
timestamp -7200
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -7200
transform -1 0 27416 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_56
timestamp -7200
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -7200
transform -1 0 27416 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_57
timestamp -7200
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -7200
transform -1 0 27416 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_58
timestamp -7200
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -7200
transform -1 0 27416 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_59
timestamp -7200
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -7200
transform -1 0 27416 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_60
timestamp -7200
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -7200
transform -1 0 27416 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_61
timestamp -7200
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -7200
transform -1 0 27416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp -7200
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp -7200
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp -7200
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp -7200
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp -7200
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp -7200
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68
timestamp -7200
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp -7200
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp -7200
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp -7200
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_72
timestamp -7200
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_73
timestamp -7200
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_74
timestamp -7200
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_75
timestamp -7200
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_76
timestamp -7200
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_77
timestamp -7200
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_78
timestamp -7200
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_79
timestamp -7200
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_80
timestamp -7200
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_81
timestamp -7200
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_82
timestamp -7200
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_83
timestamp -7200
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_84
timestamp -7200
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_85
timestamp -7200
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_86
timestamp -7200
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_87
timestamp -7200
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_88
timestamp -7200
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_89
timestamp -7200
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_90
timestamp -7200
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_91
timestamp -7200
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_92
timestamp -7200
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_93
timestamp -7200
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_94
timestamp -7200
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_95
timestamp -7200
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_96
timestamp -7200
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_97
timestamp -7200
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_98
timestamp -7200
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_99
timestamp -7200
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_100
timestamp -7200
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_101
timestamp -7200
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_102
timestamp -7200
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_103
timestamp -7200
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_104
timestamp -7200
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_105
timestamp -7200
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_106
timestamp -7200
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_107
timestamp -7200
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_108
timestamp -7200
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_109
timestamp -7200
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_110
timestamp -7200
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_111
timestamp -7200
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_112
timestamp -7200
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_113
timestamp -7200
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_114
timestamp -7200
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_115
timestamp -7200
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_116
timestamp -7200
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_117
timestamp -7200
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_118
timestamp -7200
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_119
timestamp -7200
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_120
timestamp -7200
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_121
timestamp -7200
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_122
timestamp -7200
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_123
timestamp -7200
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_124
timestamp -7200
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_125
timestamp -7200
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_126
timestamp -7200
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_127
timestamp -7200
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_128
timestamp -7200
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_129
timestamp -7200
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_130
timestamp -7200
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_131
timestamp -7200
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_132
timestamp -7200
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_133
timestamp -7200
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_134
timestamp -7200
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_135
timestamp -7200
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_136
timestamp -7200
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_137
timestamp -7200
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_138
timestamp -7200
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_139
timestamp -7200
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_140
timestamp -7200
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_141
timestamp -7200
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_142
timestamp -7200
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_143
timestamp -7200
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_144
timestamp -7200
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_145
timestamp -7200
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_146
timestamp -7200
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_147
timestamp -7200
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_148
timestamp -7200
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_149
timestamp -7200
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_150
timestamp -7200
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_151
timestamp -7200
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_152
timestamp -7200
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_153
timestamp -7200
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_154
timestamp -7200
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_155
timestamp -7200
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_156
timestamp -7200
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_157
timestamp -7200
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_158
timestamp -7200
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_159
timestamp -7200
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_160
timestamp -7200
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp -7200
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_162
timestamp -7200
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_163
timestamp -7200
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp -7200
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp -7200
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_166
timestamp -7200
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_167
timestamp -7200
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp -7200
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp -7200
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_170
timestamp -7200
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_171
timestamp -7200
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_172
timestamp -7200
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_173
timestamp -7200
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_174
timestamp -7200
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_175
timestamp -7200
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_176
timestamp -7200
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_177
timestamp -7200
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_178
timestamp -7200
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_179
timestamp -7200
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_180
timestamp -7200
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_181
timestamp -7200
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_182
timestamp -7200
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_183
timestamp -7200
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_184
timestamp -7200
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_185
timestamp -7200
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_186
timestamp -7200
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_187
timestamp -7200
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_188
timestamp -7200
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_189
timestamp -7200
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_190
timestamp -7200
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_191
timestamp -7200
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_192
timestamp -7200
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_193
timestamp -7200
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_194
timestamp -7200
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_195
timestamp -7200
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_196
timestamp -7200
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_197
timestamp -7200
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_198
timestamp -7200
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_199
timestamp -7200
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_200
timestamp -7200
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_201
timestamp -7200
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_202
timestamp -7200
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_203
timestamp -7200
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_204
timestamp -7200
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_205
timestamp -7200
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_206
timestamp -7200
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_207
timestamp -7200
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_208
timestamp -7200
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_209
timestamp -7200
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_210
timestamp -7200
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_211
timestamp -7200
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_212
timestamp -7200
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_213
timestamp -7200
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_214
timestamp -7200
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_215
timestamp -7200
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_216
timestamp -7200
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_217
timestamp -7200
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_218
timestamp -7200
transform 1 0 5704 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_219
timestamp -7200
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_220
timestamp -7200
transform 1 0 10856 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_221
timestamp -7200
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_222
timestamp -7200
transform 1 0 16008 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_223
timestamp -7200
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_224
timestamp -7200
transform 1 0 21160 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_225
timestamp -7200
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_226
timestamp -7200
transform 1 0 26312 0 1 16864
box -38 -48 130 592
<< labels >>
rlabel metal2 s 14064 16864 14064 16864 4 VGND
rlabel metal1 s 13984 17408 13984 17408 4 VPWR
rlabel metal1 s 11990 14858 11990 14858 4 _000_
rlabel metal2 s 6394 15062 6394 15062 4 _001_
rlabel metal1 s 10856 13498 10856 13498 4 _002_
rlabel metal1 s 7314 12954 7314 12954 4 _003_
rlabel metal1 s 5274 14858 5274 14858 4 _004_
rlabel metal1 s 3450 9010 3450 9010 4 _005_
rlabel metal2 s 2898 9894 2898 9894 4 _006_
rlabel metal2 s 1705 9146 1705 9146 4 _007_
rlabel metal1 s 2622 8024 2622 8024 4 _008_
rlabel metal2 s 2070 6630 2070 6630 4 _009_
rlabel metal1 s 4043 6154 4043 6154 4 _010_
rlabel metal1 s 5290 5542 5290 5542 4 _011_
rlabel metal1 s 17188 6154 17188 6154 4 _012_
rlabel metal2 s 21026 5134 21026 5134 4 _013_
rlabel metal2 s 19458 5984 19458 5984 4 _014_
rlabel metal1 s 18073 7242 18073 7242 4 _015_
rlabel metal1 s 22852 5746 22852 5746 4 _016_
rlabel metal2 s 22862 4454 22862 4454 4 _017_
rlabel metal1 s 24886 5134 24886 5134 4 _018_
rlabel metal1 s 25571 6222 25571 6222 4 _019_
rlabel metal1 s 25438 7514 25438 7514 4 _020_
rlabel metal1 s 25479 8330 25479 8330 4 _021_
rlabel metal2 s 22126 7038 22126 7038 4 _022_
rlabel metal1 s 24568 9078 24568 9078 4 _023_
rlabel metal2 s 22218 9010 22218 9010 4 _024_
rlabel metal2 s 19545 8398 19545 8398 4 _025_
rlabel metal2 s 16785 9010 16785 9010 4 _026_
rlabel metal1 s 15916 10234 15916 10234 4 _027_
rlabel metal2 s 12466 15844 12466 15844 4 _028_
rlabel metal2 s 8510 16422 8510 16422 4 _029_
rlabel metal1 s 7355 16694 7355 16694 4 _030_
rlabel metal2 s 11178 16286 11178 16286 4 _031_
rlabel metal2 s 3266 14246 3266 14246 4 _032_
rlabel metal2 s 1789 13770 1789 13770 4 _033_
rlabel metal1 s 1881 12682 1881 12682 4 _034_
rlabel metal1 s 2157 11594 2157 11594 4 _035_
rlabel metal1 s 5239 12682 5239 12682 4 _036_
rlabel metal2 s 12098 12070 12098 12070 4 _037_
rlabel metal1 s 9609 11254 9609 11254 4 _038_
rlabel metal1 s 9690 10506 9690 10506 4 _039_
rlabel metal1 s 9236 10098 9236 10098 4 _040_
rlabel metal1 s 9782 9418 9782 9418 4 _041_
rlabel metal2 s 13841 7310 13841 7310 4 _042_
rlabel metal2 s 11357 7242 11357 7242 4 _043_
rlabel metal1 s 13197 7990 13197 7990 4 _044_
rlabel metal2 s 11914 8704 11914 8704 4 _045_
rlabel metal1 s 12604 10778 12604 10778 4 _046_
rlabel metal1 s 19504 13362 19504 13362 4 _047_
rlabel metal2 s 20005 13362 20005 13362 4 _048_
rlabel metal1 s 22862 13838 22862 13838 4 _049_
rlabel metal2 s 25254 13124 25254 13124 4 _050_
rlabel metal2 s 25617 12682 25617 12682 4 _051_
rlabel metal1 s 26680 14994 26680 14994 4 _052_
rlabel metal1 s 25387 15606 25387 15606 4 _053_
rlabel metal1 s 25530 16660 25530 16660 4 _054_
rlabel metal1 s 22126 16627 22126 16627 4 _055_
rlabel metal2 s 20746 16388 20746 16388 4 _056_
rlabel metal1 s 19688 15470 19688 15470 4 _057_
rlabel metal1 s 16647 14858 16647 14858 4 _058_
rlabel metal1 s 15548 14382 15548 14382 4 _059_
rlabel metal1 s 14122 14586 14122 14586 4 _060_
rlabel metal2 s 14393 12750 14393 12750 4 _061_
rlabel metal1 s 6527 11254 6527 11254 4 _062_
rlabel metal1 s 5704 9554 5704 9554 4 _063_
rlabel metal1 s 6072 10234 6072 10234 4 _064_
rlabel metal1 s 7268 8058 7268 8058 4 _065_
rlabel metal2 s 6849 7310 6849 7310 4 _066_
rlabel metal1 s 8045 6834 8045 6834 4 _067_
rlabel metal1 s 10948 6290 10948 6290 4 _068_
rlabel metal2 s 16058 8398 16058 8398 4 _069_
rlabel metal2 s 16698 10268 16698 10268 4 _070_
rlabel metal1 s 18630 9690 18630 9690 4 _071_
rlabel metal1 s 19596 11118 19596 11118 4 _072_
rlabel metal2 s 21298 11764 21298 11764 4 _073_
rlabel metal1 s 24012 10642 24012 10642 4 _074_
rlabel metal1 s 25295 11662 25295 11662 4 _075_
rlabel metal1 s 25668 10234 25668 10234 4 _076_
rlabel metal2 s 24702 10234 24702 10234 4 _077_
rlabel metal1 s 23812 14858 23812 14858 4 _078_
rlabel metal1 s 22540 14586 22540 14586 4 _079_
rlabel metal1 s 22310 13804 22310 13804 4 _080_
rlabel metal2 s 20194 14484 20194 14484 4 _081_
rlabel metal1 s 17894 13498 17894 13498 4 _082_
rlabel metal1 s 17346 12682 17346 12682 4 _083_
rlabel metal1 s 13616 11866 13616 11866 4 _084_
rlabel metal2 s 14950 6018 14950 6018 4 _085_
rlabel metal1 s 9563 2890 9563 2890 4 _086_
rlabel metal1 s 4641 3978 4641 3978 4 _087_
rlabel metal1 s 3756 3638 3756 3638 4 _088_
rlabel metal1 s 5561 5066 5561 5066 4 _089_
rlabel metal1 s 6803 3638 6803 3638 4 _090_
rlabel metal2 s 8597 3570 8597 3570 4 _091_
rlabel metal1 s 11495 3638 11495 3638 4 _092_
rlabel metal2 s 11638 5270 11638 5270 4 _093_
rlabel metal2 s 8694 6018 8694 6018 4 _094_
rlabel metal1 s 10012 1802 10012 1802 4 _095_
rlabel metal1 s 6220 1870 6220 1870 4 _096_
rlabel metal2 s 4370 2278 4370 2278 4 _097_
rlabel metal2 s 3629 2958 3629 2958 4 _098_
rlabel metal2 s 7585 1394 7585 1394 4 _099_
rlabel metal1 s 9368 1462 9368 1462 4 _100_
rlabel metal1 s 13068 1462 13068 1462 4 _101_
rlabel metal2 s 12742 2686 12742 2686 4 _102_
rlabel metal1 s 15466 782 15466 782 4 _103_
rlabel metal1 s 17070 1802 17070 1802 4 _104_
rlabel metal2 s 17061 1462 17061 1462 4 _105_
rlabel metal1 s 17608 4658 17608 4658 4 _106_
rlabel metal1 s 18768 3706 18768 3706 4 _107_
rlabel metal1 s 19166 3638 19166 3638 4 _108_
rlabel metal1 s 18752 2890 18752 2890 4 _109_
rlabel metal1 s 18706 4726 18706 4726 4 _110_
rlabel metal1 s 15134 15878 15134 15878 4 _111_
rlabel metal1 s 14122 11220 14122 11220 4 _112_
rlabel metal1 s 14766 9996 14766 9996 4 _113_
rlabel metal1 s 2162 9962 2162 9962 4 _114_
rlabel metal2 s 2714 13600 2714 13600 4 _115_
rlabel metal2 s 12650 15810 12650 15810 4 _116_
rlabel metal2 s 10994 15708 10994 15708 4 _117_
rlabel metal2 s 13386 16218 13386 16218 4 _118_
rlabel metal1 s 11638 14960 11638 14960 4 _119_
rlabel metal1 s 4094 13158 4094 13158 4 _120_
rlabel metal1 s 5152 13702 5152 13702 4 _121_
rlabel metal2 s 9890 14093 9890 14093 4 _122_
rlabel metal1 s 7268 14926 7268 14926 4 _123_
rlabel metal1 s 7268 15946 7268 15946 4 _124_
rlabel metal1 s 6946 15878 6946 15878 4 _125_
rlabel metal2 s 7590 12954 7590 12954 4 _126_
rlabel metal1 s 7728 12886 7728 12886 4 _127_
rlabel metal1 s 8786 12750 8786 12750 4 _128_
rlabel metal1 s 21942 13872 21942 13872 4 _129_
rlabel metal1 s 11454 12954 11454 12954 4 _130_
rlabel metal1 s 15525 13838 15525 13838 4 _131_
rlabel metal2 s 13567 9010 13567 9010 4 _132_
rlabel metal1 s 10358 13770 10358 13770 4 _133_
rlabel metal1 s 10350 13396 10350 13396 4 _134_
rlabel metal1 s 10672 14790 10672 14790 4 _135_
rlabel metal1 s 13478 16728 13478 16728 4 _136_
rlabel metal1 s 18722 1394 18722 1394 4 _137_
rlabel metal1 s 15502 1394 15502 1394 4 _138_
rlabel metal1 s 12742 680 12742 680 4 _139_
rlabel metal2 s 16146 833 16146 833 4 _140_
rlabel metal2 s 18906 1632 18906 1632 4 _141_
rlabel metal3 s 18998 1411 18998 1411 4 _142_
rlabel metal1 s 22494 1394 22494 1394 4 _143_
rlabel metal3 s 20286 1955 20286 1955 4 _144_
rlabel metal1 s 20516 1326 20516 1326 4 _145_
rlabel metal1 s 20194 884 20194 884 4 _146_
rlabel metal2 s 15594 9010 15594 9010 4 _147_
rlabel metal2 s 18466 1394 18466 1394 4 _148_
rlabel metal3 s 14674 2635 14674 2635 4 _149_
rlabel metal1 s 15640 16626 15640 16626 4 _150_
rlabel metal1 s 15824 3162 15824 3162 4 _151_
rlabel metal1 s 15088 11798 15088 11798 4 _152_
rlabel metal1 s 14582 3706 14582 3706 4 _153_
rlabel metal1 s 15272 16626 15272 16626 4 _154_
rlabel metal1 s 14536 5338 14536 5338 4 _155_
rlabel metal1 s 14490 17102 14490 17102 4 _156_
rlabel metal1 s 13846 3706 13846 3706 4 _157_
rlabel metal1 s 13202 10234 13202 10234 4 _158_
rlabel metal1 s 13294 4250 13294 4250 4 _159_
rlabel metal1 s 8142 4624 8142 4624 4 _160_
rlabel metal1 s 11776 16082 11776 16082 4 _161_
rlabel metal2 s 12650 4624 12650 4624 4 _162_
rlabel metal2 s 11914 14761 11914 14761 4 _163_
rlabel metal2 s 13570 5712 13570 5712 4 _164_
rlabel metal2 s 11500 14212 11500 14212 4 _165_
rlabel metal2 s 4554 6698 4554 6698 4 _166_
rlabel metal1 s 9338 2448 9338 2448 4 _167_
rlabel metal2 s 17158 9265 17158 9265 4 _168_
rlabel metal1 s 4324 9010 4324 9010 4 _169_
rlabel metal2 s 4646 9180 4646 9180 4 _170_
rlabel metal2 s 2070 9010 2070 9010 4 _171_
rlabel metal1 s 3818 9622 3818 9622 4 _172_
rlabel metal2 s 3082 9690 3082 9690 4 _173_
rlabel metal2 s 2346 6562 2346 6562 4 _174_
rlabel metal1 s 1610 8976 1610 8976 4 _175_
rlabel metal1 s 3726 7378 3726 7378 4 _176_
rlabel metal2 s 3450 7752 3450 7752 4 _177_
rlabel metal2 s 2438 7718 2438 7718 4 _178_
rlabel metal1 s 2392 6222 2392 6222 4 _179_
rlabel metal1 s 2070 6188 2070 6188 4 _180_
rlabel metal2 s 4278 6188 4278 6188 4 _181_
rlabel metal1 s 4278 7276 4278 7276 4 _182_
rlabel metal1 s 19458 7174 19458 7174 4 _183_
rlabel metal1 s 5382 5780 5382 5780 4 _184_
rlabel metal2 s 20562 6494 20562 6494 4 _185_
rlabel metal1 s 17204 5882 17204 5882 4 _186_
rlabel metal1 s 21666 5848 21666 5848 4 _187_
rlabel metal2 s 21482 5814 21482 5814 4 _188_
rlabel metal1 s 21052 5814 21052 5814 4 _189_
rlabel metal1 s 21206 5746 21206 5746 4 _190_
rlabel metal1 s 19274 5066 19274 5066 4 _191_
rlabel metal2 s 18630 5916 18630 5916 4 _192_
rlabel metal1 s 19688 7174 19688 7174 4 _193_
rlabel metal1 s 18308 6766 18308 6766 4 _194_
rlabel metal1 s 18630 6970 18630 6970 4 _195_
rlabel metal1 s 23138 4998 23138 4998 4 _196_
rlabel metal2 s 22586 5916 22586 5916 4 _197_
rlabel metal1 s 23138 5338 23138 5338 4 _198_
rlabel metal1 s 23752 5066 23752 5066 4 _199_
rlabel metal1 s 23368 4046 23368 4046 4 _200_
rlabel metal2 s 24334 5338 24334 5338 4 _201_
rlabel metal1 s 25070 6834 25070 6834 4 _202_
rlabel metal2 s 24978 6528 24978 6528 4 _203_
rlabel metal1 s 21344 8058 21344 8058 4 _204_
rlabel metal2 s 25806 7140 25806 7140 4 _205_
rlabel metal1 s 24840 7310 24840 7310 4 _206_
rlabel metal1 s 21482 8942 21482 8942 4 _207_
rlabel metal2 s 25346 7514 25346 7514 4 _208_
rlabel metal1 s 24242 8602 24242 8602 4 _209_
rlabel metal2 s 22218 7072 22218 7072 4 _210_
rlabel metal1 s 22256 6154 22256 6154 4 _211_
rlabel metal1 s 21758 6426 21758 6426 4 _212_
rlabel metal1 s 21850 8432 21850 8432 4 _213_
rlabel metal2 s 22770 8840 22770 8840 4 _214_
rlabel metal1 s 23368 8602 23368 8602 4 _215_
rlabel metal1 s 21298 9044 21298 9044 4 _216_
rlabel metal1 s 21712 8398 21712 8398 4 _217_
rlabel metal1 s 19780 7786 19780 7786 4 _218_
rlabel metal1 s 20424 8058 20424 8058 4 _219_
rlabel metal2 s 20102 8398 20102 8398 4 _220_
rlabel metal1 s 17112 8398 17112 8398 4 _221_
rlabel metal1 s 17618 9962 17618 9962 4 _222_
rlabel metal1 s 16652 9622 16652 9622 4 _223_
rlabel metal1 s 10810 15062 10810 15062 4 _224_
rlabel metal2 s 9890 15436 9890 15436 4 _225_
rlabel metal2 s 8786 15844 8786 15844 4 _226_
rlabel metal1 s 11592 14586 11592 14586 4 _227_
rlabel metal1 s 8970 16048 8970 16048 4 _228_
rlabel metal1 s 10810 16082 10810 16082 4 _229_
rlabel metal1 s 9936 16218 9936 16218 4 _230_
rlabel metal2 s 19458 10914 19458 10914 4 _231_
rlabel metal1 s 14122 12648 14122 12648 4 _232_
rlabel metal1 s 10810 14586 10810 14586 4 _233_
rlabel metal1 s 10534 16150 10534 16150 4 _234_
rlabel metal1 s 4876 14382 4876 14382 4 _235_
rlabel metal1 s 8694 14450 8694 14450 4 _236_
rlabel metal1 s 7912 14994 7912 14994 4 _237_
rlabel metal1 s 9798 15062 9798 15062 4 _238_
rlabel metal2 s 9062 14620 9062 14620 4 _239_
rlabel metal1 s 6348 14518 6348 14518 4 _240_
rlabel metal1 s 3818 13430 3818 13430 4 _241_
rlabel metal1 s 4232 13974 4232 13974 4 _242_
rlabel metal1 s 3726 13872 3726 13872 4 _243_
rlabel metal2 s 2346 14620 2346 14620 4 _244_
rlabel metal1 s 2530 13192 2530 13192 4 _245_
rlabel metal1 s 2438 13328 2438 13328 4 _246_
rlabel metal2 s 2990 13158 2990 13158 4 _247_
rlabel metal1 s 2576 13362 2576 13362 4 _248_
rlabel metal2 s 3448 12750 3448 12750 4 _249_
rlabel metal1 s 3634 12410 3634 12410 4 _250_
rlabel metal1 s 3036 12342 3036 12342 4 _251_
rlabel metal2 s 3542 11798 3542 11798 4 _252_
rlabel metal1 s 12926 1836 12926 1836 4 _253_
rlabel metal2 s 5543 13430 5543 13430 4 _254_
rlabel metal2 s 5014 12716 5014 12716 4 _255_
rlabel metal1 s 5336 12274 5336 12274 4 _256_
rlabel metal2 s 16146 14314 16146 14314 4 _257_
rlabel metal2 s 13294 9248 13294 9248 4 _258_
rlabel metal2 s 11730 12410 11730 12410 4 _259_
rlabel metal1 s 8970 14382 8970 14382 4 _260_
rlabel metal1 s 9522 14484 9522 14484 4 _261_
rlabel metal2 s 11638 11866 11638 11866 4 _262_
rlabel metal1 s 16790 13804 16790 13804 4 _263_
rlabel metal1 s 9154 12308 9154 12308 4 _264_
rlabel metal1 s 9108 11866 9108 11866 4 _265_
rlabel metal2 s 8970 11900 8970 11900 4 _266_
rlabel metal1 s 20148 12342 20148 12342 4 _267_
rlabel metal1 s 18998 11730 18998 11730 4 _268_
rlabel metal2 s 8970 10404 8970 10404 4 _269_
rlabel metal1 s 8464 10778 8464 10778 4 _270_
rlabel metal2 s 9338 9384 9338 9384 4 _271_
rlabel metal1 s 12282 7854 12282 7854 4 _272_
rlabel metal2 s 10350 8092 10350 8092 4 _273_
rlabel metal1 s 12834 8432 12834 8432 4 _274_
rlabel metal2 s 12374 8636 12374 8636 4 _275_
rlabel metal1 s 12880 10234 12880 10234 4 _276_
rlabel metal2 s 19920 11662 19920 11662 4 _277_
rlabel metal1 s 19642 11866 19642 11866 4 _278_
rlabel metal1 s 19872 16626 19872 16626 4 _279_
rlabel metal1 s 18952 12614 18952 12614 4 _280_
rlabel metal1 s 20332 11866 20332 11866 4 _281_
rlabel metal2 s 19642 16524 19642 16524 4 _282_
rlabel metal1 s 18400 13498 18400 13498 4 _283_
rlabel metal1 s 22310 12308 22310 12308 4 _284_
rlabel metal1 s 24794 12716 24794 12716 4 _285_
rlabel metal1 s 26128 12342 26128 12342 4 _286_
rlabel metal1 s 26450 14042 26450 14042 4 _287_
rlabel metal1 s 27002 15674 27002 15674 4 _288_
rlabel metal1 s 24196 14042 24196 14042 4 _289_
rlabel metal1 s 22632 16218 22632 16218 4 _290_
rlabel metal1 s 22034 16592 22034 16592 4 _291_
rlabel metal1 s 20056 15130 20056 15130 4 _292_
rlabel metal1 s 20516 9622 20516 9622 4 _293_
rlabel metal1 s 19182 14994 19182 14994 4 _294_
rlabel metal2 s 16422 14314 16422 14314 4 _295_
rlabel metal1 s 14950 14042 14950 14042 4 _296_
rlabel metal1 s 16238 9520 16238 9520 4 _297_
rlabel metal2 s 16238 12903 16238 12903 4 _298_
rlabel metal1 s 6072 10030 6072 10030 4 _299_
rlabel metal1 s 7774 12240 7774 12240 4 _300_
rlabel metal1 s 5842 9622 5842 9622 4 _301_
rlabel metal1 s 6210 9520 6210 9520 4 _302_
rlabel metal1 s 6026 9690 6026 9690 4 _303_
rlabel metal1 s 6532 10098 6532 10098 4 _304_
rlabel metal2 s 7314 7990 7314 7990 4 _305_
rlabel metal2 s 7452 7922 7452 7922 4 _306_
rlabel metal2 s 5934 7650 5934 7650 4 _307_
rlabel metal1 s 6394 7956 6394 7956 4 _308_
rlabel metal1 s 8786 7276 8786 7276 4 _309_
rlabel metal2 s 8878 7786 8878 7786 4 _310_
rlabel metal2 s 11362 6494 11362 6494 4 _311_
rlabel metal2 s 11453 6222 11453 6222 4 _312_
rlabel metal2 s 15962 8466 15962 8466 4 _313_
rlabel metal1 s 15318 7514 15318 7514 4 _314_
rlabel metal1 s 16790 11050 16790 11050 4 _315_
rlabel metal1 s 18998 9044 18998 9044 4 _316_
rlabel metal1 s 19458 9452 19458 9452 4 _317_
rlabel metal1 s 18998 9146 18998 9146 4 _318_
rlabel metal1 s 21896 10778 21896 10778 4 _319_
rlabel metal1 s 23138 10540 23138 10540 4 _320_
rlabel metal1 s 18354 13396 18354 13396 4 _321_
rlabel metal1 s 24748 9622 24748 9622 4 _322_
rlabel metal1 s 24978 10064 24978 10064 4 _323_
rlabel metal2 s 24886 9826 24886 9826 4 _324_
rlabel metal1 s 23000 10234 23000 10234 4 _325_
rlabel metal1 s 23276 14450 23276 14450 4 _326_
rlabel metal1 s 21896 10234 21896 10234 4 _327_
rlabel metal1 s 18952 13838 18952 13838 4 _328_
rlabel metal1 s 18216 11866 18216 11866 4 _329_
rlabel metal1 s 17526 11866 17526 11866 4 _330_
rlabel metal1 s 12926 11628 12926 11628 4 _331_
rlabel metal1 s 14260 6698 14260 6698 4 _332_
rlabel metal1 s 15686 5202 15686 5202 4 _333_
rlabel metal1 s 14674 2550 14674 2550 4 _334_
rlabel metal1 s 15456 5746 15456 5746 4 _335_
rlabel metal1 s 8004 5134 8004 5134 4 _336_
rlabel metal1 s 13202 5848 13202 5848 4 _337_
rlabel metal1 s 5290 4624 5290 4624 4 _338_
rlabel metal1 s 10534 4080 10534 4080 4 _339_
rlabel metal2 s 5382 4930 5382 4930 4 _340_
rlabel metal1 s 3956 4658 3956 4658 4 _341_
rlabel metal1 s 7038 5100 7038 5100 4 _342_
rlabel metal1 s 7360 4046 7360 4046 4 _343_
rlabel metal2 s 9062 4250 9062 4250 4 _344_
rlabel metal2 s 11178 4250 11178 4250 4 _345_
rlabel metal1 s 11132 4658 11132 4658 4 _346_
rlabel metal1 s 8556 5542 8556 5542 4 _347_
rlabel metal2 s 9706 2074 9706 2074 4 _348_
rlabel metal1 s 9384 1870 9384 1870 4 _349_
rlabel metal1 s 5290 2482 5290 2482 4 _350_
rlabel metal1 s 6486 2516 6486 2516 4 _351_
rlabel metal1 s 6164 2482 6164 2482 4 _352_
rlabel metal1 s 5198 1870 5198 1870 4 _353_
rlabel metal1 s 3818 3978 3818 3978 4 _354_
rlabel metal2 s 3726 3740 3726 3740 4 _355_
rlabel metal1 s 7544 2482 7544 2482 4 _356_
rlabel metal2 s 7682 2074 7682 2074 4 _357_
rlabel metal1 s 9016 2482 9016 2482 4 _358_
rlabel metal2 s 8970 2074 8970 2074 4 _359_
rlabel metal1 s 12696 4658 12696 4658 4 _360_
rlabel metal1 s 12558 2822 12558 2822 4 _361_
rlabel metal1 s 12696 1870 12696 1870 4 _362_
rlabel metal2 s 12742 4012 12742 4012 4 _363_
rlabel metal2 s 12926 3162 12926 3162 4 _364_
rlabel metal2 s 13938 2074 13938 2074 4 _365_
rlabel metal1 s 15870 1836 15870 1836 4 _366_
rlabel metal1 s 16882 2992 16882 2992 4 _367_
rlabel metal1 s 16928 2822 16928 2822 4 _368_
rlabel metal1 s 17204 2958 17204 2958 4 _369_
rlabel metal1 s 17204 2822 17204 2822 4 _370_
rlabel metal1 s 16974 5168 16974 5168 4 _371_
rlabel metal2 s 17158 4828 17158 4828 4 _372_
rlabel metal1 s 18906 4012 18906 4012 4 _373_
rlabel metal2 s 18538 3740 18538 3740 4 _374_
rlabel metal1 s 18170 4080 18170 4080 4 _375_
rlabel metal1 s 18814 3604 18814 3604 4 _376_
rlabel metal1 s 17986 3604 17986 3604 4 _377_
rlabel metal2 s 18354 3162 18354 3162 4 _378_
rlabel metal1 s 17434 5100 17434 5100 4 _379_
rlabel metal1 s 17848 5134 17848 5134 4 _380_
rlabel metal3 s 15778 9435 15778 9435 4 clk
rlabel metal2 s 21666 12631 21666 12631 4 clknet_0_clk
rlabel metal2 s 2714 8160 2714 8160 4 clknet_3_0__leaf_clk
rlabel metal1 s 13478 1258 13478 1258 4 clknet_3_1__leaf_clk
rlabel metal2 s 2438 10336 2438 10336 4 clknet_3_2__leaf_clk
rlabel metal1 s 12374 16660 12374 16660 4 clknet_3_3__leaf_clk
rlabel metal2 s 16790 1088 16790 1088 4 clknet_3_4__leaf_clk
rlabel metal1 s 21850 6698 21850 6698 4 clknet_3_5__leaf_clk
rlabel metal2 s 18354 15232 18354 15232 4 clknet_3_6__leaf_clk
rlabel metal1 s 21160 14994 21160 14994 4 clknet_3_7__leaf_clk
rlabel metal2 s 17618 8449 17618 8449 4 net1
rlabel metal1 s 11891 13362 11891 13362 4 net10
rlabel metal1 s 4324 6970 4324 6970 4 net100
rlabel metal2 s 21942 8602 21942 8602 4 net101
rlabel metal2 s 3542 14076 3542 14076 4 net102
rlabel metal1 s 4094 8942 4094 8942 4 net103
rlabel metal1 s 2065 8330 2065 8330 4 net104
rlabel metal2 s 26450 8568 26450 8568 4 net105
rlabel metal2 s 2622 6460 2622 6460 4 net106
rlabel metal1 s 2806 14892 2806 14892 4 net107
rlabel metal2 s 7958 10778 7958 10778 4 net108
rlabel metal2 s 8418 9214 8418 9214 4 net109
rlabel metal1 s 16330 16694 16330 16694 4 net11
rlabel metal2 s 7038 8806 7038 8806 4 net110
rlabel metal2 s 12098 7582 12098 7582 4 net111
rlabel metal2 s 8510 8228 8510 8228 4 net112
rlabel metal2 s 11822 15742 11822 15742 4 net113
rlabel metal1 s 12967 15606 12967 15606 4 net114
rlabel metal1 s 8970 8058 8970 8058 4 net115
rlabel metal1 s 2346 13396 2346 13396 4 net116
rlabel metal1 s 7866 12342 7866 12342 4 net117
rlabel metal1 s 23506 6222 23506 6222 4 net118
rlabel metal1 s 17618 5780 17618 5780 4 net119
rlabel metal1 s 17802 17000 17802 17000 4 net12
rlabel metal1 s 10948 7922 10948 7922 4 net120
rlabel metal1 s 8096 10234 8096 10234 4 net121
rlabel metal2 s 24150 8160 24150 8160 4 net122
rlabel metal1 s 17250 9894 17250 9894 4 net123
rlabel metal1 s 15962 13498 15962 13498 4 net124
rlabel metal1 s 11270 13396 11270 13396 4 net125
rlabel metal1 s 26956 14586 26956 14586 4 net126
rlabel metal1 s 14950 16014 14950 16014 4 net13
rlabel metal1 s 3864 17306 3864 17306 4 net14
rlabel metal2 s 1518 17527 1518 17527 4 net15
rlabel metal2 s 874 17527 874 17527 4 net16
rlabel metal1 s 9200 17306 9200 17306 4 net17
rlabel metal1 s 6624 17306 6624 17306 4 net18
rlabel metal1 s 5980 17306 5980 17306 4 net19
rlabel metal3 s 15962 12291 15962 12291 4 net2
rlabel metal1 s 5336 17170 5336 17170 4 net20
rlabel metal2 s 4738 17459 4738 17459 4 net21
rlabel metal2 s 3450 17459 3450 17459 4 net22
rlabel metal2 s 2714 17452 2714 17452 4 net23
rlabel metal1 s 10580 3706 10580 3706 4 net24
rlabel metal2 s 12190 8772 12190 8772 4 net25
rlabel metal2 s 11914 9282 11914 9282 4 net26
rlabel metal1 s 17986 13396 17986 13396 4 net27
rlabel metal1 s 17521 13770 17521 13770 4 net28
rlabel metal1 s 8878 4012 8878 4012 4 net29
rlabel metal2 s 16790 17102 16790 17102 4 net3
rlabel metal1 s 6670 5134 6670 5134 4 net30
rlabel metal1 s 20562 14926 20562 14926 4 net31
rlabel metal1 s 19039 14518 19039 14518 4 net32
rlabel metal1 s 11638 4046 11638 4046 4 net33
rlabel metal2 s 19090 15334 19090 15334 4 net34
rlabel metal1 s 17981 15538 17981 15538 4 net35
rlabel metal1 s 7130 4012 7130 4012 4 net36
rlabel metal1 s 19550 16558 19550 16558 4 net37
rlabel metal1 s 19591 15946 19591 15946 4 net38
rlabel metal1 s 15548 14450 15548 14450 4 net39
rlabel metal2 s 18998 17306 18998 17306 4 net4
rlabel metal1 s 14807 13838 14807 13838 4 net40
rlabel metal1 s 18952 14926 18952 14926 4 net41
rlabel metal1 s 25484 13702 25484 13702 4 net42
rlabel metal1 s 24375 13362 24375 13362 4 net43
rlabel metal2 s 19826 11458 19826 11458 4 net44
rlabel metal1 s 19177 10574 19177 10574 4 net45
rlabel metal2 s 12466 5202 12466 5202 4 net46
rlabel metal1 s 22494 16660 22494 16660 4 net47
rlabel metal2 s 21385 16014 21385 16014 4 net48
rlabel metal1 s 24564 6834 24564 6834 4 net49
rlabel metal2 s 19550 17153 19550 17153 4 net5
rlabel metal1 s 25760 5338 25760 5338 4 net50
rlabel metal1 s 14122 14484 14122 14484 4 net51
rlabel metal1 s 17388 12410 17388 12410 4 net52
rlabel metal1 s 5198 4692 5198 4692 4 net53
rlabel metal2 s 21298 13129 21298 13129 4 net54
rlabel metal2 s 21385 11594 21385 11594 4 net55
rlabel metal1 s 19642 13838 19642 13838 4 net56
rlabel metal1 s 18947 12342 18947 12342 4 net57
rlabel metal1 s 24932 16626 24932 16626 4 net58
rlabel metal2 s 24982 15946 24982 15946 4 net59
rlabel metal1 s 22034 17136 22034 17136 4 net6
rlabel metal2 s 26616 15538 26616 15538 4 net60
rlabel metal1 s 25801 14518 25801 14518 4 net61
rlabel metal1 s 22080 13838 22080 13838 4 net62
rlabel metal2 s 22406 14450 22406 14450 4 net63
rlabel metal1 s 23414 15538 23414 15538 4 net64
rlabel metal1 s 19274 9520 19274 9520 4 net65
rlabel metal1 s 18982 10166 18982 10166 4 net66
rlabel metal1 s 22954 14450 22954 14450 4 net67
rlabel metal1 s 26220 12410 26220 12410 4 net68
rlabel metal1 s 23506 10574 23506 10574 4 net69
rlabel metal1 s 20240 17102 20240 17102 4 net7
rlabel metal1 s 23828 10778 23828 10778 4 net70
rlabel metal1 s 26128 13158 26128 13158 4 net71
rlabel metal1 s 13524 11662 13524 11662 4 net72
rlabel metal2 s 13657 12274 13657 12274 4 net73
rlabel metal1 s 22678 12274 22678 12274 4 net74
rlabel metal2 s 22402 13566 22402 13566 4 net75
rlabel metal1 s 3726 4624 3726 4624 4 net76
rlabel metal1 s 1886 9078 1886 9078 4 net77
rlabel metal1 s 20470 12614 20470 12614 4 net78
rlabel metal2 s 26726 16796 26726 16796 4 net79
rlabel metal1 s 21574 17034 21574 17034 4 net8
rlabel metal2 s 15410 10404 15410 10404 4 net80
rlabel metal2 s 15506 9078 15506 9078 4 net81
rlabel metal1 s 14858 13294 14858 13294 4 net82
rlabel metal1 s 16284 8602 16284 8602 4 net83
rlabel metal1 s 21712 6222 21712 6222 4 net84
rlabel metal1 s 19913 5814 19913 5814 4 net85
rlabel metal2 s 6578 14620 6578 14620 4 net86
rlabel metal1 s 17480 10098 17480 10098 4 net87
rlabel metal1 s 15778 10132 15778 10132 4 net88
rlabel metal2 s 25162 10812 25162 10812 4 net89
rlabel metal1 s 20654 17068 20654 17068 4 net9
rlabel metal1 s 25801 11186 25801 11186 4 net90
rlabel metal2 s 17986 8568 17986 8568 4 net91
rlabel metal2 s 24426 10047 24426 10047 4 net92
rlabel metal1 s 2622 12240 2622 12240 4 net93
rlabel metal1 s 10120 16014 10120 16014 4 net94
rlabel metal1 s 12696 10574 12696 10574 4 net95
rlabel metal1 s 12466 11288 12466 11288 4 net96
rlabel metal1 s 7498 5882 7498 5882 4 net97
rlabel metal1 s 26266 6834 26266 6834 4 net98
rlabel metal2 s 9430 16490 9430 16490 4 net99
rlabel metal2 s 874 1095 874 1095 4 o_digital[0]
rlabel metal2 s 18354 772 18354 772 4 o_digital[10]
rlabel metal2 s 20102 908 20102 908 4 o_digital[11]
rlabel metal2 s 21850 942 21850 942 4 o_digital[12]
rlabel metal2 s 23598 1078 23598 1078 4 o_digital[13]
rlabel metal2 s 25346 908 25346 908 4 o_digital[14]
rlabel metal2 s 27094 534 27094 534 4 o_digital[15]
rlabel metal2 s 2622 942 2622 942 4 o_digital[1]
rlabel metal2 s 4370 874 4370 874 4 o_digital[2]
rlabel metal2 s 6118 636 6118 636 4 o_digital[3]
rlabel metal2 s 7866 636 7866 636 4 o_digital[4]
rlabel metal2 s 9614 636 9614 636 4 o_digital[5]
rlabel metal2 s 11362 772 11362 772 4 o_digital[6]
rlabel metal2 s 13110 636 13110 636 4 o_digital[7]
rlabel metal2 s 14858 772 14858 772 4 o_digital[8]
rlabel metal2 s 16606 636 16606 636 4 o_digital[9]
rlabel metal2 s 26266 17187 26266 17187 4 rst_n
rlabel metal1 s 25668 17170 25668 17170 4 ui_in[0]
rlabel metal1 s 25300 17102 25300 17102 4 ui_in[1]
rlabel metal1 s 24748 17102 24748 17102 4 ui_in[2]
rlabel metal1 s 24012 17102 24012 17102 4 ui_in[3]
rlabel metal1 s 23460 17102 23460 17102 4 ui_in[4]
rlabel metal1 s 22816 17102 22816 17102 4 ui_in[5]
rlabel metal2 s 22034 17418 22034 17418 4 ui_in[6]
rlabel metal1 s 21252 17102 21252 17102 4 ui_in[7]
rlabel metal1 s 18538 17136 18538 17136 4 uio_in[2]
rlabel metal2 s 17802 17425 17802 17425 4 uio_in[5]
rlabel metal1 s 16928 17102 16928 17102 4 uio_in[6]
rlabel metal2 s 16514 17425 16514 17425 4 uio_in[7]
rlabel metal1 s 2392 14858 2392 14858 4 uio_oe[5]
rlabel metal1 s 10442 17306 10442 17306 4 uio_out[0]
rlabel metal2 s 9798 17248 9798 17248 4 uio_out[1]
rlabel metal1 s 8326 17306 8326 17306 4 uio_out[3]
rlabel metal2 s 12742 15861 12742 15861 4 uio_out[4]
rlabel metal1 s 7314 16218 7314 16218 4 uio_out[5]
rlabel metal2 s 15870 17255 15870 17255 4 uo_out[0]
rlabel metal1 s 14720 16218 14720 16218 4 uo_out[1]
rlabel metal1 s 14904 16762 14904 16762 4 uo_out[2]
rlabel metal1 s 13938 17306 13938 17306 4 uo_out[3]
rlabel metal1 s 12926 16762 12926 16762 4 uo_out[4]
rlabel metal1 s 12190 16218 12190 16218 4 uo_out[5]
rlabel metal1 s 11914 17306 11914 17306 4 uo_out[6]
rlabel metal1 s 11316 16218 11316 16218 4 uo_out[7]
rlabel metal3 s 14030 16643 14030 16643 4 wrapped.o_busy
rlabel metal2 s 9982 16864 9982 16864 4 wrapped.o_copi
rlabel metal2 s 10810 16864 10810 16864 4 wrapped.o_cs_n
rlabel metal1 s 13837 2448 13837 2448 4 wrapped.o_data\[0\]
rlabel metal2 s 15594 11577 15594 11577 4 wrapped.o_data\[1\]
rlabel metal1 s 14766 10438 14766 10438 4 wrapped.o_data\[2\]
rlabel metal1 s 14766 10098 14766 10098 4 wrapped.o_data\[3\]
rlabel metal1 s 13570 10098 13570 10098 4 wrapped.o_data\[4\]
rlabel metal2 s 9246 5831 9246 5831 4 wrapped.o_data\[5\]
rlabel metal1 s 12650 3536 12650 3536 4 wrapped.o_data\[6\]
rlabel metal2 s 13156 10676 13156 10676 4 wrapped.o_data\[7\]
rlabel metal1 s 14122 15402 14122 15402 4 wrapped.o_data_valid
rlabel metal2 s 15042 2244 15042 2244 4 wrapped.o_digital$17\[0\]
rlabel metal1 s 18124 1530 18124 1530 4 wrapped.o_digital$17\[10\]
rlabel metal1 s 19044 4454 19044 4454 4 wrapped.o_digital$17\[11\]
rlabel metal1 s 21160 3910 21160 3910 4 wrapped.o_digital$17\[12\]
rlabel metal1 s 15226 4046 15226 4046 4 wrapped.o_digital$17\[13\]
rlabel metal1 s 13892 4046 13892 4046 4 wrapped.o_digital$17\[14\]
rlabel metal1 s 19918 816 19918 816 4 wrapped.o_digital$17\[15\]
rlabel metal1 s 5934 1734 5934 1734 4 wrapped.o_digital$17\[1\]
rlabel metal2 s 15134 3366 15134 3366 4 wrapped.o_digital$17\[2\]
rlabel metal1 s 7130 4692 7130 4692 4 wrapped.o_digital$17\[3\]
rlabel metal1 s 8510 1530 8510 1530 4 wrapped.o_digital$17\[4\]
rlabel metal1 s 12834 2312 12834 2312 4 wrapped.o_digital$17\[5\]
rlabel metal2 s 11546 1632 11546 1632 4 wrapped.o_digital$17\[6\]
rlabel metal1 s 12190 4624 12190 4624 4 wrapped.o_digital$17\[7\]
rlabel metal1 s 14260 1326 14260 1326 4 wrapped.o_digital$17\[8\]
rlabel metal1 s 16238 1734 16238 1734 4 wrapped.o_digital$17\[9\]
rlabel metal2 s 7866 15096 7866 15096 4 wrapped.o_sclk
rlabel metal2 s 20470 8092 20470 8092 4 wrapped.o_spi_address\[10\]
rlabel metal1 s 18676 7514 18676 7514 4 wrapped.o_spi_address\[11\]
rlabel metal1 s 24196 6970 24196 6970 4 wrapped.o_spi_address\[12\]
rlabel metal1 s 25484 6834 25484 6834 4 wrapped.o_spi_address\[13\]
rlabel metal2 s 25162 6324 25162 6324 4 wrapped.o_spi_address\[14\]
rlabel metal1 s 26220 6426 26220 6426 4 wrapped.o_spi_address\[15\]
rlabel metal2 s 24978 8908 24978 8908 4 wrapped.o_spi_address\[16\]
rlabel metal2 s 26542 8092 26542 8092 4 wrapped.o_spi_address\[17\]
rlabel metal1 s 22448 9010 22448 9010 4 wrapped.o_spi_address\[18\]
rlabel metal1 s 22540 9146 22540 9146 4 wrapped.o_spi_address\[19\]
rlabel metal2 s 3174 8772 3174 8772 4 wrapped.o_spi_address\[1\]
rlabel metal2 s 21390 10336 21390 10336 4 wrapped.o_spi_address\[20\]
rlabel metal1 s 20056 8602 20056 8602 4 wrapped.o_spi_address\[21\]
rlabel metal1 s 17572 10030 17572 10030 4 wrapped.o_spi_address\[22\]
rlabel metal1 s 17112 10778 17112 10778 4 wrapped.o_spi_address\[23\]
rlabel metal2 s 4186 9690 4186 9690 4 wrapped.o_spi_address\[2\]
rlabel metal1 s 3312 9554 3312 9554 4 wrapped.o_spi_address\[3\]
rlabel metal1 s 5106 8398 5106 8398 4 wrapped.o_spi_address\[4\]
rlabel metal2 s 5382 7140 5382 7140 4 wrapped.o_spi_address\[5\]
rlabel metal2 s 5474 7174 5474 7174 4 wrapped.o_spi_address\[6\]
rlabel metal2 s 6302 6562 6302 6562 4 wrapped.o_spi_address\[7\]
rlabel metal2 s 18814 6749 18814 6749 4 wrapped.o_spi_address\[8\]
rlabel metal1 s 20332 6834 20332 6834 4 wrapped.o_spi_address\[9\]
rlabel metal1 s 10166 2584 10166 2584 4 wrapped.player.buffer\[0\]
rlabel metal1 s 5934 4250 5934 4250 4 wrapped.player.buffer\[1\]
rlabel metal1 s 5014 3706 5014 3706 4 wrapped.player.buffer\[2\]
rlabel metal2 s 5934 4930 5934 4930 4 wrapped.player.buffer\[3\]
rlabel metal2 s 7866 3876 7866 3876 4 wrapped.player.buffer\[4\]
rlabel metal1 s 9660 2550 9660 2550 4 wrapped.player.buffer\[5\]
rlabel metal2 s 12466 3876 12466 3876 4 wrapped.player.buffer\[6\]
rlabel metal2 s 12512 4658 12512 4658 4 wrapped.player.buffer\[7\]
rlabel metal1 s 13662 6800 13662 6800 4 wrapped.player.received_samples
rlabel metal2 s 15502 13039 15502 13039 4 wrapped.spi_flash.address\[0\]
rlabel metal2 s 20286 10880 20286 10880 4 wrapped.spi_flash.address\[10\]
rlabel metal1 s 20424 10778 20424 10778 4 wrapped.spi_flash.address\[11\]
rlabel metal1 s 23138 11764 23138 11764 4 wrapped.spi_flash.address\[12\]
rlabel metal1 s 24426 12648 24426 12648 4 wrapped.spi_flash.address\[13\]
rlabel metal2 s 26266 12036 26266 12036 4 wrapped.spi_flash.address\[14\]
rlabel metal1 s 26588 11662 26588 11662 4 wrapped.spi_flash.address\[15\]
rlabel metal1 s 26542 10778 26542 10778 4 wrapped.spi_flash.address\[16\]
rlabel metal1 s 25024 15130 25024 15130 4 wrapped.spi_flash.address\[17\]
rlabel metal1 s 22724 14790 22724 14790 4 wrapped.spi_flash.address\[18\]
rlabel metal2 s 21390 15028 21390 15028 4 wrapped.spi_flash.address\[19\]
rlabel metal1 s 7636 11322 7636 11322 4 wrapped.spi_flash.address\[1\]
rlabel metal1 s 19918 14586 19918 14586 4 wrapped.spi_flash.address\[20\]
rlabel metal1 s 19274 13940 19274 13940 4 wrapped.spi_flash.address\[21\]
rlabel metal2 s 16974 13124 16974 13124 4 wrapped.spi_flash.address\[22\]
rlabel metal1 s 15502 12308 15502 12308 4 wrapped.spi_flash.address\[23\]
rlabel metal1 s 7314 10132 7314 10132 4 wrapped.spi_flash.address\[2\]
rlabel metal1 s 7268 10778 7268 10778 4 wrapped.spi_flash.address\[3\]
rlabel metal2 s 8142 9316 8142 9316 4 wrapped.spi_flash.address\[4\]
rlabel metal2 s 7958 7684 7958 7684 4 wrapped.spi_flash.address\[5\]
rlabel metal1 s 8832 6970 8832 6970 4 wrapped.spi_flash.address\[6\]
rlabel metal2 s 11454 7004 11454 7004 4 wrapped.spi_flash.address\[7\]
rlabel metal1 s 14306 8602 14306 8602 4 wrapped.spi_flash.address\[8\]
rlabel metal1 s 15042 10132 15042 10132 4 wrapped.spi_flash.address\[9\]
rlabel metal2 s 13570 14620 13570 14620 4 wrapped.spi_flash.fsm_state\[0\]
rlabel metal1 s 6348 13838 6348 13838 4 wrapped.spi_flash.fsm_state\[1\]
rlabel metal1 s 12052 14042 12052 14042 4 wrapped.spi_flash.fsm_state\[2\]
rlabel metal2 s 7590 13702 7590 13702 4 wrapped.spi_flash.fsm_state\[3\]
rlabel metal2 s 6486 15640 6486 15640 4 wrapped.spi_flash.fsm_state\[4\]
rlabel metal1 s 20240 14382 20240 14382 4 wrapped.spi_flash.shift_reg\[10\]
rlabel metal2 s 21114 13668 21114 13668 4 wrapped.spi_flash.shift_reg\[11\]
rlabel metal1 s 23276 13158 23276 13158 4 wrapped.spi_flash.shift_reg\[12\]
rlabel metal1 s 24932 13498 24932 13498 4 wrapped.spi_flash.shift_reg\[13\]
rlabel metal1 s 26772 13362 26772 13362 4 wrapped.spi_flash.shift_reg\[14\]
rlabel metal2 s 26266 15300 26266 15300 4 wrapped.spi_flash.shift_reg\[15\]
rlabel metal1 s 26312 15334 26312 15334 4 wrapped.spi_flash.shift_reg\[16\]
rlabel metal1 s 24886 15878 24886 15878 4 wrapped.spi_flash.shift_reg\[17\]
rlabel metal1 s 23000 16150 23000 16150 4 wrapped.spi_flash.shift_reg\[18\]
rlabel metal1 s 20516 15878 20516 15878 4 wrapped.spi_flash.shift_reg\[19\]
rlabel metal1 s 18584 15674 18584 15674 4 wrapped.spi_flash.shift_reg\[20\]
rlabel metal2 s 17066 15572 17066 15572 4 wrapped.spi_flash.shift_reg\[21\]
rlabel metal1 s 16054 13974 16054 13974 4 wrapped.spi_flash.shift_reg\[22\]
rlabel metal2 s 15502 15300 15502 15300 4 wrapped.spi_flash.shift_reg\[23\]
rlabel metal2 s 13202 9180 13202 9180 4 wrapped.spi_flash.shift_reg\[8\]
rlabel metal3 s 14122 11747 14122 11747 4 wrapped.spi_flash.shift_reg\[9\]
rlabel metal2 s 3818 14756 3818 14756 4 wrapped.spi_flash.timer\[0\]
rlabel metal2 s 4186 13940 4186 13940 4 wrapped.spi_flash.timer\[1\]
rlabel metal1 s 4232 12954 4232 12954 4 wrapped.spi_flash.timer\[2\]
rlabel metal1 s 3864 12818 3864 12818 4 wrapped.spi_flash.timer\[3\]
rlabel metal1 s 5750 13362 5750 13362 4 wrapped.spi_flash.timer\[4\]
flabel metal4 s 27256 496 27576 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 20540 496 20860 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 13824 496 14144 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7108 496 7428 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 23898 496 24218 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 17182 496 17502 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 10466 496 10786 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3750 496 4070 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 27158 17600 27214 18000 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal2 s 846 0 902 400 0 FreeSans 280 90 0 0 o_digital[0]
port 4 nsew
flabel metal2 s 18326 0 18382 400 0 FreeSans 280 90 0 0 o_digital[10]
port 5 nsew
flabel metal2 s 20074 0 20130 400 0 FreeSans 280 90 0 0 o_digital[11]
port 6 nsew
flabel metal2 s 21822 0 21878 400 0 FreeSans 280 90 0 0 o_digital[12]
port 7 nsew
flabel metal2 s 23570 0 23626 400 0 FreeSans 280 90 0 0 o_digital[13]
port 8 nsew
flabel metal2 s 25318 0 25374 400 0 FreeSans 280 90 0 0 o_digital[14]
port 9 nsew
flabel metal2 s 27066 0 27122 400 0 FreeSans 280 90 0 0 o_digital[15]
port 10 nsew
flabel metal2 s 2594 0 2650 400 0 FreeSans 280 90 0 0 o_digital[1]
port 11 nsew
flabel metal2 s 4342 0 4398 400 0 FreeSans 280 90 0 0 o_digital[2]
port 12 nsew
flabel metal2 s 6090 0 6146 400 0 FreeSans 280 90 0 0 o_digital[3]
port 13 nsew
flabel metal2 s 7838 0 7894 400 0 FreeSans 280 90 0 0 o_digital[4]
port 14 nsew
flabel metal2 s 9586 0 9642 400 0 FreeSans 280 90 0 0 o_digital[5]
port 15 nsew
flabel metal2 s 11334 0 11390 400 0 FreeSans 280 90 0 0 o_digital[6]
port 16 nsew
flabel metal2 s 13082 0 13138 400 0 FreeSans 280 90 0 0 o_digital[7]
port 17 nsew
flabel metal2 s 14830 0 14886 400 0 FreeSans 280 90 0 0 o_digital[8]
port 18 nsew
flabel metal2 s 16578 0 16634 400 0 FreeSans 280 90 0 0 o_digital[9]
port 19 nsew
flabel metal2 s 26514 17600 26570 18000 0 FreeSans 280 90 0 0 rst_n
port 20 nsew
flabel metal2 s 25870 17600 25926 18000 0 FreeSans 280 90 0 0 ui_in[0]
port 21 nsew
flabel metal2 s 25226 17600 25282 18000 0 FreeSans 280 90 0 0 ui_in[1]
port 22 nsew
flabel metal2 s 24582 17600 24638 18000 0 FreeSans 280 90 0 0 ui_in[2]
port 23 nsew
flabel metal2 s 23938 17600 23994 18000 0 FreeSans 280 90 0 0 ui_in[3]
port 24 nsew
flabel metal2 s 23294 17600 23350 18000 0 FreeSans 280 90 0 0 ui_in[4]
port 25 nsew
flabel metal2 s 22650 17600 22706 18000 0 FreeSans 280 90 0 0 ui_in[5]
port 26 nsew
flabel metal2 s 22006 17600 22062 18000 0 FreeSans 280 90 0 0 ui_in[6]
port 27 nsew
flabel metal2 s 21362 17600 21418 18000 0 FreeSans 280 90 0 0 ui_in[7]
port 28 nsew
flabel metal2 s 20718 17600 20774 18000 0 FreeSans 280 90 0 0 uio_in[0]
port 29 nsew
flabel metal2 s 20074 17600 20130 18000 0 FreeSans 280 90 0 0 uio_in[1]
port 30 nsew
flabel metal2 s 19430 17600 19486 18000 0 FreeSans 280 90 0 0 uio_in[2]
port 31 nsew
flabel metal2 s 18786 17600 18842 18000 0 FreeSans 280 90 0 0 uio_in[3]
port 32 nsew
flabel metal2 s 18142 17600 18198 18000 0 FreeSans 280 90 0 0 uio_in[4]
port 33 nsew
flabel metal2 s 17498 17600 17554 18000 0 FreeSans 280 90 0 0 uio_in[5]
port 34 nsew
flabel metal2 s 16854 17600 16910 18000 0 FreeSans 280 90 0 0 uio_in[6]
port 35 nsew
flabel metal2 s 16210 17600 16266 18000 0 FreeSans 280 90 0 0 uio_in[7]
port 36 nsew
flabel metal2 s 5262 17600 5318 18000 0 FreeSans 280 90 0 0 uio_oe[0]
port 37 nsew
flabel metal2 s 4618 17600 4674 18000 0 FreeSans 280 90 0 0 uio_oe[1]
port 38 nsew
flabel metal2 s 3974 17600 4030 18000 0 FreeSans 280 90 0 0 uio_oe[2]
port 39 nsew
flabel metal2 s 3330 17600 3386 18000 0 FreeSans 280 90 0 0 uio_oe[3]
port 40 nsew
flabel metal2 s 2686 17600 2742 18000 0 FreeSans 280 90 0 0 uio_oe[4]
port 41 nsew
flabel metal2 s 2042 17600 2098 18000 0 FreeSans 280 90 0 0 uio_oe[5]
port 42 nsew
flabel metal2 s 1398 17600 1454 18000 0 FreeSans 280 90 0 0 uio_oe[6]
port 43 nsew
flabel metal2 s 754 17600 810 18000 0 FreeSans 280 90 0 0 uio_oe[7]
port 44 nsew
flabel metal2 s 10414 17600 10470 18000 0 FreeSans 280 90 0 0 uio_out[0]
port 45 nsew
flabel metal2 s 9770 17600 9826 18000 0 FreeSans 280 90 0 0 uio_out[1]
port 46 nsew
flabel metal2 s 9126 17600 9182 18000 0 FreeSans 280 90 0 0 uio_out[2]
port 47 nsew
flabel metal2 s 8482 17600 8538 18000 0 FreeSans 280 90 0 0 uio_out[3]
port 48 nsew
flabel metal2 s 7838 17600 7894 18000 0 FreeSans 280 90 0 0 uio_out[4]
port 49 nsew
flabel metal2 s 7194 17600 7250 18000 0 FreeSans 280 90 0 0 uio_out[5]
port 50 nsew
flabel metal2 s 6550 17600 6606 18000 0 FreeSans 280 90 0 0 uio_out[6]
port 51 nsew
flabel metal2 s 5906 17600 5962 18000 0 FreeSans 280 90 0 0 uio_out[7]
port 52 nsew
flabel metal2 s 15566 17600 15622 18000 0 FreeSans 280 90 0 0 uo_out[0]
port 53 nsew
flabel metal2 s 14922 17600 14978 18000 0 FreeSans 280 90 0 0 uo_out[1]
port 54 nsew
flabel metal2 s 14278 17600 14334 18000 0 FreeSans 280 90 0 0 uo_out[2]
port 55 nsew
flabel metal2 s 13634 17600 13690 18000 0 FreeSans 280 90 0 0 uo_out[3]
port 56 nsew
flabel metal2 s 12990 17600 13046 18000 0 FreeSans 280 90 0 0 uo_out[4]
port 57 nsew
flabel metal2 s 12346 17600 12402 18000 0 FreeSans 280 90 0 0 uo_out[5]
port 58 nsew
flabel metal2 s 11702 17600 11758 18000 0 FreeSans 280 90 0 0 uo_out[6]
port 59 nsew
flabel metal2 s 11058 17600 11114 18000 0 FreeSans 280 90 0 0 uo_out[7]
port 60 nsew
<< properties >>
string FIXED_BBOX 0 0 28000 18000
string GDS_END 1938054
string GDS_FILE ../gds/digital_top.gds
string GDS_START 383892
<< end >>
